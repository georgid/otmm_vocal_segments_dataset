BZh91AY&SY�6� �_�Px���������`?�ML��E P� ��`�6�Ja$MFT�h��&����4 h���M!P�茀 `���2b`b0#L1&L0i�)��2h  �  �&��&�j�&M �h2 B�����O&C F�i��Ѧ@�
���%"*9 h �H3��)��x����U@���7�$��K�*h��=�(�"�d��io��C���~���+����moږ$RI$��I$�	$�KQI$�ĝ$��������Q������t\��(���EK�N�!RtQEBJ�I�B�RPvd@Y��n�jA$�Ij)$�X���J�P�IRIJIBI/�q�޺ES�59��U���F_'�+���N��s�����[xZ���(\�|��C9�v6%nL,ORvC������$�1��0K�<H 0vޢ��3'kC��77����C.k�#a<�XR3���c(U�2u���->S���;�n��­��/w�2ŭ<�d��8[2�/���ѹ3a"nH�
��\�Iiġ���x�R���ͧh~���
1����Mi1�}b�0����K��N�{	��b�7.۸[�)Hgi(q�!�Qv�yc�U�^aF����Z���}חX�X#B8u"��κ�_O�����$�I$�I)���[��I$�I$�I)�S��nܗ���_f������Ǥ��>C���v��UUI"���Ȝ�(x�އ�Ȳ,�# H
�����k�o�ߞ '�e�.���`��@:���������zl�a���X�&|�K��� �Uݷj2jR/6�%�|�}�ۆ�`2����`G���RA�y~6.Jϕ���'f��D'V�(P*1�j�]]3M�X����<)e���v����p 9��Y�є��;,���s�,�u��q�qsQ\�`TD�'X$�Ě�@�2�����3��`4B��O���wadP�'Ha�fQ�|N;^��9aT�H@�����j�q� s�zjI�3���Z�O�&�`�M�m�E+�ѱC��ŭ*\-��tGAb�i	�"���f�|��UUJ�O�4����$8��u�n�Γb8��_�-�pQD�圞�2r\dQ�Zr�����YIW]����B��5�KKL��'M��c �)��y�Dh��6�_���v8s�-��]�;�����͏W�y�y�C�����]\�5uS��c��# i���q�Y�Z�Q&85wn� ����3�s���]�O(��W�Ȕ���ǣ��+�����r�i6���?(<��!��G�~m��r��bH;{=�@ʫ6]y�.H���@�x��8�����T"�J᝼���䦥�wK��g��q02�By��l�{Ȁl���vVwf�~	�y���{S������|�!���g.�+�FD�'���DU�;�r�z�o'<�Zdz. �(�eVV��ʚ�ײ��50�f�K�o��������;ص��[Z����cr�dT�)�[�fbi�x�<]i<k��C�����f:)N)lT��X�؟���8���ɔ�c���ޫ���^��S�)�v�OS��nޱ��	 ����/�k�w&�To������4����r�|f7�k:��"f+{k�o�0��fBNgј��󚳪6��{q�m����)7�Y��X��u�o�r��%�.:m���I,�3T�.�w�qS�*<��A�+Ψ�\g���t��y�<"��梶V�h���ܫr<���&�=]R��p�7u���Ð��������}����j�찇��>���濷��i���y&��.z\�9�?+؅]Cڌ[~^���=�d3���=�>d�Ȩ�d��Ș�����W��Q���%ޣ���:���P�G�6Xa+��*;ݿuz��׀}O:�_3�J����:��Yݸ��}Y~�2��g):¸���Ezut#�'���W��aD�y����5����]w�z �AWu���|�ʈf�C*���|�[۰{�H��^����i�c���1�u�,лԶ}]_�_=���"�}���G��Ec�A�]]�)&�W��g{�Ļ� Ep  
��J�i��>^��� ���� /�̯{�d#�y�g7Rڵ��R�Vj�i���� � �`  
j�� �    M��6  @   
b�L���B�p�7�Q`D,��R[2в�^�J�Y
b�u�6T�(��1{�T�*�)EXH7��.R9@~Q�p..8�����*q�M��@II�MW���c�~����6k��.�>~�N��1���ۊ:(l�ҥ���LQ�*H��W�J��M���'�uTXʖq$�/�����:Q��U��Cّ)!�-؛���Sh�k��B���b� W��9Ϩ72'�dL��Ъ��pT�ʘ7jsV ��Ctٱ/KO�#�=���O�=�Ē@�-EG���D�{${l��:����X�[�H�}�rѴN�.^e����(���- $@	�C�P����@��	�dd��%)�\c2�+8f@��o���e��<�7|}'1�6j5 �*@��UB�
H)) � )-�43���05������w�:�!�:��İ� ,�}=�7���dp����W]]��f6�_�p�7��� 1�&�a��f�hжA� �ݬ6������F�|y&�U^�������P���ZI̟\�P�lN�$���Η���2;Ht�/
0:�� ��MfDGqdv� �p��a�ZIcv�y��d�`:!C��p׼.�!�j.��SDͧ 4��5�h���^f�1�-�jY� B��-���(E:î���	:=םB���u����\:�t��f\�Qb��ݶ�,�߽7(�#d���ۺ6	� �D�����iUXp�@
�<��ɣU�H�㴒C`wM��&@� ���
,B��Yg�Cs��M26kپ������b����Chj�uT>����HTx�]�� P� op6Nͺ���A������b��?��n�fǬc���bc����M�� �a��u��~�� ,�xh�3.i�'-!����|֐�갷 ���-��H�
F�!�