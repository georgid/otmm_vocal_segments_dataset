BZh91AY&SY�J� <W_�py����������`*�|`  �z "��WO�s��4�� I   	]X � ƹ�h$ �  $ ��r�h�6BP�*��d�UQ4�d��0#	�L�LL5<@)JTi��h@`��� jy��*mM䑚@  4  S�jS!j�� 4 @���T��6ɔ��i������d�A��"P"h&&�&Jx��)�P�=M@��?n�D ��@ �q?�P@���u���{}Y_�f��2���o����n���i"�Q2���}���������L������|?	�P� �  :����$e��%9�#,
9Nw���yRu���Z���-;ΰ� �Hm2q�Õw}泫��\���wx�Ю��s���{S����ovޛe�p�B:Ī�t뼻�����s����:����B�!�6�84	�KX1YB�P�r���u����i���뮷�2�8B�B�u�iV��;�Me�!B	K�t$����;�.j����]�h�Zk9�#P� �%�22�.RY�7��)A뤥*U�ڳ�^u{���K���j��8D��!�FDe�4�m��9Y1�!F/w������<l�M��!��!F�٧�eU�!Ga�N;��T���Y�.��f��ޙe�u�!B9 %*rBv��g�Fa��b���!�q�Q�l�)���z�!�Zm��F42���_�R����\�^fG�n(�J��T�Lv��!y���ءm (mP��l?\S/9�w��`��I_�rL�SY3����
G���
�L����'��V�<v�t������tUS�ӹ�DN?L=�ܰ����6yH�ж/nKe5t�*�x`��"���j�J�4�]�8�B�]���۝�5U��3XF��\`��en�����q�R����1�B��^�T��I�Jj*\O�q�̮�,�)x�Y��L�+�}
{,bH6�r��F�@��RS�P�+m��^����ۊL#�ov�x��kZpDe�{5L�k#ec�Lkq���PPԥ:E�f&L����)(���Zl\*��g��Ǘ�=��f�lT�ڔ/�v��su�M!a�qi��\�ɑ[�ml�ܚ�X7Q��Q�&�4�P�ڢ�2q�b�J��rL\�R��.��)XW�#A�,ѓ$Ye��R�.�0�M%kkٮ��m��=Y��Q8�.Ķ�ʵ�M�jL���\AE%����:c)�uL���z�R�W%��o�I�q'1�Z�r�kM���y[���oOn�⋎����M�}�3�g����("}�Ěb�臶�ől�L붬�(�T�[�`8�ۥ�
�"i��v�Id��
IUɒ�#�<��
E���e�v�u�E����8A��WFĤ�.��8Dwm�qI������H���c�B�@Fڕ�:�c�$�5�u�?0�O�����>�}?�v� *��ʊ�f�T�(P�����(��(��(��(��(��(��(���*�*QEW^�oH!ϝ�y��]�bU���\A�qW@�0�"b�\�L�0Pq�==.�Íg�����S q� q� q� q� q� q� q� q�F8 �0 q� q� q� q��`�I�f�d$�X�c7tq� q���~�WWu-.�-y�(��K�`�uD���}�pv0[�A®HU�\^G_J@P ��o�'r����t&�Î������� �!�D���\555�\�\555MMt�����^Ÿ�ݜ<@��WZ�N�~׶�M�PTb������mg�0�@"���fV%9u�6�ὐ6hb��J���T���˕�9L�)ƘT�{[ekj∹00ؙ�EjHI�\8��F�.�7v٬�'~_��&�F����(x� h�r��gyI�qE@�!i�Bi�c�I�Vɥq Ңf�.ͫ&�;��=Cffs�g+����&�� ����#���b�£�b0g����
*"؊k&���	�m�M�iz�P6��!�I@�*�@�؜.uV�I�4qE�i��f���1gH��cm^�*n���Q3l1��9��鞚,��i���C�U����r�KT��| P�=�˹�qdQ��0E'uB�Ü͜(^���I��L8��������R�6������6��b��*��YNwj�R�W��������h�gEL�Jw�*V^n�`�/0�\�5X=�p�ݼ8*�z 	5�F��8y:�0������R�JԩZ��x�N'<N'����q*T�N<x�N=~�d�r�B���ߖ%G~-�79�IS3p���|}"4�FV����lE�d (��O��ߖ�y�_+���ل|��ƾs[
�4����{Q)܉�"�����U�?f�����cH�Ͳ�I�e�Ș��؜W������jA�D�؉�͈��|��k���)�6��L�b��H��`*k��|�۰%7%ͱW#5������u�#V�).����O �ǀ�UM���v>,�rɪ�� O�����>���A�N>���/U�]��T���Bc^�l)��`�Л���q=���T���2���s;_���VCD�������#�:�����	\7&c��\;cGg4| ���j�؞�s?s_?epr���Sىc^fU�'�][R�Q�����{¤Զ6�PJ��xI�D�>��&F�p�������q�R�Z�*W�ǉ��q��8��q�x��T�<N9�<�|		o�y&��A5E~Ϛ˝�VTE�Cyo ��W`�Di�C������X���ɺ0�����4�#$iI#��EZ�W0�߯~�_y����hU�#�>T �}���Z�~vz⧘}��U(iwa�y���~ o�?\��{	��1�H=xD�Ҋ� W��`��(�%z����_�'�*"f���#E�����"������-.���˂"�X/+�{~�֨�H$I�RLx{�%��0Gݮl����.*Ns�V���ϕ��v�`��Oz�v�$�:5��[<#�������c���EO�x��?9���_}�N_���S����}�xT �ﲁf�$ݝm��
j%�l�����P����T$CEu��)����M��~� g��;�� ����.���m#dxO	u�=eހ��B�]�T}��}��J��r�}<N'�Ǐ�ĩ\�J�+S�''g�0:��o��Ӯ�ބ�2ݕV�o#\m�İ�{����� ��?�91<]!���Y��|`:�$���ꭡ�#-�P | ^��{׸<��~����&b&\O\.0�ͽ���Ə������$���0��b�c��U_l��d����#�j�6Z���� oǿ*���ڙ��e�0=���I;�F�_}�X�!w2��V8�_��"��� ��Y#l_�D.����CJm�eG����>T��ݜ��b����">)f+fr��<Ǽ7�i6	�cT9f[2OJ9���a�V�Ң�	�w)��������E�p~���_]*u�;��FD��v��Q	}�W|�'�8�f\���?Uݿ��N�K��T2\@���=�{�� c�m0<s�u�GkAz͔���m��������\��Z�J��S�������x��\�R��z0��]�z�I'3��31�2>��"Kq'�M��5����u��%�(+�����Ec����������?l���q�d�\d��&$�E�<�]4�<��Sw��>wk2m��عs�'�a-&���4�Lژl� A&���?Q�A^�F�d��b5%W�I���S����d`��\�V��I�W=�x���ݱ��d|�v~�D h���+,|�� ���Wg$/�P��"+���	��m���{*$j�����'r;���Y��'�1|d�{� ,��=՚!�,��5�ܢhfy_O�s݇�z�lt�	�R]1���vdx���5c�1'C�]ո��	Z��W*]�{;"ھk7jd�e�߻�c��6���_�ڂX�H-*�h(p���]j�������%r��#�M����d8cf�z��h�<�~B����vr�P6IC޹���DJB��2:*����+/����)�Ӛ湩����R��9ǉZ�jW+R�R�����*z���C*��hӷX*v�D���'���/s���٦�KG+ɧ��i�F���ɍ�2Vl6��W�+6��FL��p	Q!�����CC�3�/ L�a�$�ɉ"��`?O����^��C���M����)����V�U-�=�W��G�.k���b��3��S{��1�ܣ�cX1f:A'���*�����7%���:�n��;��;lg�d��+�Õ����z7�1���Tqa3Վ��^�R�1�Xv^w*�\]f����"�2NV����)b�aS<.F/ӹ�$>�\���P���BX���|�U�/g�X&�Q��cR�$�ӌr�����u^�?�����R��VުP<''���2&�.�f϶�pٳ���F�!�r`8��x�BD(0n9�&с����t����ʺb�^�꩗�G�*'(Cl+���SP�Z�*T55�+R�jW+\�W�|��B#1ATD�c$21����H��׾�����d~���<����Cqу��6oʆ'Vş}�n=I&v񫴃N�<Ti��D5 �A��D�+M�B�#V���8��"��Fo�4�CqsR� ����� ܇6��-uf��z�ػ;*l��%�ʸ���n�LA��x�au.�[u��T�E�w*4v�h�����������%��p�Ƿ�'64E�ē&���UFe�� ����HA��a?ei������gޓ�{$W}[�a�SV�ݐ��q��M*� d�v�G��6|��}|���y:�)	Fb�.D�@���g��;�p�B1#0(�_���	˱b>��鏄M�d,H �1���tm�K�f��ל�{��ή�������,�̸�=`q�Y0�nm׹r���+f�C��נ��3 �������Lτ�����555�=�jT�R�Z��V�JԮT�Ns�5�9���h�"^���3�5��܄��
��v��=�L�.V�U��B&�l
�{�@#��)`׀�7�v�t���cFIJ��Ar��>��q����FJ8G�����hb(�(JP<ES��H3�m���R*z�ۜ�վ�U��0u�Q�{b6��su|�d5��ɇqCv2iI�y3�p�,,�t���Rc8]�uu���f2Ɯ*Q�5�@n��u��:��v�����<�!L6�����2��F_fG���G�w��N��O)�"h�:������ӳ,��DE\�}�v��uEc�[$��C	�H��zɗ���a���i?yP�;���:&T]�ۍ�G��l~24������\�+R�J�+R�ʕ+R�r�*y�'[��iqې�m�D�TJ R��
�<���������wS{z��*��u(�|�D<&���ɝ�\_G2r1Ju
�b�I#��� �����o�{��/>YlQ�3k�}��8cT�p���G��'XQ�o-U�SB�P�mbNpBOf�I��I�L�b�,����|	i3Z2�v� ��O&�"�.�}��'�� X>���>6N\=�Cpsy��4"���O8`�?�����N��I�a�H,@"Cɩ9>�6*���P����q��V#	:������/��w�}�F���qt۞�؍CV�#�I
`�9��`.�����h� ����޾cE߉������D	��ʔ �Z� ,� ���G��l��6rxEĄ*�	)n�����(�]�\' k�Ve����Yb�r�r^	�,�3hb콾|��3='#�>S]s�T�J�+��Z�r�+R�r�;����9�2$��⋃���Y�Z�vK$�;��:ifż�p���<a=DѣaD�%SM�8*�*���/(9̩��C�M���SB6b$PN���Q��#�Qº=��t�"
 ����gIS�2�lƚ��/��[�+���}����ڛ�n��k�#���G��qV��{�.��ۋȳ�{;��v�:X��y�TpF� �e����+7�T��#����ٻ�"�S�*��!}_M<i��z�r�fk��3vG�{��w�#����������d�.&N����b��S�iwV[���O*>��m̅B>�?zDNp�>�F�S��q�[��D^�aSY5@���t���&�uUU� 0y������%�Z0Oͥ�r��_
!�t�w��z��!�p�E�s ��1^؊�����"���(�2�� ��d��U�]*)�p�q \U�q0s	1Z@	D�R�!|���ŀH�*�0�.,���@��HQ(��
�!"�(IE	�bQ�P�cdT2��[�`� �"��!`��
�%�$ J�J�@Sc
�!U@�A��V�d$��@�Ȩ�������KE�:&�2H���`�)" I "��&�������<�S6�9P��Tܠ��A=��muḷ�N����7$�������Z {ӓ"��w������� 2���A3��oo�POo� =[1�����I$�I$�I$�EUUUUUUT�UEUUUUUUUQQUUUU1���Ш'z�r�]~�;�6�X7��}6����5j���~��m��,eHl2�Π��@z��ݩ��u���* d��w���8}�|�=#�@i����H`[��M'=���ۤ�L�Ԛ=��p�g(> �d����o����[�����f�jHb"*j�
��~A6�*Ot�.q�r�����˖O��-������yF���U��^}��L>���7{x�ft�EaE��}sn{�<�BB�b VH��"QR`*�!$��B�) Q$!@��̋
L	"�@g(��E܋Z��)q�1�x,/�S43	�F����P*f0�DGwT����"�H�+�lq�ϣ��qק��׊<Cnκt�f,�8�d0��}e�<;�������5ve����V�2���K�t��3���
��"���v_l����հ�t����l��t|̍���I��a��]�4�#��P ƽ	�
Ȫ!BA�Ӎ��I�9�X)^�^�^�O8{�A�8�eR��p�Pp� ��zAׄ��n���	�Q�dU��*7}�����8W|���&��Jsba�E��T ��P�w�nQl�҆��T+F���@�D˯$-�Y%��p�V�:�]�X�iD+�f?3�B� Jo7�:s�]���u6���ʏ���4�"d�ɣ�p���3}��|�\�VGbv�6csg	A�~�P�a:�c�æ^wr P Ǔ���OyR�
���C�N�P ��\朇�2���t���Wf�6�Im��P�0����-r�uibYd����|N�.�����c��V��]���N����kv�ɇ��FA����YpP ɚ��b��1���4��Wq@�2z8p�sju��;"��*�v-�L��&���@ϑ��T$	�g/Qc�=���}���(	ۏOn44w�` ���r���A��<`���p���E9�{k����6��G_�rE8P��J�