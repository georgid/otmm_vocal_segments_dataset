BZh91AY&SY����r߀pp���f� ����aj_  �`� 	}��   
 )��f�
 ����f�  �� ��                    �A@                  �� ͓ǧv�eV��t��ˮ�U{-�U�uZ�[Y�>���+F�q�2��7�in���/z�π�� R�E)IS�N��\T���:kMV� ]��Mm���C�� uӱ0�R�M&�5���v�PҌ� � ����Fu��-.ݵW���Z�l��K.�*Ӵn��tݭ�כ����E��G�W[�z��^7L�[[�ݽ�<U �@���ݩn;{w��ס�[{�٧���sU[m��f���z�{ݽ��Uջ���k�-��Wk�� Y.��������宖��4t���z۽R�omWosU]��8�sJ��S��+Kj���(P����קKqE�Y�n�s���ۮ�j��J���΅�:Q�2nUmm��ݗ����[�3u�WO �A����[w<�=�u�k��Or��h���oS�������u���{��.�6�ʎ����k�Dx�P� �Ig�v�'���j��:�*��j��u+7]F-K�M]K�Lթ[Xz��������� ��cN�+�sT7������ӗ��V��uQ�^��خ�;�Q��ԹNN�Wn楥�� xT�(�(Vq���]Z�۴7R�u޲�v��׷���wKv�m؜�]t:;V��Y^xS���x        E?����P d�    
���b�R��      D�2�J�)�� � 4�� j{%$5Jj�0!� ���4 O�"�*Q���b`a
B�#M&$�!�hd�4�ڟ�K�?�����������G��=�^����AW�� ���US��U_�?�U]+�����S�EV�ʫ�ɠQUW�?�e���DU��?��lA_�����ID_�����Q2AJ_��2@R�_��A_eA2`Q�AhW�QL�_d r=���Ur
T=�E� W�����J#@)�
>��H#J�/��>¨�*��)��)�)�)�)�)�)��)�b��������������Oc$J�T�X�b��d��`4'�B��>ڑ=�%}��=�!(=�=�=�=�=�=�=�=�<�<�<�|�<�e
}�=�=�=�H��d���4��"{"d�"e��j�r�eOu���{d)�b4��H�� {d)�{�ȯ��S��=�}�=�ܯ�K�+IB
 ��׏����?:E�գ�g��u�I��}��;�����[��#���_�x����U�2��ߪ*�Ɵ4����n��S�����n��C�c�	�O$�j�[;u��86��;��#O9�sv��Od�w�47i��to[7�5$t�4�������bxu�@Y�ouӽ:���gw��vu]����Ǯw�ϭ�,���C�US:��*�u�O��qz�����7G]�z��	�NBP�'p�����C��2S$3~=�]u�u��Һ۠��ވ��<;�ݷ��p���<�7`d�&F���	Br�
N��JvDd9)HP�%	[��J�BP�%&�,C0J:�w�2LL��'<5<x�3[�7��2ujd&���9���j�4����(2͸������]f��s�f�t�\��f7tv[�����S�rr6��F�rM�A��%:[ 3!��2prR���drt��:ڴf�4:�#(rR���JC3�I�]9�V$��C%�do�Xo�w�n��ӆ��^h��.�fr����.�̮��N�1������Q�+9K���_N��Ĵ|V�L�{5 �JS3� �N��8y,^Fp��;���e������t;��L��d�X�Rd�A<���a,��隵3�Q��Ԇ�!|�����zG*[1J;��`����\2��12�%�tf���6�A���Gq��י�]wo�s&ǡ�N�+Hdγ�RGOF>��T��N�#�:�K��'E��(���i�2���o���÷���Gg\5��z��Ϝl�<�`�^:��:�,0-kF��֮�����O%)��M�a���0���}�u������h �N�]n.d�o`w8h+��7AZ�۝���u�k�&ζ����y��kgշ��<f�^C��cZ�M>XsH�3�f�J�U�v���|K�r�uQ�W�f���C��}�;|��:�:�M�Zdt$�D㪘("<h �#E���	�0BR�r^��R��Ґ��1p4)�!Bkx&P���)vj�;��`�	����!5�0rC5:	�J^K�`aN@u�S��12���m���ֳ:<"-fs�'����C�DYL���2/'Oy��R�DD�
$�9��j�gP�.A�������&�p2�$(z}�m�sBXd�AO�g���`A���P��R�{xwg��w��my{��k��D	�Č�!���r�׺0�&��Ɉ�Jq�;�t�b(�ms�<�z�Z���B��kRA��k#����p�ڠ����j�$(J���	�̻�N�3D�2�N�5"f�h�Y�=��C�Nk�(JR��9)H{<^�<�C�J{$(JR��+ٵ��s9&�Q�sQ��Ԙf�Yh"�	BP�'J#L�Pd9�ݢq��`8��f�HP��!BR���PL.�%��HP��!BR��)��MHP�)�	q�&;��M��oG��%	BP�%	BP��Hd%	���$:���:�ب���Д������0�a�U���w&N�֧!(JY�R%)ԛa(�6x�y�ӄ���oX'P�9�&�(q3Ӷ�jvɐ�`�	���%�9!I�>�OQ��$3��A����n:hM@MT;���'���vk��f<*;��8t�v�݉����;��i��K�3��ݭ�wc\� q��jq*X����j7���ΓC�p:��)
�Ԇ�2S�ƫ
�z��U*��W�8����N�u�xc�i 2
�;��[`��W3(og���:�z2r`�k����I>r2u��d�찱�s<�� F��n��՚;N�~�_Ҽ����%(12�N6C�!���,*ϸ������⠻|�YMl�珝��Ϛ8��C�7sK�	"h����yּ�\�μ��Y��t�(��ʝD�a].�X���9�R+�p�y4��Α<���x��h^Y���&	���ZxM�2������'.c�Awͦ�d��� ȝgq��y�뽆�F\'���U��̷�0ٴ5���'%)
%5!B{nS�
�JC!2|��f�]��J�^NU'RÜ�>W<B��;��#�12ٳ���\�GG6u�c�Ö�n��05��,8�k�R���l�Q�=���w�&���T�lp��d{�ĲR�i��A/7�����p����̃���P�)�oF��ӌuy����nӽ��u���h���F��^'PabA��`����$��䱱�ɛ�u���.{�z_��w�A�8t��Ѣ�ՠ�|�t�k�%�3�Y�3I�^D�ϓ���#"� �=�Z���"0�( �ֈ3F�J�`��G�ߙ�"3�8p9�J04���
B)
Y����
H��u	Hj�N�:���7��{��0Ѵ�p�r��[���'xq����-�/��,��3����b�%2�@i�͝r�[��6Z��A��P�!BR��	JR%HP�%	BP�%.��0�8l=����f��zw�P`札��]��h�\6�7��fy`Ж�&2H ��"�VHP���a����U989`aA�o�9�`Nda�C$��F=����5j(Өrr� �n�X��uh�<=���ČM����sn���Q�u��z��o<C8B�Mu@d6F)A�`@K	JPC!!Y��il�r.@fI�f���0�1�u�[7��Y�މ�7�Ѿ�u���:������ڕC������]�U��qNK�~�I���/W�����M~�[��w�ۧ����[� �L�o�˲ �B�fj�۳F���[BDꀄ�����`�j�Za`�tA�Y	�:$)Ö�k�ѣ�ȋf<4uX�	�"+NJM�d,�X�c8���������f�,�o[���bd	BPU�ҙ	�L�ή�9���e*wR��2�fV>V:�Њ�T�YT}�bl����$��.����/xYI��'��������t��_�
��(E��
U��Lwk���r�՟��3�]7du������5��}��s��S�v!�> ��W�����)�]���9&:5�$2
I'no���W]o	�/�V���IUyW\��,>}��9�~$��%�%�]8�g���<{��d�enӲ�i,�Oy��GAei#mp��F�YUE"�}�����E`�bz��=|�d�u5�ɞ�����Y���W3�]]VT,�Y-���fK�p�T�|�R�}�o�oy� ������`	X�5�P�
���7R�C�!,R�]A��X0P���4%	JR��I������	K�M��
BՂd�&&.%��Gd9�[4atv΍vE��NÅ��=Y��A�e�0��M>o�:�<u�	�	̃���r4�W�`;��L��2\��3#v:�ӓ��C�ej�.�(JR��)JB�{Y]vl����׼Ce.HP��!BR���fh�����9��F=9	N�1�FbY���1�;3�7�������%,L��(<M�0w������S�氹��Ef��"њu!Bu���øJR��+�C �15��{^�(�)I���0���9�	����^��k6�h�jzx��(J��R��(N��2t;�1��)S���W���,l~M��/%���8vq#�/<�hֳ݁oD[�����,��P�Ԛ�!3Y�u��0 �F<��>K�	e���}�$���n��} J�P��8�����L�}�l}]��5��z��d����P�%&>kq�1��l�������`r�C��M�6�!������ꐃ�����m�jB�ԧ�%)���i�R��	JRg=�^�u��#}�k�wo^fxgz������5	v�%���Ar1��8O��M�\J9.V�!Ԇ�#�ѫ�;cX�:5�!;�:\��[�;��]��o|����������b�"`�p�Zt�AD��x�!C⮹�a4�'S��0 cA�0������d9Q!*u)I�u�tI���Rt�pHFA�ζa�1ah���=��(JR��%)HR�)������ײ��9|�1:�<W�W�Z.�}w�tt���mA����rR�\�5�t�ĴkaʋVư2�y_����{��{įҟ����.,}��e����^��Ω���,��J�)���g���>R6�� q�ECqCr��ƎPە����������w��?����S���������{��u�&����h�������������������������rA�F�b���������������bI��7$��M��AAAAAA	HPPPPR_IАPS�𐄅��AAAA|(((((((ܐm� ؠ�����������������蠠�����Ē&t��`:�绗pܹώ�v��fY��rŉ����Z%��6Ɩv޽���O>h�X�d�kݚ�T�lPPD���Ӝ|ȳ2l�AAAAAn�+���t��C;����Fs�#����T�wp�ms�R�N��fd{wt���z�gJe�6$��n6�r�!�ys�n��3�wt�&)/��H($�$����K�6�-���6x_IАY�9�������O,m���C�iw���$nkݚ���������y�ޱ�gH�c}[���޶���.��_O���h�
�sH�ӹ_E�{�Z[���b�ՙ���F�S����ROu7ݵ�As�7��v���P��r�3sT�-á"t6�ĒU3$xm������n,�Γwk���X�����XH�nOV�&�o7}.���Y��]ҭ߉�@h����D^)hW��d"Q�V�j��Ro"AUAu��szI�a_�������HB旟ws{�������t���ה��1.3�8���g1�AAUAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA@�H�ؠ������������������wt�((((ܐm� ؠ�������������5蠠��������������������5��


��/�����������������������������������





Scm��


























��5��


















7$��׭��𠠠������������T����
PPP~�ޱ��AAC��nH6ܐlPPSٙ���������������������������!v,� ������������rA��b��T�yY�




0IC�����*����������������3&�nH6(ܐlPPPPPPPPPPPPPPPPPPPPPW5A�AAAAAAAAAAAAAAAAAF�yvܐLQs�|Ԓ�

































~��
� )�P�yc���$�R�ſ�zI��J�Ի�R�v���QK:S��%3wV��\ݪ��$����Tk�鷝��.����U7���L�(6$�$���Zk;�7�i���̋#HK*
n+ijGC�ˍq�LY�;5fn�n�*Hm�1g:� �8(('iշ�]7��(KQ�PP^��3$�&u�n�mn����W��mU,�R�� 1@�1��6�8���{�c��lBD�����$� �s9��ݫ��(8(�,��S�6((((��Ď����{�PPPQ� �rA�BS���[w��l#&s�����.���rA��.���̇J�s'�5�|-ݪ2gx�P:�c�Ax�~��I_H�����7R�޵ܲj�F��[���uH_{�}{�}�3�{m��Zs@��9���	�"��n�����q�W�`!of�tA�·1n��mg��Ut�˻�w^�n�� �1AAAAAAAy�d����w
:l����9��9��t;�w`�,I }������n����ď�|��o
v�p���k�]������ݱ3���=cb����1�{wD.}�n������1$�wi$��`��wM��];X��*M�[:O=��.s��1�*�	����;wwM��ݕD��s��7jWu͗���%~M��{�c��|ߘN��q�Ty�N�&ܻ���S���?������\��˃v�o伯swo��Y�^�w^�=`�گ������s�V�Y�����:���*vמ��2v��}w72Enl��*^U��z�BMoz�q��m߳�uI����b�.���R\L}�n�wPI7����� ö�y���Xw��woq��}��o�֎,~q�_j����P�⥷���Էu]���k�=we�����A�AAA?Wpj.�U��[U�*e����s0�Է����[���8��Rݬ�g�z����q��wy���r�To�H>��>���b�� ����-bӟj�������k#�ܽj�|��J�������M��@��q�w:��.������;�~F'�X���y�� ,I�!z ��(��m���%��"��vwl���H((�P�@M�>c�c��|��b����"�GHWwwkp���J���I���ۺ������[n���M����WsS�
��]c5�ּއ!g�ıo#[�k5�݋�L���E�����v�߯���wR�	]�.+Kc�66((��C���Y�L�N�2PMd��6�	���|NS��T��[�sUN�{)�%�¥V���b�z�cm�wR����g��;��^:�H��w^a���jȄg�s�mAAb��-�+;��껥)t~�ˬ0^K�]Ш�R�Sm;�wBX{�w~u�V�
�ꁚ��xy��l[�}ò��Zȯ�^um����g�1nNޓD�Q-�j��9�kծ�ѷ��]��+���U��i��ًvnw>���5N�����zM��,�@|�Ux�9D�
rɵjk��;����;�=��sb�O� �����vj+�����C� ���]�/T�s(�{�Qs4(�$����[X=�1#311]�y5AOW����u��N��wvb�����u�w���� 9�C�绱w



7�m��ڔ6�]�U���F�p˺�ż��Vx�c�Ε�z���sr��b������V�fh�s'U)Z���AAF䂹�Y�fK7T<���2��H)���������PPPP��㸻�/��O/R�qv��LPPPPIbI67�ۗ�ɫ!���{2^=�ٛ'q����4Ffg11N�λ�6�$���<(-�'(((ܐlQ� ��k�"����y)5LI!AAAK����!�$�m�-��|(((g\��껣t���}��I		�9�3������vvww_c�bK�w�N���Mm߶�M���̇��$���ܙr��H��7��ݒ\��b�̂𐄛��=$!�����X�B�S�QJm�6&k|���mAAAAAAAAAAAAAA{��e쬃�AAAAF�M��ַq76s�[m_fzfkG���L��(�$��;���PR^�揅�6�rk���RqS�lMLQ�Q��fL�ؒ2�3�^I��[�ZA���MGt�il���in2�[���bIAABgD���I��q�Ÿ��t��TW�N�ض;m��L>�~MmwWwnuҫ�vvYcD��w+��ɩ>̏��-ܭ��65ƭ{��y�띝�Vʻ�<z�\���$��,۫oK��ڪ�����:�wZ���I/��^�M1+��L�Z�ui�URXIM=B�Eu�@M�Wv�_YW��7�eJ��d9�.���̸�����3��/f���1�ޮ�}����׾R��W&t����=�!n��uz���=6�F�.�%�n:͓��;�լ�����]�˼��g��=���lHXUԷ�Ã��*aڜn�.q%<��%B��SX*�u㦛�/�wυ׻q��.{m�����N>g9,�uQ�-I���g���ޛ7ϋͽ���Wj�k�*��{��^繆O
���\W˓�G*��Suo�q�gj��ꗻUJ����u*�9�ݽ���d��Jn&��������]�l�t����n�z�N8�伭۸��g��Z�̣Frq��M�<��Y�4����<pT�@��Z���gWC��쾾f�E�,�X���Ӫ��{�U��園EU�]�q���E��亮�ovEٶ��f���۹^yy�˕E��;8���j�/�G"�3�_>�	



PPV͖��.���V��	�[���:g�p1���u��lY��o��lj�hjS--/��g�7�G�]�3i-��I�$�����xTc}�(j�F<�����y,#�c~�t�2�m&�ջ�vԶ��>�N��}�/D�#Ryfk�Bg*+����\��(#�2OI��tn����/�T��[���AAAC�o���_


[�����HX�BI�^[��ےD��wu�R��Z�W�N���6!!N��ܜ3]�ws����oݕ�r�W�6s#x����ɍ,��ܻ0�ֶ�
�3Xؠ��wwb�wWv誳8�s�g11AAAAJ��f\��e�{�%S�����,Y�%)��%��r@���lX���3I�T��((x PP򂂂�sX("j���'��M�UH]�:�\��P�n��u��+w:BU









�ǘ�������<��k��wwvR���W)�$��-6�jݱ>g1<ܭP;wL�M�llSL���$�|Y;�ࠡ�M31:�V�]{�6�lLPY�9���o��lPPPPPPPPPPPPPPQ�*���$������������r6�Po�co��ؠ���n�^�����I�D]���5�>�m	C3GڵC)�c�����Z�ٙ��$(L�&t��z����$�o��:Ǜ��I�x�e�d�tv��Z�t�	�


7��ƥ|�cm�ے�	�wuU��l��`ؠ�޷�i,i����$T�(���އ7Y�����/���ESb���� *���$&t�HBB���\��t$n2�]��y�f
:E���Az�BX��"6�7un�J�����UP29G^_%�wl/]gB8�����MP��AAAAF䍸�s9��
]ؠ޷�lPPPPPPR����AAM}��8<��o������������˽swON�&Ul�)�����-�1#������]��5���'
7$;�k̳0�ūw5����w&�ؠ����������6�7t�7M���C��~�ū_=}���& 
׵ZA�AF��ے1|((U.�	�$�KޭGn�]��PPPPPPPPPPPPPPPPPP���Ŗ�_W�]V�֦�q\�m�ë������1!@Z�鏳��As�fǉn�g��']9�H���z�M�B��z�������$!!AAV��PPPPPPPPQfܩB�˳W,�sfd�Ē����K��[��n�N^;�wG�1	
:En6(ܙ�{�[�܋�����㠥݊PQLP陘I���)ݻ��]�J��9�җ��i�-`�ΓLP��v�I��Y���frНRv��k��mޛ�pl�vz�G�w#9�����[�LR�o�՝�ǀ�n���@�0^H����p�7.�oj_wwP�#�|�x庥��ﺷ��|�+ۼ��	����X�<j 6
�;ns�U绻��0�)��y�nf�J�!���@h�B^���Wǫ~߶q�PR_U	�7���rı�{>yدb��6�7`1shv���ff@k��R�7�D���׵\yn��ɦJ���}�%�k؍{�Pm��Ww16����U�������[����Y�7rn��o&`((gvwV��]��ɗ�c��h�+�~kg����f6�ω3;\΋�ә�˻�����ӷ����T�n�&K�ܛyZ��ʵ+I��l���oa8�t���w~<�U4���Av���{#2�6z[��֣ymʔ^�k�AAAs�mn͛7wtkfǯdx�g{og_Y�@k�t��̹�,MUR�nH��F��n��雒���f��%�$ 
»�enog3�nu�W��X�� ���4�9;�}����vT[iR����h$����ъ��D�OR�'��c��Bz





HBER���������`������B���	V�)���Bt��Y��\zޥ�c��_g����Q��O�;噗o_n����ؠ��+��J]ݙ2���'=xٯ`� 
�-��M��u^�Z�\���>��KJ��Z�/u5�+3꧜cyٙ�q���f0�җuĻp��Ȳ���Au�w]ٙφ�h�H�wi��I�U�SWe��f����x��;�ۭ݃����n�@�m����Q�)Uy-4� 	�A��V���ۉg��Y��Xm�btI���Nÿ��7m^��bQ	2<��ě�q{6����}:�9���P�s����b�;;;�  ���rl��I���p�v��LPPPPPS�����Wu�;��{2�q���Z�B�����u��[lHLo[�6((((((.����g:*�-%ʭ�����Ė��$����OKkv

7$ K�ů3���繑K��̼��Cd���G� ��ΉjDcb���%���_Z��&����������/�s9��e݈J����n��'����v,�����Ē��6ܐlR��>�|}�;�kTlu����7�#: cX��LPIbIwwwp�TI$��t.G��(z��b��\��*� d�S���{���m��#< (.)�7���BCT�k�����߿~��߿"��g���A}������������� ����H"��_������������+�9�w� ѵ��"�ب�b/��x��U;Q�t^/`��G^
	a��"G^�o���
2"���YB (�OAl=@�JfFA��A4�� +�4%)CLL�
��-"D$$R*KJ@�QD10�!CJPH�2�!�K�o�_@Q�a�1D��mQ|4
�A(b��׿Pb��ׁ��]����үH;��\B*=v���肅�bb#ۊ	�� S�WAU; DQ�TC@�^����3$���B�@��J�D�HA,���z�>��4�=
����4 'N��]���!�Ȯ���U΍`���+��u��h���4!�'�><����v !�*|T:ڣ��?�����բ���S����p?�*a��A�� Ȣ �H� �(@�� R$�RФ`�l����g�[w��<���kÔ�g��|]߇������[��� ��]tF�,I��#�j�͋��M�\����*�UVڪ,*��]R�� TPuYp�T��V|ip5LT!�a���n!�ggU�j��*�H[���;"����������'Z�(73��s���d�n/-;��55���I�8��=�ôd獻��DC�I�=UW���G��]�a�WJ�Aad���[խ�a�6���r��t�=�i\\��ڻ&��v�s�Z��%���bMv��!B=�ΎF-MS���U!�c��s���ux���vӵm�rk��@�/F�g�;^�'3�ik89%��bő�F\���ꡍ�v%طchьj��f��>��2U�d_���=Ћ��U@�U<;@y��������z��y��36X�BP\r�|�3��y��|.p��6�G
�-����2s���N���a����83u[k';��M3n�H��4WB?y$�d�5杶2[�XJ�><������9�؂󝺰1xﭜ�.���I:����Ev�g�8�޶8��a���W��O��E8�.6%���ypsr��Jڗr۪ܽ�O&�5��/,�ӗ�Ӳ7V.�z�{���a�vx�1p�������t�R��J�բ�sݿc��q�t�ϣbO=�0p�v�w.%�ab�q,s�Ϸ�ﭾN�����a���A�˹v5d����<�Ѧ\l�v�<�8�}����u,���VH.�j�4�f)M�J��EEʎ�`g{�|��}�p}l;����Iqu��l��]�S�R��7�M��h�9=����T�CSy���Iv�@�\j��u�[n�0v�,��֍�9�P]e]�����X]���T�1�
RH�Տ3��t6Eq��y�=��nf�(�����eZ"n����{vnx�#l�S(��=w��0��*��}��5��U=6�Y�����(�z��'jJ�i�ƕ����2(�I� ��X��s�J��.R�۔����h1s�v�u�������j�.���X\���NW_�8��+�*���$DDKk!�U78d���YF��{4��u�m9v��.A�X�����R]N�PbJ��a�s����D�h��Q} ��;�� ��|�:��g��x�۸��@!��  [�U㚄�8�3��vz�`�p�A-�Y!��U����y�Ғ�j![��VÜ��|��Sc[�|��۶�ez��t��JN�Ձv₤� ��YAի#}�}�ӥL�u�9}�Q�L��Q���nz��6�ԕ���(;�h�ꈈ���2!��*I
K.��pقaÝX���c�8�f��F�N�:h�c�[a�UA0��Q��.�l5��z2Y�j�;����dyf��:����6U2B���\p-)nnYӪ�Nͧ8K�t�4�$�vA��vws��T��We��oɴw�k��=^q5QEvتݩB������of�Y�v�,J�f]�n��Q!u����ָ�ϟ�=.q{�Ý�Z+��2��%]�j�0r�ݱ�7���gu���ّV�,�����OR���R�vy	IN9m;eȝ��ίZ/���=+փ=�i,����D��-�Y5�wv�d�g�VIݴ`��d���hr��m�HQ�5�\����v# ��ed���`-*jbn3.�Iɸ����{���}UT�V�H�1"��WT�
܂;�X��&�����2&E�p�CgT���&�q�i���rI'����	�mV����E&���rp�v�[�+8�uJ�Et�{T�رIa�k[�����#�MM�u��m�r$cW����m�*�O�gwG���X�c�\��w$9(K(6z�`�`s��e��4�w=�tugK�~{���
-W$9:7��+�[�UsSwSVe]��ƛV����V�����=+ր�*���΋�Q��Z�T]:�+���`v{��AOR�/^C��eM�%U�Hӥr"��,Ik�ܡq��jT���)T3�ӒL�D�wwad��fL�vр��b��t�8�eδ�H�� c:�
�0���h����;�`s��,.uz�U�J��"R���Ց0���͞��
^�
҃A �*�� @J4H����O�_(E����zX�ezĽ��6�n]�:�:-�����{<f �l8�{��;G��7Q�R�S�*R,Zw6ꕧ3j�,������r�����#��K�M˰�{<X
�VF!@{#x8D��m������wU\�D�w3}��4��,�]V��~ܷ|���Z�=Q�Zq���K�J�G�\=�a�{�V:���Wum���="�:�n�v450��΋1܂�o(5+f��M�~��RD�ˢSEȭ�����3˾�$����ua���y���r�sWe�`)ꕄ���S�l�K(쥔p�]Ez��۸��ӹD,s�ŀ����&!�cv��.�g�6X�$�TJ0i�]s���0�>�Xuw����Q4).�ʥ]@P!S��Hj � dR���s��Հw��H��L.�Y�"�Qd��\�^���ԛ�J�ܜ�%~�㞙S+2���i��g��5n_�No�8{�'7�ޞq49QE��n�nQ����+����W�{�J��Ia$���F�R��{�֢s�R].�-r�]6��q0��A�Ӧ�n�^�)��A���-�������T�:ͦ�axh�����m��\�AGr1ͳ+jgjP*��b$Վe��C(ĺ���#���m(�������
�+�|�bNQv��n���yV�_Z��v�"U.�8L���BZ��-h3��{
�r}?Er_�'7җ����=�� ���H���Xe�_����G���I��p��T�D�]�3ySU��ov��$�4��js|��Y���g�˺�=A���9������֬�V���٩�Q�us3�Wq�����Zw�^���ڄC�Ry��-(C`����v�Zv���Maw	]{��B���	K��f����&���J�r��g��i�:L���/$ͦ=qΖ�{NV-һV�:P ���ݗ��h�����S4K6e� g]���M��]5c	N�U׍�b�?��~��}�ӋHY�#f[��$�s���I�ϟf�m��jM���^Xe�Wy�xy�P����|i�s�o>��Z�Jf�&�Mڿ^�O]�L�/�ӛ���~���4�L����2��x����9ɾi�ztsk�yw;ԩ�5NU�� �H�����lY��VY�4�`�(A�m�$
6*I���{��W9�^+9�����~���-L�.yqcs�a�33����ee��ߧ'7�n�97�u׌�y�ڃr�J�զ���=�}W����݊M�����d�u?T��3�z�/Ǭ����'7�Nuɓ6�R�.���vͽ�W���������&~֜�s���$E$cQ8�
��]uVeU҇����&zَ��������~&`(���a�uZϗR��[��?|����k���歽�ȝ$�b�hm���_��s޺�:��s#��O�!��X{=�@]�֜��<�un��-�O����'���u\�Ve��]�vg�m��ū?DD}���b"=^�	Lz�[c`��A�e�K4"Y�c��l{m��qbfa����s��fm�rtQJ[�4��d���5��/R'P��"G2n����t8�ԁ�kZ��T�;��5��(ئCA&dm0�`f��͒�٘Q$Y����('H��Ѳ�$.A��[N��������8V�V�m6�H0yb� ��e��+5�,��1�# �����EJ��P	�]�df)�(��j�b�XfB����ϟ]��f�y\hܸƎq��1�c mm���Wh�[�J�]�8�;n2XSk�$@�pV�
Ц�rh˥�j4��`Q.t�S�0�&0p�LcɌc� �Lc֘�%���m1�Q1�`b3l��� �c�1��Zֵ�sěv��N��[��]�\$�؄MV���r;�,v��x����:+��U��Z�/mcu�.��pF8��VB�wZ,Gigvݷ�:B����@ܘ91K�s	�����U�,Q��R�{mi!cD�M��8��V�VK�q�硱��ݥ�g��Mrʘ�9J��-V�K�]s��z妫m��O/l�8.ڕ�ZAv�F� �EC"�+*馹�^2Ί7��.�`��a���"]�B�[�T`Z2�Q�4@��
��7�l���m�p��vݓ�C�)L<d�3��u�k���\�AFՆ�����Ƃ8�9����Dv�v�N�:��kt�jڶ(b]p�Yխ��3��r@P)X�Pjפ��\f�vC��t󺺙�S8خM�ŗZ�T2�!��3v��B��Z�ķ��I����CS�^��V���q�ڧq! �]tr&aF�N` �Vj��#�A�Z�@�DZ)s�^�����tu�mٮ��LVݜX�6�4�m,���ŝk3�L�]m�[D���Ε+e���O�/�ۊ� ��_Qe��"� �Њ�i@!�4�!h;��R�����JO�{���)�=�r>3[5�p�{�����JO.��߰:��;�^��R����5��=BR��{��-"�����Ҍ�X}P�n�IJ˿�	�	����P5f�w5��+5�SYt��ۏ*1�:6�+-Y��y�������JR�~�߹�(Ol��7���:��ｍ�����9�n���=u�"p��\��k�b�g�):��w��HО���}�dwg�`p��r���k_�kBR��~��ֳ[�ԛ�3������R����o�L�����~���)Jw���قR��w��~��R����\�Zټ�p�s��oz�3�R��w��J����يQ�I�������=�m��#�z������_�U`�R��W�JR���}��%)Iמh��N������s�䄇��C�
�Ѿ����ʗfzv[X��n)(-V�����[�e�;\'J�c�1�ﺸB���v1g�{F]\�lك[���w:�N��W&ѫ�!�I.ԓ�Ϣ���кU�ۣg����lr��s;�p�VD�8���e�9뱣V�o�I�����I��||fZ�۲J-6��wg!d�|����s�9-�^I������ڢڷm�3�u�.�FW4��e���>}���':����Kߚײ��{����3{���)�t�t�	m�J��K����)J}���	JRyy����%)ߺ���r����߸=JS��~�V��d��uowe�vr���y~��JS�=��R��￴{�R��%��}��#d�}�����4���g-^f���d�@О{���A��h���=3Z2S�~���JR��ϳ߰z���̽m|�� ֵa���%'^��~������o�L�����u��JR�y���	Ht}祣�f�|:�:�Ff�ftn�'P����5)G���%,���m�t!��!cH�5s���3SDK��9����Y�ל�S�}����Ol��y�߰:��ߏ��u�Lm�']{=��&�[(u���΅E��(;�M�0&��kg��O�����Nx6"XmA��)]�1p���Pkt�zy	���/'Z3[��>������N��!�e����&�-�{���eꔥ'�~���JR���_}�jR��|׿buB^y����3ꥺ/jR�R�aT��t�Jˢ꺔��>�o�`��'�}�������>������О�I�����n�wd�v��=����d�����'����f��4%)I���{�R��<�����W��"��mʺ��) �&��R��L�ϵ��2R���=��JR�y���)JRw߿o�:�������\�������󑳒�O�??��uK���h�fa�����Z����*�x�,t$/RQz}��\R��뿴}�R�K�����}A�VwZ݊�Pn]a�av�9�%\��q&r�9�0Y�8���%)ߺ>�����<��buBy����	@�uy����)�</O�do\Y�o9�fsyqJ����g�u�����%�f����}��Cԥ)���'�G1|��g�6n��I���3�z:�f��N�)O�����%'מ��ǩJS�tk�MJRu���N�)����W7p�Fo�kz�W��'W�{��:��>�_[�%);�߷��K�	g���)�}���{��\z���Fk\��Z�7R��~{��`����������'�z.���uu%W,if����߯�I�(���kW�iMBRyyy��N�h�=?>�۴�vI��{ބљ�.��	F�����Clvr6N['�ߟޜ�U)O<�[��(���Ͻ���BS�o^�}H��;���qF�������R����K�U'R����G��:��<���8ː�Y'{�G�`yy�o>���:+�&꽗�vWvrjR����~�uBw⚜�x�>��)�ݡ�����ԥ)�kX}A�WMݤ���r]a�A��]e�u�BW�����_�BR}翷�N�hK�}����Oǘj}�\�Hu)O���f~�f�s��s��-8%)I׾3��'�r[$�g�y-�v�Д�U�1�.1ݗnЀ�����SR��^O����R�����>�}U���k��T�t��E�e�9B�ie��c+4��^rR�y����)I���{�'R�'�澷��JRyߟo�:���>��V�������淚����;��Iԥ)߾��%)I߾k߰z��/��~�U�T�Z{YLM�WXW�0�yW�N�hN�ѯ��5]O~�����%/ �ϵϬR�����>��J=�g����%;�3;ݞ�N�s^B���}��R���������~��=K-��y�<����,��Gki�[3ڸ�ږeA�ڍ(l�F�����&ik4K���e�L��M�%Tq�*%�8�� w�#�8S�Ϡ}��D��5�vp�k��J�۬�u�4K�:�xu�ӻM����:���a�"*�iIQ�����o��
���%!.����r��.�����7��w{������z��nV�7]G�qmK�[�1�MN������'r��A����┥'���߬���/?>�V��ӲCw��N����
r��R`�@���7g!y�o'W�{�Ǩ9.J}揾�:����~��JR��{���k1��>�}�͜:�z�7�{�f�������w���);��}�'P4%���~�5A�y��؝JSy�g�Z����kY�\�g�);����ԥ)�����`2�g��؝JR��ѯ�`����ߋG����u&k��fovgF�S�){�o�Ҕ�w��>��JS�=���������}�W�^��eөRK��5.(�FN)�<�#߱:��4swY���n�n�6��zw�ĎM�&Q�[�q��5��Д�'�y������Ϸ��S >��=�3F�6p�Mu�_I��ߊ|)	�)͊���h;x4=a�Ss��s����N��8Wv���>o.\�PqźuU��&���[c��sP����b:X���9	�ͥgx�)eٰK��_��L~�������P4����R��w�0JR����g��	A羿���k|޹\5���|s������pz��/}�{�	�JO<�#߰:��;�^�}A�W{�ʴ����>�v��5�RuJw����-9)I߹�}��	��=��j�S$�ϴs��)�~����e4���ӣ�g%�䷓���K�%)߾�f)BRw���N��7&��.~�5��R��߷��G5���Nu�]u�4o�ԥ)ߺ�k������z݂���W[1��6u�P����>�g�NO��Jy��>�A����hz������įd��[س�@��h���icX6jVm���o9-����~���J_y��9	I�{��:��;��5*����������V]�)�J��:��o����E�#��m�'ﳨ���)Ok���2R��}��W9-翿�u��gln�[{9�������)O�־�Z����=����z��/=�~��j�Ͻ���:���.drL�	�����
���]Q����_}�ԥ)}����Ւy�y���%=秺�n�l͜z�-pٛ��BRu߾��:���]��M(�V�Җ�iQq�MH��*TT�H$���_}H���8�V���*�޿j�����4��t����������J�V�)n.� h�]�<�䷜�����r7���~���qz��<���qJ��|���J[�O��	��ݽ�ݜ�������=_� |�_[�)�������'P4'~}��`�!���e���������îfq:��;ϵ��Д'}���:�־DXsF�/=���@���>�g��)Oy��g�,��9��vr�F��)I�h���)K�>�|R�����>��JS�u�0����Z�c���RfJ�:r�����%;�߸qJ�
:7�Z�fu��-]v�.T�깻[%8�5�z�3V��'��}��JS��_}�	KA_s��U}�}A�{�m�qH]U'�σ�� 0�/cxx7����k\SP��y���:��>�����(=�_}�ԥ){���R����o�Vkeé:�7p�9��ԥ	ߺ���~�R�������JGϾ����'^���؝BS�zz}��ٙ��������y	I�h���hK�3^��j����Cԥ)�}ÊRw�m�����ˎ��#�.�
�����׿`��d'�y����JS�5�2� e��e�$� A��D(��!��z��u�Z�Yfa;�Z�ov�jz�\�*�n��4�©K-�Hʦ��ƶe��=Y*�/l�o=�N���s��W+�T�{v�x��g��Y^���6�-�jx4�6D��ʲMЖ���zt/f.��i	�1�ג�W�#qƙ��Jjrp>�?zV�Xs��{���jۦ������v�d�^���}}�P��r³�:�F��la�;)qa��)ލh��8��־��%'�y�������=��jC�+�t_n3g�޹����;�[Btr:YTlNrn���ԥ)����4%)I�����N�)K�3��)<��{}'P4^y���mo�kZ�l���MJRu߾���iN���R������>��JS���U}L��}G�:�d���y�����=JR�~f��ԥ'�����:���F�5�}�	JR{ߺ���)��u��	%�Q"wv�]FK��}A�w�׷�u&��N�׷�S h;��w��JR�����	H{��}�Zt��u&�������BR��׿pBQ�Pg�󗲖^'�R�-D�S3rʓj:�vY�W�|������N[����`������=��J}��뙽�V��g��lsVg^�~�m�)�kQ��6����-��� ��XB�0�5����$�W
�b@� `�$1�!�	`jO`� ît���!,�11�$4���I�pp�0 $�������,����:�7�6��10c�(���PLF��s�7G������
���>k�RE��2$u87R�HTe����S�
Cˮf�|*��H$�Ar����9��fF�&�k�Ĵ�<!����[%��tƵ�<ލ�N`�Du��30E!CQI�6��"�
X)�
�`� $�jJL
$��'$%��c��ԆKdXd4��T�ւrh�E�<�ItN�&����dR�ad5�4�r]a�w�F��Y�e�ف4�Av���J�C,λ6����:�s{��3�o(M��	Lݮ�4���AXJ���Mu�#ؙ#l���kQ�F%�8m�J�u��DB���5�6I���s[�=�����_~�UZ�5Uz��Kk׊���h6�7n
�[:��9�"�Pm-J�U*�A*�U+n��<��~��j�x�N���Ok\\����¯�2����!��k{��ñu'�I6����oLu�eܜoV�.�Y+��B�y��p�}�Sے ������f�t-*�^�e�kzZ)��Jv�����yܨk�`B�.��Ġ�Vc-�G$X��(�շn'Z��}��w؈9�\��&��+ѽ���ʴ�J�;�U�2c]�э\���T� ���u�P{9�L:���a��bX�
�3@v�Ÿ�5b��qlبj��p8N�b��;f�Sb���@[�7ED������ږ�6�3m�M�����Nrrx��>~�Wb�hN?����&�T:�-kZ�eaf�-�{5��Nb����ݮ���{�:������6څM��v�M)+6�)nI�@e�7LL��-�&iζW��%�WǏ''9��	�ncv�X�:��r���5�Yk[�l��)I��{��JR����`�����=���)Jw�Z�쯩�Us���j"�«2d�<��u)@��o�%)I�y���=BR�YI��EDp��t��">5*�\VQӲA�w�=�&�r�=�}��9<�R�}�}�BR�����R���ݺ��U\�U�/�*�1�;�N¹'P7;�bf�׿oBR�����>��JS�=���):�<����Wh��7�+�.˫���A���������V�'�;�p�8�ɡ/1
_ST�P!�*4���M�}=�ú�U�w�����3�l@�F�U����WJ�YP"W]����{�P=�c�gS��V�(mI.&�⌥wv�M�H�5�u�}G�@�A�`9�f��b��fDO�0A��FT�V`���A'i�Io}���Ir��S��y�w2����S���$	�yA��c�h���*T�r%,T��z���yku�5SI�DT8�����)��+nL��{���M
t�t<��n�Nf��5��t���]J�����l�I�y&��̓��sۺ�'y�/��;��Y����9|��`$���:�`������]���NѼ[����t)1���dVNp�ǒG�o]���w�.։����(��rP˔2X����{�{�5�{�ʝ�E��ܢ�z_w{8{j��vު�Ѱ�0o2C)�)���G�C���W �*c�A����o�6S��YvZ�Ӑ����n�{� 5�\PU�H,�ix�)�$��S�8+�w������`��,=��6���eǊ�F*��"�. B��k�_~�jyAλO��W>��s�h�C�n$���X��	`w�=���^�a�>�^��iwt�!2��r
<�p M;�{����G�2��w'u�s��S�mIV��}@�Q%+G꯾)s_�/؃������6{q���Iq�6�Tk �-yg��2�%��`}��k�[��+�-�[WL��.[Uuۦ�MOY�fEW#2��eti4�B�)c�v�n�J�������4Z�~
J鍆|iE\��h���-۶vXh�r�[Gl�m�[��+1�$�ϒI_Uz�߿7��[��6��cYm��L��������q2:iT#�BR}>m�Ia�3��ǆ�]����$��{ u�x;���#�2�
yS��Mk�$�/*0�#yrA�7Aδ��;���Hrz�9���M��7����&[�w�C0�����ܭn�u[0Z��~���軻�������� wm�to+�*�^�s�w�+���<�a)��Lq])FU�Y��>��߽8^�{��O(�">�WkS�(��i#J\N�ժ�X�}{�����#mҼ���j8p�Q��*'J�Lb��_��w��`sݚn ���s���dF]�����+�N��;7�8�f�[��lʶfk�bb�F� `�s/.���u��	Ǵv��Y:�s�dhScs��Q��Ù��{n2�k���I�Aѣ�R�"?
��;t�I$���~���\�<���G#ﾐƽ��h�{�L���d�Wv�$w�}��+��+�ݺ�;����l���fƮ�m̻w��9��:½�o���}���ȋ ��(O���6W���P���W5sd�}�Tf�sR�?�X[>����uQ~�>��W���}��P(?�B=��G+�}�*�|(���
�2��=�{h]�t�N���d^0[C.F��?�
A���i����v�sݞ�f���ܦ[wi�7�4���[��Y��\A_����u֭��0�)z}����'�D)5�ϣ�����}U\ �忭�^���)NV[������w[����}���}�X�<�$��Hs�}��_�G�	*�����ͻٳg5�����^Y�����P-V�?}}ڈ��DG�EԯO�r�:�~�cT�8�����M@fuw<�\��	R��/#��"{���
]�F��ڔGd�c-9N�s��ӼAu1`�9N��J����)�72��`a�������d����O�C���(7U�\�.&p*�e�A�U��(*THq�C��Np:���O��[Ͼ��}�@պ��3��ԏͥ);nA�(d���O���">���>�MײC�<��6R��s�U���S���u+*��`W{饁������f �@�H'W�h��5�o����)�H�R��܌VϾ�������|E~�z}����F��O�~������]�~���Y.@i��b0�~����z�Vۇ�8�5�n{Cn���F���h7b>�w~������wǽ������Rw���rZ���e�gx[��.��CEӫ��~T'|�:7�7^}�ߺ��>w�R��n�fd�d���n��s\�Vk�u�]��o���@ H���~�q�e}��5ʼ�߹�X���W���8��e9(�$�h���0��򓨥t�9`=n�9��P�nf��\�k9�o]nκ�@? ʤ��s�ʽ��ߺ꯳�﹪�+1Q�9,A3QYW9�����o[���;��{m�9P�
�W�A"b&�D�t`	�	��VݰTl�����NC��ׄ)\cK�)l��W!6x�8�'����x�f畊�m��Y'��WȺ�)<M�mqCs��wgus�l,e�0�E�Ьqd����z��U}�n��_�_�K�ߚ���������{���.�(�"�#�<]s��6���$p���&�y�CwRl�n��CyCp8QAL(�/|�s͹l��S�&`�S��>���g&k�}�O׀9JS�@wU�>��� �?s���M�vT]�N����A�Ր����oՀw_�ܐZ�~	�(��~����l�F��Z�wF˜90�Q��;�����w�)jS�owQ�)v������������?s�9C�Poud3�}�DG���~��i��ܣ%əW*䙔�m��#�HBY�m�@L��2�R���8*��os��0-=�ÝV�*IU2๹.2�1/�舂">(�U��p��F,��#T���ŕ2h"��$�dd��!Ea	P+�������al��WV݇F���e�Y�]ޝ��a)���F㯻1!�C�@�O1�ݒ�ֹ������ e).#y��uǞ�3�a��mf� m�X�4t��_g9�O�2NL�ǔ�r���<���|�e�7V�=6;c-���ZyVۻ�����"��}�X5�߹�<�q�2��k|�W�_Q��5���[-4\�3��|��j^H)i;�j���d�
���u�o��뙝u@��DBG����\�����~��U��k�������	YU`�%I_��~�u�?2�j�`�B���l�%���W�9S�>�\�&���UZ�X�4R$�h��*nH�}����`f�n��ym��]�����}T�<D�Ir5�oF��v�ٮ
	�@eT����!T�$k}uj�{����;�d���|�s���}!�v�rOG���[Nv
GE��o�37�Uj� ,�
�2kC
�C4�f� �5�a,@%�#D *f���V�c�I� �$�D � C�WEN������ ,QS� B�#)��w��d_g߳��w��=���/�VQ I  �H�/��s��?|�K�O0�٘[���ν��?�UW���z�=����Q�7UC��n�'g.f�f��E?�!B���ew^3ܐ��l��]i���"#�i�z���ߨ��Lyv�1)f�w]��s^�F�[��K	���NN�vb��-)�	�#���'�9/'9/>�"u�ޠ����Ki���!�\R?M!����8�����$��Ǝsf�0����种��U�~���#C����0�m�z�U�ɚ�7�:�|�g��:����~��^���秷ǻ�i)�9E�v����[[�ـs�4�U]:����`���&Ă�:4� BbF0���F�#1,�h3o4	�E�H���m�&��z$���N���Zd#]q:�rx�w�̰���;����Lv�0���Jvx8��&�5�4�D���9�1�D�Ħh�~����t=�cX��}�/�����_}�06i��c��1�`c �]������%͹\�a�=�W#Qiˉ�؞n��u�XG<�D����Gf��c�Ɍ 1�c91�c5�kZkZ�kZ���Lc�0+�6�S*&-kZۉ��kZzJz�Ơ�Sst����մ��4�YXv��\�v�]���0իU�r�)����iEf�65�V���y�i�Ӷn`ڬr�hv-����a%0Z�&�2��dɗn�l�m�Ѹ�Ƭ��`�4r�M��7P���&܉�ͻ7iZ"�9ѣ�A���Vғ�`N�c��u�b`��� t-�,�^6Ɓ����k:��a3�m�6�갛0��l
��P���X��l�%�q=^������R9݇';\��n�U���:P �oҁ�'�+ʋ,�WV-��I�a5�r�����79��\g:6اHO!v�&��Y"-�����.��p�֜&�:����ځU�c*���Zᶦu�H��.P&64Ż�ba�c��
X�s�\�u�)O���/=&��U��[%��a���|��n�t/.Dp��a�)� �ܜ�b�C�5��iֶ�������^��m����m�Jr�M�.�>b�V��ˏd��)Ю�j�of��k,�����Q��t�;��nR�f�Zٜ��J#��G�a�N�iDO;TCJv�و�C %G�uV��A�7���Z�gy����Y���0NQX�<Tٌ�-b?�W�-����� �[0>���ʭs��h�9���]����Qp9�{s ��U�"���h���rnv��E)BRT�ӂ�=��;�qq.��v��jF@rd��2�Z����48�j	�I"N�v�-��}��;ֱ�%l�D}�}Ϣ?�>����w��(���'!r���JJE�\��̈�Ѽ��m�l�/0�>���DY��C�J��x�Yn�x������f�0��v�G9�^��%�QM�R咜e�G�@���(7U� ���D}�/��s������~]�0��t��%��.,���A���cL][��w�=F���Чl�Ҧhw���Dۚݰ��e��Xک�s�D���=��6)�t�f�UC+m#���;&ni�gq���E�RMK�d��̼B��9�����NI�H�O�Ϸ�zߟe�?q��N{�eZĜs��|��B�i�I�溑5f:�e�d#�f��e�⟈���k�������r�w�{��nꍥ�KJ�>� t;�Q�R���
[n[��/99��t�]�:���l�v�/�i���Ok%��<v��&̠��n�}��Ü�0�ym�Ż縏wڈ�iK�r����qK�������g�U��+��swo�V��ņ�w�S�J�s2�(˩E󀶛��\����>�>�A��}T���ف[��?%D��u�D��ž��GNb+8�����i�Ql���fR9�[0_>{� ��>H9Ѽ�k������d9$��r�s�|�n��bb�ȭYXy�\A���s�`��	�DҸ��@R[D�������b_�ݘ�gn�W40m���(�2�D��f�t���,�{/w. �l6�Ŗ��F����Ao�kZ�/�_Ͼ�Õyߛmv�j�7�:���(�W6YU�9Q�ќݜ�^y����*����W/}��*�?~�_���>�>����"�����>�"|(e��U����o���ݚn*
�}�V�w�m��R�v�Kd���5 ��(�A��)@�g|�|�=��i�Ry
4m�]I<��㺰�VdK�}��U�t|rWs���rF�ػQ(a�F�k2��	�� ��@d`�!Q~���~��{W�A�zx�F֛�����}��P��-)[B� �L�����̧*��w��j������y����!#( �
u~ϯ߸������?:ȌV��YN�x�����]}R�����D�]Y��>��Wy��2��Ͼ��	�eRH�}W����k7�o7��Z�����������d�����W���(7]~�l�]��l��՘����m~��@�A�P����z��~���Z�=�T׸���;�R�)1�N*V�������>���U�s��$�85��ش!�wnk��I�S��uϿG�4�O�ֽ�8��0��������m�nk�+Y*a���NҰ��#1%�:ݶ;�m��ۯ�e}_}H=�f��wt?�mJW.�N�n�p�i�PvtO(7u�p):��QU_U*9����L�U���;Vb��� [����v"㏜UQ�e ����p���9HNY%+��K
�|}U����v��׆ q�y�;,o"����]̧&G/1�����A���`+���Q5��ɚbb]�nŖ�$�������G��>�j�ǶC}��-�0;���8�cu�<��ԂJ�QB�b�q�;�d�����<m�Su��'u�s}7l��A��RJ�ǘ�G�� ��v�w��� ��k�;�m�⯊�ߍ"���r�dW�u>p�Cy[2v���P9M�pl{��E9���4[���}]������
��v����\��c��*J�J��o
���*�oVH)�hن����m-i��80�>9�W;��E�:��h,�%:��sZ���,��rp��\�G��>��U.8t&S�$e��[=�4]��l��mhM�t���	�-�)4]7MrNNrV��_������o�F�!-+�\%4�w}u���xW2� ��"�*%(W3uݗ�(�`λHO�З����8UCyCݑ�.���ŞI��f��0���˵-ŖJ��p>r���Z|��ԭ������=�j�9�d\����l��):����!U�#�}
�·�jVK�N�jTd�i���8��ی5{�ms�=���|�=Q�R�\��t�d����S��i�@Aλo�R��o�zlv�[s�I�D��饖��`�,��B�e殶�e��w�)cn�/y���r}�~�����k����ޭ�f��-j:q5+v���r~s���+�(��]��&��i4`�M����;�����3K���is�ŋuͮs~�]�5д�A��D��X���yŻI�t��0nJ,��H��CiP�Q�JC���vnaA֭���9�">�}��DvCg��fL�Q��)B�`�
�E�����L7���]u�?y���W�����B�%Y%J>�{��_�6Ԩ+��#V��~���九Տ�;*ف��ܕr]�u��Z�7��zٮ�����F@�I�[��?��p����:�^y�}��?���y����,&�*j�p*�������>T*����
�(�rc��lK���׻��TbfQd���~Ϊ�=�?~�U�{�{��~�޵����=j�1�eA�)��LJ۟FD�"�0{�K ��}֫�����!
2�J�����?��/ʗ�i),�(:N�VÛ߹��jd
%$���x+Ó���NzU78s�*\�A7|�0X4L���嶃���0�W�}U���� Ȑ�	n�~��*������֯�=2Z�&;��2�5NX͛�ë���w��}��J��!/�������p�����Ħ	�VB�`sηm��vQI$��.uHXb&�,��Zr0C���j�[h9���}���`7^�%%%�{�T%�-cw�V�W, I�����q�]����r�N��:�� �Ѽ��5�(&�EW��'f;P�{�u}_W�H����c�߭�w�z`p�j8�RZ��m���wߟs��_y��9/H)	�V) -�aD@C�!I�acQDx��W�V}_S����?.����o��┤���2*���p����s�:�� k�w���$����IĤ���9�]�����咹:i�Z]�h��lF�KRtC����~����Pw��� ���Xg�|�iD�b��O�<s��%��RJ��ّ�G�s�\�9cyI�G �Ѽ�������տ:{�R���#QB��vn�?��p�Psu�8�-�G�'���31W�;��)�̠�wn��M�QZ�ݶ������%Hˋ[�.�y�D}DDJ�S�r�|�� ��|�G">�^Y�K�{� �떖&�a�&+PK��K���κ�X���ٵ�|㴦�W&���]r����5�B�T������/(\�\cw=C��(�&�b$V��ڸ�F��V�6�gB��]f�B�\o<mۢ\v��]r�LIN?��������:o�v�Y�^�R�4�����v� �V����Q�w�y��s��y����Z���E:uR�}U]�퟽t����X����j�9嫸����}#��R�����6TMIR;�����[�.g��[�@n�f���.���eL���	�Z{o������9���"�����R��,������]�<�L�/$��8�|�l�O/�����nf"��Zc�?}��.����^^�8��#㛶��D�M�\�WjЉWW@s�������}�̥��XKo�d�I����J��$�53173�ޏ ��s��/$}���*cʾ{&�	�Y��@��r"A P�I�j	�/R��X�! ��
�U	,��A�$��&2�@$��e]�d�"T��SA�		���w��άú:��opJ�u,�Ut�71ts�m�'�:5N�����,ueV�X��j�­]T�n�6�uA<�ub��]5[���-�J%#�y��a��Q&kf��[n�$Ӝ5cfm�klM2��0�3D�%Mv#s��g<����s맍�zƁ�9m�j&�u0Φt�'˵��X�UOBYر%�yp�� c�I9��c[x:�=�ۮ���u�ծueaɑ%%�7TiX;bH,�vo.Hy�Ec��3�Z�̐�0m�RY�l^�0��9�3���K*��u����:)��jAc�fێ��j��*���γU���{l�ʾo&;i}Z�L��b�R��J�kj���3ַ@�v�ke��7���f�� �E�5�� %��:�{E4���QUNk���s�f6�6�޸�Bچ�2hR��n��6�z���grv�j�?=��e����lx�5��6�m��Q������v��.2���z�r)	J�l$m��ߞ�/߿����O�����}A���p58��T9Pw+�#�c]�oM�;�;��(5�������3�=r]���d���.�ޟd�5�|��Z����ی��P����+G�_�~� S��(7�l|�7[��tS���Q㶦D�fw�ug��1U�O*!'��1ֺ�=D���]&�D*A%�����5n��훸����0v����֠�,� �(Wv;���-����Ҷ�o���V��fj��Z�4)�̪�cDÕ���<����!��!�f,)&(��1�r<�##PҀ�D/�m
a*�HIS4I`�&de�(��L�IABY(9�8d��	�/{P��~�y֫�=�X͛�O{��;j帤���8���r)V���O9a��IԦ���LJ�dU��������V��;���V���$���m�9�3�7V���dD���ATSj�v:��O�r��r�����|�S�yC�)ԕW�;�>Z�ٜ@+��F\�W1y�7U��kWd�s�wvٸ��@FJ��ݥm��a�wۘ�`�!�P9��k�Nf����'2�A���˦���}��V���UJ4%�!��0�@J"BM ˂�3����W����޲������o�6�RK�-'�%a�����~M�q]���9��u�p�V���:�����$�\�05wu�7�,���BuŬ��E���qBR�J�U���������a�}�xZ�6Է.Z�(#�CY��� �K�\�o��~����2d��c8 ���7���3UƝ�9`練8���]�vn�n>�ߍ�Њ2@�j	]��w�����n����6�ܐ����hH�qp����
�Lx��[�Ü���;�oom󓜞�<� �g;`���2C	���*I\B]m��н�� qucSՓVB'v�.wZxĒ+�`k��k�ûm:u�Ckg���3�eS���nM3�"�{e��sUÓӺ\�m������1Ԋ�1�Qɪ�ۮ����iRmO�d�Wֻ��W���������2]�+�%7`s�=��3-� Y�̴&2%Wb���e#"T�j�&�Λ�Ü�����k��H6�d�y���ܢ跔�bN��Q�l�LP�W�$9�����r��|��7e��Z����ݗ5G>c;�
�A޽/q�]=��7}��ytݶn���iKML&@�yV�Y����.�OR�����ֱ���֣d�V�D��[>���ww�ی��7�:7�$�@�
���DMXf�ݷ䲯
RH���TJ���W<u�G��$�oWP����Ic���ff��\�����uπ
�d!
IdX �$Nr�yխZ޷��X��f�<b�.絊�o��Ik���m�����CPJ���Ƽ�@uB,��fōa�=C=�y����ڨ�E���(�0�'9<�<+e�ML�i �c4���wW%�$O<p�O$7�m�������V���~�M5�e�$YRD�WF�S� [P�Pk�'�5�ueM����V&<�E����qwҶ�}�����~07^�7A(�h�
�l�
3#��#2d�kE�Pvto(�:�O��F�]7���ۥt����w_�n>���?��&Ӎ���":xm�GaJ$)��MÝ���9��n0��J�Fqwi���19X�U*} TT�a(!@�R��y��=7yAԞF���Pľ�R]eNT��fk����ߺ�E{~�G���\�,�����m�3�T/V�a/���s�ڸy!�,g*UH�;�7u��7�ZJ��Җ��]I�9��׀)�<��O�\����M�Q5w3S����c���}+m�X$�oD����wc7m5��I�p\�M��{�`jW$5%��'F��st��W��[q$8��ʢ�!�Q7�;���s��X��k�5tݶo7����d�'��c.���ns�}G�2'L��@���Hou>p<o��BJ�[���%Wa������9�bf�}�}�Ls3$5�fL�C�Q)X�3K���%�~���~~?~��[�(�s���"_���(a��z�rӸ4Z����fR�J*2��uţvvL���55U5d��=�M�jO!�@I;����3�oo�v��]Y`Rȶ�AQ�H:p�{�K5���5t����n3��l	K�һ%Fݩ�]!�z>����{$��p�	��R7jR�2��E�t��/{]���^�wf�q���Ӻ�D��r��"��`oz��s���ī��nc��~~T�Of��Mg��ж�����0�4��$&x�s���Md��:q� k��؉ή��)���8��N�T���0���D{H	%��S���Hcl���#6wk�]������%�sZ��x�Rn��)�Ϩ������[v�V��hE��*+�������D�:*U>n�7'/W���c[n۳U7?�7v܃���0u��$��7����r�Z�&���E:M%$ ]��rx��.�9��������h�O�5�L�#*�Tl�������|�[I�����${;B�\�j�j�Eh;�����i`g_�n0��k�#}�Xj'Æ52�I/�\�)�/$5Rn��y!ݴ�G7�*M��N�pJ�FՁ����ry�Gm�+*Z!�3W.'�Pt�$�����i�o;���٥�4�x�r�0YrƢEJu�
`bgk�\R[�ޱ4�LR��v��A`X�`7#*S&�l���v}�qC����IL��)�aX��[��wx��9���@��Q�I�9Q��������On0���ڰ9��pjP�Z�M��'$:��羏�/*R�zp�{�J�gW��[
lj}��4'aY�H�٥��Z'�t��Ƕ�(������*�#����h;͞Չ#����秷{�ڬ3��C�I�b����J�]�a�~���y�N������/,���x�)R�)�T�H'@9K9���=ݚX��یӿ���iX�|���UlZ�����h��j/{o�m>PU<�+nӞ�I�:�	q���]��%d��m������}�ɝV��[�`ݴ�_}&�d��J[�IT��2��_�n0��l3{��%�綎��C���y�x[�3���"&>����rfE���P)�<��]n����#%F��q\i���v~����%��Gj�v��k�� �I@qF�
�"�}�4��ی5t��7�z���j��ڷdI-҄%�R�d�o''6z=�� Z���Z$7i9���V'��z�)J�+(�Y ��g��� ��i�3��O�Aݤ�"#�HN����rs�8���v�3W�m���0��Wj�U|?TG<?؞�DHd���d��2���2� �d�N$DRQ1HR4�d����C� ��B�ة����k�#h�2�(IGR���5-)X�c�`hR�A��G��1���"��Y�)d�eHIP���i%F%j,�Zĉl�V*)F"�#%D�S�!����D$���P�%���$%������?����N�Ÿ���nh�ֵ�k��X'"�����^�thL^GPV���m��<(�E۵�ny�pU�:���R�3��Zִ֙�:ֵ�s:ֵ�km�gZַZְZժ�c��b��ЮZc@Lc�101�chK���M�6h\�4�Nؚp����KJ��ݛL/�Ɨ��ݙ��[D�ŗ�����Lݥ3��h\��ԛ�01�K�Wix�n�o	h�ԡ<����{$��G`G*��;�Τx�ۚǭQ��-�y�:���k�\X�۫�:کQ�Λn2݇M;GVaӪ�7����l�kl��;np&m�F��b��Q���	��u5�b�ks�L7@�b�Ss���]5c������&�TG��X٥ܺ:lr�KeXB�\���+����k�QU$
��)��r��n���Q��c	�]#rے3l�l+&Hu�m�u�kZ�`��ᨘ��5� &2%�)�j�� �k��!��5�����4�e%U��IY���s���TѸLc`��F+ix�U��;l�����4%c�����XP ����(+4��r<���vݛp���l��+i5���ڃ�燪琑r�Nv�2�H�h2mfіan�JMAAҼ�A�`j@��1Y���R=k�ۭ����͜Ƌ�\Z�m�;�	d������<T^�G�8"�؋��������/Z�TE��ך�^s-g�y�7�Լ=����9N��=���N��V�g ��5U��P骘��l�v,��_�XAP�>�;cv-2��K�	���B�馅���a�M�a��n`sO��n4ͻ���a�1d����vѦ�O�CI�J��w�<n ޽�`s����˧�ٞ�v�$���	d��p��0ݴ�AݨO(;���GMoTI�7-݉Er�Û�n`��¨��񸃫�[h�m�G+#��wug8����$:��W�}s���{��)eA�%�%�fGC*�8���+:Ѧq�;�L�������ݹ:�n{;)<n2�g�[`����ð�H�Pj�%�:c�����ݰ�8�;!0�6"Ӻfa(q�s���X����gJ���P��Q���s���9$��~����ޭ��H�R�(vÝ{�x��&���ԛJ�2��D���_IQ4U�jS��i�jy���jo:w��Δ'{��
��c�H$�*Gkuw�m��s ��,s�ڰ7��YJ\Rۧm)A�(��g?_�j����N����R�M-����R���j�&S�{�u`g�p�+�2�3� �����L����+.�&0������Nxi����|����sM<�iʌ�f;�D���_����99�N|��:��AX�D�f�u �-��`�R7]n4�M�v�Ry
z�C�(��ʛ����ow�(23�2@@M�n�,�ʭ[]u���2M��з��,-��fswͮ�����m�����.�,�`M4pta��n�hȞ�>�m�b9�;P���N]��]����{1�$�N|�
k�\pvH퇷���uw���g ԞFz�qeQSrs9S�|�p;:'��m:��'�է�_UV��{RW.
��Voe7��C���8)�������4:�.L�Z��^�{n�sg�qt��+꣞{�x{�u(Ҳ]Л�RH���0�S|�����UM4��\B���d�L���u :��~���^'=���TS���]_y|�>�{��`1Ɂݹ��� f�X�g ԭ���>�DD��߿f��_�u��bWWRG=�}���y��A�!�������k �w�r�ej�`j�7D�Yg2���VM�p���X�(�ﾕ.��`����۠��)wn+�7��Kz����{�Aշ����r:��b�1��2Ӻ�0=�M,�%)SL��i���6T]�σ�:;#�127)A]W�Y���:�{m�;ݿ|/璘�8���t؍��Vb�Q
�*M(�r
X�m�{U� [����G�Ds�(~�=�<�=W3+̡[�����~�U}������f�{�u`t6���������۰���|ˑΧX{G���&��}���ͮ���SU1�iQt� ���#��yA׷	򊞻Np9#��:��Jq��wvJ�X��Հ];1����v2\����|�k��蒪�E@u9�נg;=��W}�Û^U�:J���?W�����e�a󂑨ܒSlϫ�-����nߌ�O�������7�:9sS4슫ɬ��.���>p�l�8�ެ���U|���Ѓr�[ǎeB�<���y@���pճ	�[��(��m	���d�J;�5`s�������A��b"�ޏ�jəUe�L����m�Y�����8I�`3������l�t�pL�(�m�la��*�iH���d�	���v�%S�n|����{V���&�nf�#�P��R����f90e:��4��Ä�gvSdx���:��,d�󜌜�/�?�-��:�Z�ƥe����](���k�3�}z�`8�%]ˈ�5(
��t���h���:��`n�m���+��ki�wa)Ti%Q�?�_G��RT2
���o�?~���`ݸo���}�=*i��o�'���Iq�UQ������3���0��������UE�iB��PP��2 z��pT�#��W��>~��"�iDJ�̬�.�����5��A��w0�f�g���gt��8�J]�c�v9�wʼ�r������)�-���Fӡ��3��=S���D�[o��V̩���8�����ý����������j�Y\�86̖Yu3I�=z�Y�p�d�whz�*p윗�%�Gm.�@��a,׵��٧!�V&� l�n���7�v�N�4��@Y����U7e��T��{p�(:�&��jT�R$VK��lP�3ޕ��8��v9�wqtݶ{�{�Զ��e�R�R�p��ə5�������R��=񺣡�N��'q&Z?}�WԿ{�����F3Į��7�kDʁ���$JX9&`]7m�Ֆ+T��V�� B�m�	nhY��q3PT^wv��4�0���	�f�3z���GMe��c�.QE*�&�ԑ̰��w)bk�5��ȐI<���
��8]�#�\ds]u_g��r�y�����xt�W�ߺ\����ݶ瀆��qu7�979ww8@5��(6P�Pwu�G �;h���5�E%&[�]�t�諾�m� ��C�ԧ�)s��]K����-8�$��J�;��\��|�0��x�1o7Wmb,��e�.�f���9`n���'�q!�YsM<;�΃��f�P%]1�@Q2���F��]`�����׸�Ry�}G��{#ܓAĿ�XUL�Me����`6�9�췔ݸo�i5a��֭R�S���$,����w����՞�ӤL�E�R@ix#ռ���������u���[Jq��.Йu
�7��[�w�m�ws =��a��%[Z�%#ĦSLş,��]{m�諭�lÔ ���x��$���㎶kI5��T�\���~t�7�Rwu�GG.Jwkt��Nrv233�cv)���]LQ6Ae]�d�$�ܐԞF ���� 7u�a��un�M��o9���-n���}�ɺ�=�P6�=��|�W:��M�YV8!(���;ٺ�(��u����x�A�<�!�u7S�3q�nf&K%^պ���w�������v�anvbj�X�kmAj.�	A�e���x_75vV�ێ.�*Xʣ�i���ɴ�e�v�L�*=�����X��ۡ�dt;:OLM�:�6��b��tY��-�Ʃ���<�����v՛a#T� ꪾ������v����WI��-�}��]fccBJ�ӎ%VZ�%��5 Ě\������]bn���vu��Q��E����5-9��:i�M���6�N�����{w�Ձ��L �׶�����sۮ�q���W)���"�9�C|�I\<�oS� R��,�EC�T��I�� ^���`s���a�쭴��遽=�2�*��v(I"��m�Z���!�Q��W$�F��>���j@y�j�����3�yό�\F���bm�m$Ңe4��o��]ԃvl� ����2��嬐�H��mWk+���?8���"j�z!َ!o'K��Ll$`^��n��0��(�!!�H�!0�9�I�2= h��ӈF���#ăBl�sA7ѣk�&	�_g;�<����o�Qb��V��Qb�/F��g[gl�bΎ��aފ���kT�k��L�j�/&*U��mWU+v�[���*1��lj���z�J�0��*K��;LS]���;m�v�i; ��.�ln�i��@˱`Ì]*;�;[:͎�
���ƥ�a�e�2:YF��Ac]C@f2����N2c���l	h9�!����(�ڙ� YF[r��`��(�!�6-��LU3���lE YZL�V-��72 �c��n�K˶7X��̶�S�.��E�	���Km ��KB0��ڽU���'=���6x�F���V*v�['�J�3��1���F$v��Y��
�q��s��XG�AꦑA�70Þ��3��߿���ߨ#`!�	��}6 #������m����!vظ]c�a�s�9ĭۂ��	�gOEv����a�i�������n�ue��Z��#��USխ�;$KX���ܚi�A���߹��w�w�y��G��ۛXM�[�21nA�7�8ηX���"��8��q;���Z�+��3����h�wS� �� {����rˊ��2�f&r�jg(;�o�u[0��$�u���K�l�w�^��35-^&�v������6u��rE�W7eVB��HK{ٺ������q�fa�V1�����H�VO;�۠}���7]��cqU$�`���y�ӥ�W����#X7 1���D�
5wu�͞�a��w�Ր;׿�<?~� �J��-�i]9�����t HJt�8+���)$'pk����o^���e߾�Հջl���ߕ%&&Ը���n�f޻��W2�[���F��[J	J��)$��J�9�MՀwޕ������j�~�a����V+��#Q�/ 9�v�wn&GN/�j����J�O������5�)O{���`�o�F�Ĩad�'q��ņ�/*F.��2B:�n��m�(6to(9�m� J��3��ձ����Ȩ�)%���V5�g :张�����8t�쨼��Y��9W}����{�_}�t�!�|�D�b��f�j�	�H�κ������W����5{�xm
E�e��V|��}�|���ߵ�93�Hy'��螶�������WUS.Z.�*H\s�w^VQ��?A��Oo8�+�ȼ��\�;��`u+��C�tO(�(�l,�~[��Ə�Ҹ΂3uCNI*)"�����>��ΣޚX�z����I�qv������|�z"">�����[�(R�<�i���j�R���őZ��]=���m��>����\����q�r�P�&��E�^e�M�ݘ�X�!�Ly!���yo����M��X�|�a"�a�e�\ڭZ�^�&�Ѻ���魝6�r�gM��@,ز�)u%$�]�!��#TG�N�w&7Ect�6	VV�?���efҎ \�BdDݵ�KV��bɥ��\뺼i�k4s�\)��va�Z3n��7��?���߾�����<{Rt�[x�*+Q���wn�W��/X1g�%v+8Ƈ�ͺn
�QAJ�(�g;���z�m��۹��{U4H�W�%(�򨁦%%�

�g�P�d��J��ճ ]k$����N}�a|�����N�9& s|��g6n�wv���=6nCz{TbJU���u$�\s������ܚ:��9r������;S�y��O09���{}z`w���>���c�(��~����2�!��Vq黌KX �pQ4��Gm�y�;�ƍ��:�$�VL�7e7A������nӗu9wc����_C��!$T�
N�dd�2c��i�7:]�J뷥:����+GE�%9Wm�V��N�e닋pu�)�e�25ef-�f΄�䜓���Kl��px�B���([0E1p[a�z�����Hy!�K!�Doڞ�:J]�j�v$X��� �vi`qSn� �S��}������eryx�Q<X�[��9��wR^���A�ww2��ZI#cuj�@r�\��!�@�N�4��C���
�2�1̼�U�N�z�������D�m���sX�u��-�Cm�l�o{��[�v��n�<n�E)S�%�v�w�Sd
J��)S�5�&Lf��M������=�^����mi����)1�1��3{�]W~}��f�0�1+�	?J@L3f���L�J���a"j�C�)`��#0�r�sȲIA�	�$�&��-Y.Q����Mb8�ь�b��2��8��a�$��	��:�s 1��;�"�������x�/m���{q�=��DIJ����)K[�[�a��Zķ�w0k�m�;�yk#��QH�yx����V>Hw]�Ov�Nv;l"�&�H�����7q�L,H�1	S$]�LҖ�#�Mp���h�*�St�㯓��Y�s��2�O/w���%�<��jGK����2�t�!w�{���`w��X�3�~������`���Z�-8�*Q`s���=J����C%�s�0j��9+���v;�9�J�A��{qٟR��I �����('���kmKA�vx���z��n��r�V�*I�{�#��Ey��x�_���K(�S��s�����c��ǙD�L����omz����̰[i���9`��m% �j��t����Vw��j�{ٻ��u/!:[��
��u����5����N�}��g�+$I��}vC}�����[�
V;���iHf���H�^�������?%��0c�S$�.UԄWy ����[3�M� �mz��Ѧ��˒P$�� �����u�l<��;eԥc���JH��8�[� YmK$� 
γp���GL"��m�MIm�Vn�p�h��[��6��;f����I�4���qk���嬁�t�YTc"�
 e�W����h
ӊͶ���3��p�Α[GC-�؟q	�'%���Ly������MPˊZT�F��k����wS��l�&�61VZЖX���"@�(�TԉM���P{ݞ�m.y�W��{��+��b��)�qL��yB�a��Ft���߿}�`����:ݳ ��%�.��ʺ%)WrZwRI�=���a��[h3�ڬ	�v�`s�<�EJ�%e��FK����� ��fޫ��k|�F�\�$V[%�9Xqu�[�^���R[�~��V��h�<�lj䃩����2�˾�dI5�&"P�RJ(Ԭy�����j��C[Q��W[{����7�ud`h�J��������
�Δ˜3p�zݤ�D�]\Sb�P !Y��NˊE��.�?�n��2��:aF1=���tk8��5���ۘ�/]��\|uۃ���A
@���A������w[��;�	e �)e�r���\s.��&�r�p)K�m!��uV ���3���I;�WR��5���X�,�km�Pu���Λ
\�tc�X��V)�PoV���ۘD��嶃�}6����E)S�%��BWN)m#y�w*�V4��P܉1���%4�Ж�YQ�v��u��������0��Y"Q��vD���*���&b�,�(�!Lh.v��)��UBY@-��,X���9)��͛���a�3\�s�׺���q����V �<|��o(�։s75%�$�d�G��GwҶ�f�n�n�,u׽l��"�^�Q,v�H��+���|�	'��q+��=�Ys+�ḫ�+�
�,F`w��m�	)�i��.���w=��Ay�7S%�70]�wm[m��uk�f�׳�t�u���S	X�#ck���bu���A�z�{������XwC}C�r<�����:�����@T���џ��"#�z���',�!��E��~��9���f8��z�ge�x]*���嘑��!bXi�ZȖ��f�R�mh�wm�B�f�s�i,���^Ed{,ұ-� �X��C�Cl@8� ����P�Es�Y���l4kV��%GZ7�:�S��	'#�8�����|ߏLc a6p1u�quc�00 Ԕ����g��L�u�hWKu�YY,U���g��v����8��M�9�rEv � �Zֵ�s:�m��kF3��1�3��5�1��gF�T�0��[�m.	�\�1�cT�1�cFf�T����6ڈh)a;]�(�n�a�vD�N��6��������v�\����k�sG	y���E���Q��M14 ��cr��R�.� �֟�7b3�*��Ѩ�R#"͋,(a/L"���:����l]��u�V����T;�ˍ�ĝ"z�O�mf�p���vXՉv�f6:�u���mS� @��ָ��-Ƨ4�[mU�[ l�:�Ƴ�D�0���f@���-����	�kh�\�0����t)�(����]	��T�.8y�K�;E�n�f֢�`�t2[j+5#u㲳���J�6�חO5c�H댦�^�n�u�y��66�f*��3�Ƣ�A��1iPT�6kWe֠�P��gl�d���f�۬^�M�6ε��m�ns`�؛v*�;��q�k�:
��zu���qTcݴ���5�ݙ���;��b��u��NPm�@�[	�iXp-M�Lv�[ͅ2�4��aӷ��.�8u�uN�� ���v:mn��-�u��?��A�Ef���2�ٵ4��|��$�9� �(��#������7�^b�ß��4("�39�y�}׻�͜ �yGccdLI��6�*)�?�weXݕ��(��W�_��sU�K�N�Ī�H �r��秋\Eee!�R�O�M�&����6�����) ��K���ތ���]1�
[w9WRM�+9ﾉ$��{/ǗF7;k�/)A��V]�����@�m�P$�F��x��/P�^�ImKUu$I݆�����٦<�]V��m���9
���Up�&�"����jpl��v��{��MQ"��*�F�X�[��˞^�0�{s01崖8F�R@������z���V\�d���,�u�v���dJ��~�����ε9���uA.�C�;ٍ�TN}���c�@4�gh 0LV�/m�v��A�p�$�v�B`�Z��m�D�2T�(�JSQ�rs��?Z;[F�քx��O#��������j�Sa��9�C�b�6nR',�"H��&{����6X�Pj�S����X恺��S��,��#��)�:i��$���ٻ�7�۫���a��^�s��V���%��NA\�T����">�7]��:���-��2��j�UV+�Gp3��,u+ó+nۮX$���V�.�梢e�%fV��<�n���sx��~�`.�F��jTUL��M���k��-�N���eh�A�\�:����rS�
p��P*I�:{u��ۅ�ԯQS.j��w��G�g�N�v|>;���-�&���,��9�Xt���w�j:�]i��n�%Z�f��ً����ؼPr��7h�O9�ڭ���ceh�1�|�9�K9�Izj{w�pA�.;�K�^S�5gt5����np�����ec��D�0v��S����
�=<[H��W��۹��^�fp�yhGx��2/�O8M�k��R�y!�M�{�P�JNYZEӂ���3��x:�:�H�h���M_.`]�3 9��l%��?�ĕ(�J�vJm��G;����!��!����݅����9*v��5�L���������(C��SZD��8�X]\�d�78�D���Vߣ�>���]�n��ު����V$����s���ݟs`�� �|����{��uA�m��{+֌8���*TK�M4\+ ]�o�����'U<�g�V���q2�+-�*��&���^�����ŷ$<��p��TT;"�&��ʑX�ez�(J�I |ѵ(T�Cq�������-�=<i����*nC�[� Z�I���M[㼝�2y�C.�m�0[��vE�[�u�y�vS��l���/8�',���J�KA�����DD\����W$�K��b���	&K�$�$��i���s����ʪ���$��`wޛ���䓡�*�B�"�.�(�}D�_�S�y!��3���Ժ�~��=Z�~��Хe���eٟ<�����Ky�����H�¬�̘�-x�Dh��𱛈����}��0mBYG:���T�]�M����ct~0������p�髒���~�(6tO(S��G���rC���ѽ����*l�oU�Y�Ż��=ۇ�ݥ�j|��J��XU��Wn����"�κ����{�f%�I������l�p�6����wBr%��svV���ی8�u�z�;KX�R6����G[���ꁣOO�f���:rv7�vD`+�m^ۗpm=���-�.��u.��S���p�n���\q�Mk����͒!�m[nq��mgQ<GS�t2@�<�Y�=�<0�qhK��YG#���d+w���~��1�|�N1)j��;�$r����������*
-8���u`��EJ��r!D�ARM��{v��m��.�����/V��Hq�ǉS�W-�ڜ2��(b�i���yo��O(8���8��K�i�[#���78NNQ7u���0wid�Z����ugWzߵ�r91�R��]06P�PG^��3��yAͤ����US%�M�eFL ڴ�A�Ѽ���ua���y�t��
'R��1ʊR�ň���X��J8)1�myf<�J�l�큕����ߵ�A���l;���{��QH��P���d��R�Ɍ�5�m�@i4��W|��<.Ȇ3����rдs�JtA�c3n��<�ك"Ntr��T����/j;&�֧�ww��x�x��YPZ�\}!u֊�ǰ�����pmj��i�e��鰥�"K#���e`��m�s���A��um#=�^�p�}BR�7,�-�]H��խ�l��PrtO(9��p8�T���Nd��[��]z{m���]X8��g��3�^[DD�c��	�i�o��i���﯐n[3�諳�k���,8e���3�����ѷA��� ��<�R�ꋚ��,��h��n�,9D���mݐ�+��Np�i�e���Y;2����Y.&���������W�}�*7c���>��r0�p�C����(u��
V[���&� ����n����n�ۘ����qTvݒ�IR�wm���m>Pu������~�$��D9xV��AJ���I��F0��p�P���Y5u�ć�tj�mP9i���<�O�a�ek�M��ֳs[.ͪ7�6eU��J�D�n���WOm��{<g؀�|�e{ަ��9��ǒ�G�"�u �rt�1w�m}ٻ����:�v�Eӕ$V.��a���s>�@*��S������ﮊ�ϯ~�=廱[�t�d��d�Ix��e���ʀ�O#?}�GӺ�YRUK����q���������+��\�!Ҡ<��x�d��n��/q�jf$�.��j~��Ѽ��v�d��9g�P�V����@�)kb�(!( �J�0-=��{٥�s���7����n�(r��$T�(�Ӵm�0;��A-��A��������F�����m��{ۘ~��艗>~�%l�[���*Kɻ�3"��6}�9A�v��V�G�^s�8r��U7=sv�[�\ڭQ%x6���Ѻ�`�:��A��ݞ��GI�ٝ�:2��-��ˡ�fu]��=m(Ʀ�+���r�)�������rc��Pl�vW��m��(ѝқ/\�7�E��z�v�ڄ^W^������~�;�ֽU�f\yq�e����`�]9C�Ӣ: J�w�lb���lu�K5p~����Z�z�\�55��(�+��p�p�m�pv;j8�I���7vр쥔��8u�04�շ#���+��x]]<���k�7ݛ�ë���g^��u��N4��p�J����������h�ٞ�Y��Z���Ԭ�M:WO0:�쭴�Y@�j��G�}:�糔%���swTVJ��t:v��ν�`~�-V4ĿD"�u�ֳv��9�S��]�S0QW)7���|�:ۼtJ����]f�։9�w��_GrF�j�i�0�0Y�a���d$nE�,�dVoiNh��l��3e��(��F��+�(J4r�2�BBAڔtm�&��w"@&���`[I�F���0���4%�Y`��C@a�ŃP�KBszVI	0��1����7h�h�H4�lb�٨3Z���0]kq�0,CX! �E����I�9ofr��nL �V�]$��߷]����c�~v�
�*�E���qc �[N���i�\gsu)���f�8Yz�KR�UJ�PJ�UmڠU���(r��jѵ5Z,R���m��q�	���(a�mY���qe�~������:�f�A�nO�\V9vywm������pv��6#�ҫ��1�}�ɵLn��!�j�Җ!��D�Gt��b��s�=s�t+HE��q��WF��
ƒ���جw���wfG�	U��\�9 x��U�f�j`}9�s!�JV��*��61��H���,TT��Rj���ت�� i��@��nθ�۞�k�2���8[����g��#��pXu��Qz4b�Ol]i[� ۟Z�۫R� Z�7)�zD5�R�sk�%w|}y�A�|^ 
?�O��d�O�[�R���)���\�Lb�0��f��Ø��ҿ+�G�d!Q���BA��K�7[jsk(���̱��T�A8J���f�I9�rs���|�屗l[	f&�	N
��ʸ���o(;��8�y!��{����R����ĚV�"v�}�o�R�Psi9��N����*w����I̸�yhrV`����;��,�^���wۘ��u�JR��qՂ�Zv�,�;ԯ ն�(��Q�BuD��V*&�5�������V�>�?6P�+�8����.�x(��&b�b����{߶@���Id`s��᥺v-Ζ[U+�@��)��QE��}��w�4�3���b]k޶{պ-�(R�ݕ�9� �yŔUT7���0ֱ��}��|��]��*;J�v�Jv���u`��+�>���A�V��P�i�L��V,�ө��n�{������8��^�Mx�l��r�L�0��X��� �|�)"�����n�
��ETԐ�%�j���ߟ�֛=�z��9��[3��5�̍���1�TQ:\hXmi3�ƚ�[�>yo��ـs�	e��YA���$T8�˛�������V��,x����IsV�U�W �rK�K�K�������^}����x���=�#�4&�1��:Q^s����U��>�����^E9,m�j)l;��� oW��{����Ի�^��~Z�$�IL�x"����mԗ"�%Qӌ�(g&&v ^��ڔ�6:r��N쬐}�O�jNb����r���l�i�,y��n��<�n��9ڍY@w��VL���s2��V���o�<���YM<f`w��X��n09�����z]Xs�L�(�%�A\�����Z�|�֮O&V����W���ֽr�ƜHN�#� �}����}�W}���e����8��iC["�G<P�@�ږI�6v��k<Tp-γN�����A�u��r��E���ӹ� 3Pd,�����咼�X뷧��b"�1q�%p���Hl�m���n�:�qJ����1J��3��s�DWf����w�E}UN�U�W�~�O߰+�F��QX��+cq�1w��Vُ(��`�YB�/f�ͺ ��=]4D���\��Lic�[�y'N�/��:þn��	�٥�X����5>Dd�L� ޭ�a޿{r���b�]�g=K�ͪq�.K��TU-��rd��<�]Ց��'��"�(�J�əv)N�`svV�q����Wԑ�[�����_������KJX�+"o �Q�(9ݸY!ǩ�)Ѽ��w�-�9�;���e^��k�.�h5�*��8k4*DL?��R�J����=��A�l������~_��:&�q���y�Z��2�VZ�2��1Y�/	��A�)�\���ٝf��9�=�lg֜di�^�v��*c\��kg�Y8�jlVhDՋm�ń��#l��H	(�����2�{��(����?G�}_W�^Xs������_�
JI̒�wWts�)Ѽ����\���`:�`ڳquj�ք	,��Ut&����, �e+���|�̺n�7v�.&��"ϢkXL���V��ws ����K�}zXs�^z��U�v�$�R]���ۘ_��s8��M��F�@Q1��3&��ch跛��g��!ݤ� u^PԸ���j9����N|3���yK�қ��ߟ���/$�s�oU��=��˗�U�#{浣z�l�g*�7������
<��9�H{�����<��u
&����	�œp�{��ٻ��UW�[}^���f�~V9�^��c�b��(�k�s�Y��)��vрs�p�N�(�p%&8��N�,Ƒ�l���%] /7k.|nU�:���mM�b`����� �[�IP�W�ov��� <�fէ-kȭS�*Q64�p`� jR�*T� �x�=�J������]��iw�wU�W �c����Y�u\<�֓��Ӹy!��j�ѡ��S���[mE��vn�.���ӂ��$�@Ē�@�O������9�4�9�J����j64�������˾�`o;4�3���A���0;�9D�8է!V�F��u�޶�$�䓳��ȶ�Dβ�6�F�\�`�3lƬ�	ie�o�߽��	�O��R�M�����s.��}�0����	�l�Z�3�k�F
g�[�(�N��N�.��R��K��#C��s{��ER]��� �B�P)�(�l:we���"$'t0.�m��l��������ی��OX���M�#�\�}u`g=+փ�ٻ���x��Q�_(W;��t,r��p���d�9�r{u�&5�81D�[G3Ξ������@�����NXx����e�L��Q�dN���l@�5�0nؔ��igL��X3hb�=�Ө�x��^{<J��ث��5�|�$������������(�<W�������{m��F8���co]�5����9�BjGM|}]�}��j���m�9K�ͪq�.)e�Μ� �b����12��:�n�n0��l/y�e`�z��x�[N�cS2��Ue�8���F��gVPou���}Z�۔㸛n�W���V����<|�S�xT�5@苒�U�%���W$���l����l���P�*Sr�ur����w�<���x�	b� �t�&5�5�,��t�Ѕ������K~wҶ�us�v��V�II9���]���>rN����4�#����s�2)��c6��{ol��;6ݢ�c�a[�m�@�[�ӌ[F^9MS��v�\tŋ2]v0k��;,f�L`ď9��$v��а!n�;����R7�Mil;><�n���ۅ�{m�;2Z��m�
:�l�{��w[� �����+T?TU�W��F7%�p�O�C�Տ�
tO(�Ȱ�D����U��-5p�9���Î��C�Z� e,�T4諺���egV]��`s�۫�*�$Q���T*$�g�s�uIu$q]9^���O�a�%l���m�2�
���ۮ����gǝ��g��cYv&�nTI��� �zT���X��������G>��B�P��;�w1��5tݽ�~��>�舉��J��[y��y֫ݔ�%7�r�WqJ�-n�s ��'�-+� n���(�_�]�.�˸���s<�e��PuV���K(vn�+�Ey�ͫWr�Q*TaVy������m�����3Z��J*ddQ���`���M��n��?h���W �c��<���#r�G�k�����q�-�=��g@ն�(;,o(;��p�RUJ�*�a.6��������mՁ�u�l9��֎�իTm	ɎKn�,�;��o+�|��.����1�d���"��c�����lH�Ss�S% '%4P'�I��d�u$�Bd	�C��儺��
T%&� ����F�qX����q�)A�"�Z2'b#0b�&�!�(I�� ��"RP���C"�`$$��"�$0B�#��3D�2����:8�j"V��L
��	��Q���KPBY,�I��b %Q0B1#�'P�hI@��3�)��(J
Gd� da�A�QK��у�N�d��"CBP��4�E!J�A#�%��r�N�9"����}>`]��:ִ�#:ֵ�m��m�ڦ�竳��z觴:��uA���Ѣ#���ɺ���yz�q�qnu��Zz��ٸLc�Ɍ 1�ck��ZְZgZְZֶ�����SŸ� Ǝ&0��1�9A1�c:8a�2��&:�����z�04�൶�m���k�����V7-j���k.��<@r6���朻��"��UƵ�iWbi�wh���6���\V'`yD$��n��ʀ��a]�m[Nr�]%�]�.�����.�{n�]Za8z�j�M1/-cpV��n�N��3��zހ1��Wm.�n4���6TR�Χc��g9����ַ	�v�!I�Pe[��4�8�N��3���!�q4���H�6�!G6��a�i�`��k���- �&C\��\�Ýawi��M�h��g5Z ;Erd�Fـ ˶�\�"c�
^k�f�k�jmk&�
gm�W'f11g���n[Z��a�.�j('j�5U�8�<�a����6��F�nDa�Ė\�lY�m��W�K�I���G6�FY�;{b�]l��w�6�Ჽ��Ŷ$T��y�/j<������'��UvmY�y�A�H�u�����r�"i�*	��\[����q��R�2�{p�����u��v��v�6����'#��I������� 2��E�@!U����f*�UP7����p�_w����_{��JR�8[P*�Tl����y��f�0�4��hmz���Ʋ������]N�m��m���tی� .i���&�xL�9�-\�I��I� �m�%*&�&�t\]:�:c��5t��bq42Xqj��`]7m�9�^�E\�����粛�Fco�,��`sޚ^�.?j�9�^����׹�W<����qXܲ9�V��K=�^����Ŧ�8�^���M�ɔ[�V}��vX秷sޚX/���3V�R6���=4�h��472R]<��@Xhf�.�Pf�P�i:�%��5nzm�y�uc�κ�[g�Ⱥ��"4�{d�&�zs�ڪ.Wt��n$�ku���3n��-�^��s\ ۮ���˫�jj�ݭnc7+5�9$��s��W�U__�b��R��j�iK�b����w׸���y@��/�$%)�HT�&8X]5�n73���uQ�~�������F��Y�z�r�n���W�����K/��Z[�]]Ɩ������6|{�Aޫ���*z�{��~����&Ԕ�n&����=�`oj5ez��P%I�z#�~��QWE�)Ǌ�������Ł�wۘ��Ü�Z+��&�R���ݸ:�����(5+fͦ� �j�:���wI9��o)e���~�`\���S~��RH��p�;�wG(��SE]\U���8�Z0��8��e������I9$���xN��c
֘�s��6�h�K�¶�C4Zm)�&�6���ѭMI�l�&���K�	Z��4n�d ���D��n"tܬ�����R0�(���uS�ր��,���ݕ�	m����X{���p���i��N�x��V)�����@�!�z�07CeM��ME$�7���Ëw]��ez�yw�֎z���#��e��t�$���� �j5e����V�(%PEE8	.6
+a�ݺ��O*"�E홱�$v�ʺ磭�n��E���SL`7��(;-������\]��6|��Y�ߒ�q���4�t3("ꋩ�*���;)K�i�p������A����\ݧ�S7*�e�u(���7����t�pu�����;7����V{�ŉs��1���;�c���s��m�ޫ��s*wed���M�2�&�2
����0�By@�I+9���]=����*�
VZ����ym��{��nvniqe��U�w/ٱg���n4L�u(��}���u�s�p�E�T�R���³-����R+��۸4J�ڋSs����̙5���s��Oi,���D�'Gx�r���]=�ýݺ�3ޞ,�f�3}��JR��P*��z��W]���e^y��t�e &RH	"&I���Ih���5�9���諿���+����-�'��1�'�%�Zn��}��6tO(�#��>U���Ԥ�Y17�r�C��;��w:��yD��4�'/����뷮��*��ŗs$�{�n�^�� [��D�;����;�,���-�	n8�vi��)`n�n�q׶�qx���w����ymhNF��-[r��v��9虃���y_���7�w�����˒�E����=��{�7}�V=�[h�)u��M\�����:��ʤ<����o�����vbc�7S�j���؇��ͪ�W�`��ۭ��v^� 5x�M��\d�n�Y(VG�@�э�;[0����1ʞ���]y�ggԔ�8t�3u�]T�zXi\���k5 v.Hg~��w�ۚy�m6��B�h�iY�b��&����{�����7J��AԬjf9���f���m#�ܒ�h	�]�@��12VۇqRY�Jبo>~��}��}l;���F�ַ#��[����oG#��� a\1]��y!��VS��o���(~�:���Jc��X�R��e07��_��O߱����A������ ��&�2�2��+07�����$7n��v�Yu)����II9����H�`~�����^{�� �C�P.�ͯ.{ݡl���de�V� ��3�۫3E��B):K��R��R�omt/L�1eTLO�s��递x� �<���Ej�x���&��^������m-t�oS�-\m�,q�+�V�fb���qW��������u����/�.]���MM�ϛ�E����Y�X�����ӓ�˞��f֔-��鋝-q���-�����h3�������A�׶��W�A*�8X���+A���`�o(9ݶ`���θ��UՑ3Q�o��$Y������#9����d�p���=����tSДIq�D�t��ꪨ�"|���j�y�&�[� !9O(��u�jncw��������` �t���5��K��]��i�v%D� ��G����w�u`g=4�П[��Mi�o{іBu��\�g�E:���
�El3���aŻ��޺���ezќ��s%ݧN�����ݾ��}�_UUUÝ�e����;͞�gO-��ڴ��C�T��u[0&Uwed�g��(�����O�)Yk)Gx�q���W�}UK���������0��m�9٥��ѡ��$�N��mD���l���Y��В�:rJT{pC�N7.���6x������zA�[0�쬓�	�nj&���~�w�z���-�Y���\IUs���� ݨo(���z�8���*5��֬����;4�8�j��O��p�G
%ē\��O+�T��p$� �V�+�F�D}�U�_}��[�k���\������J�nP��;������H�}*�z���y��%��lĳG��i�K[�;P�6��7#�K�c�r�ƃkB�/�>O}�������B���M�UeVNQͭF'���Cn`Lǽ
u��2d]ۅ�	���������J�#��Z�JeY�8�{m�����7����8�v��R��j���%�nRpó3���e���N�ݸY&�Hդ���K��mUŘ{�o�z�u�^{�[ �>��J�4F@p4�7�Pl�4�� %���C���X����L,lsN�L��;@�"0�� �3E�]d[�f������f�46�&kz���9yx�$�ϓ�ӵ�[M\M��!l��,�86�J�ܕ�4j^��^�7<P�5��cIIe;���Z�����;6�\�7Mf��	(�ѳA
�DƎ��!�LD���V^8�p`�Wo
8g�W`ϴ����R��[��V����mkq���ݧn�	%��:ݶW>��5%$��ٚ68:sE�l'Ջ�&*��i���7��'�&�Njb]4�x�vR�+|����ҥn`(�b�����@�\<�KV>H��s���]�^�Q�;!V�FYh]i���"&F�ǲC�Q�eޥx�������~@�D��arI�Zo�a��� ���
�z��&��:"K�'+*��r̰�u�`�j�֟8����m�,?{~t�V+ʶ�5�ݹ�~�����s��rs��tHX����PE"xF�H%��߿�����o�}�z�s��y���̋F���P�?����d�O�"����UQW���������_���(&'���Ą�P�$!UA�` �Tz�EDN�t"*� 0 �� �� �)�vb��J Ei@�/\�)J4�JEA�A]� WP*�r@�E^ �  �X���) P �ښР�!U$AG��޻��	�Gz�����EDh�D���\�������������������}?����������s���'��~�/��ޏ���C��U_��7��_���x�DUz?ȔX�����;�BG�*���(�����C�����U_����k������n��?���}t���P/��B��_����F�TA�rAJPUZ�)Hd$)��$"B%��	BX !e	B���$Y	 d(DYFBA��	@IdE!%T� @��YBPd!F�XA%!!%(EJR@XE	Q�$�%U!(HEd A$	IERBd!U��!$T$"QY
B`!B$$�B@ !�Q$	@��HE T%	Ta	`H@IEB��YBQTHJDa	B�D� �� �$�!BD�!HBIB�$HB��%Q$H (HBU�E�$T�� $	 $�! �%@�%
BP%	 �$	F��$�JE)@�@�
�!@�F�e	 c
*A �H �0��(�B3 ̣B1�#2�J2#+ʲ@�
H2����0�K��#+J2H0��@�� �����������������0@
�/�O�?ܟ���?���4��Ht?�P?�����8x~7���*�?���M���G8����?�v�������*���2�C�!�_�_����*����W����vhP?��R"�����v⠊�������?�;��M�"���7������=(��������������TU_������qǯ���q����7���"����?��c��*����O��x�h<��p��?���������9����/�/��@EU�;	<;?�1���Ϳ��
;���������_��ʀ����?�눀��Q@�����7���������]������_��PVI��hq���5W��Y������������A)( Q3�        :  �������Z�J���|Kp� )�
 �0�ۏ ( {�@-�  S��a�+����=�:(�;s�� ��s�pС�: �݃@9p�=�( H(�P�gq[p�C�t:��hӜ=}���k@wg[e������C�:և��/���נ}u�n��׎��   S�`U*j� 4      0�Ԕ�4�4 �   �Ob���M�db4@hF� � �S�j�	D       � 0�=�O�?J4��=Sd�<(!H@��� �� @  ��8q�������P����A���ȁ�� �#
�� ������M�P,d�&;�<�_�����P��M�w��~|�e��^��d	2�~�V�[�G�7D�� �
�8��?hoR��-�k�D)�J�8�4��T��l)κFeD�$�m��XV�ԄPTEH���m�|���S�<����q���]�>�qE!DHb-a>��T�B�g5�P�e�����s(�����H)$��XY��%�"oZ;ʗj�73��b05J8���
��J��ZA`	�Pڠ�(=l�����]�2�N-�	�9�`���P`L�۠cZܛ3��	�ë.1ը�!El7"CA�b��(�1# �U7@8Cx&;7EPc��;j�M9w����c���E�\�<#Q �4O
p-ӕ*a0N��
Ŵ18���y<.�=��qРH6�XNm�Q��,'���͘�Q�r��^n^l�
r�
����42���bk���4���Z#zxt��ۦÌ�p�����F��,-9�4��de�83�P�*@�)$�h�#ѭ�fg�����w
��f�%��B�M��"�� ���Շ�f<�#("�@P@5h""#� �7���;��w�3=��*�H@��uLXTPYKV��~�Bq����(MZAD�nD��4FVk"u�����(�f�!���j��H]�!W�n����#E��� ����o����5�Ak���f$���5@`R$�!T ���:6N>l�f�f�dg�(4�拪c4!
��T:�qӮ�,7�q�~�o�{�o]�<��ڲ�س-5E54@�`�PF���L#�ED
a �	���N&�ۧE�K�,Av��;4�c��H�m<4�$�kLl�q"$�N�\ �H�a��Z��cӷI��a(�(j��4�B� ��e �]xs�;��,z���g��:t(ХF���F�j��kE掳�O  �X�!���b��b�0��%�:3gQ�x�HqM,�(b�&DP�0���
�B�z�z�\/5�c	'��B� ����n/ǂT���x8����!A��B����4:�A�/��7�U���r0! ��1h#:�C�%����$9�X�~3@���A�}�Do�tl�c�x�ծ� 媔�Y+Ⱦ���|��߉���lC���t:�C���t:�C����$��I ��:�C���t:�C���t:�C���t:�C���t:�C���vKh�;%�H�C���t:�C���t:�C������l�C���t\�)�]��d����S!�A.��i�����$�d��1�+�}u����tY���|��"PԒC���`� �sq���r�@���e�a$��t>�� P�t:�D�I����w��7ʒH�Hd0H�C���t:�G�����O���C���t:�C���t:�d��$�����t:�C���t:�C���t:�C���t:�C���t:�C���� vKh�:�C���t:�C��yZ�t:�C����=�=����U?������� ݑZ���ؗ�+wU%hln>�8{�D��S��N���{��l<^�s�9���[�S���F��C���j�"J'X]����g��ӹC
C�[d���C���I5�TxR����4�6D������Jұk$�U.[z�ICJ�R�P$��H��@{�̮;�WT\{��{���.�nIg8c:��Ű�ay�H�=���9`M��jj����x^ٻr�=�p�W���I<��jtI�*%�t�nak{�SD����9����7~��$��,�oZ��+�7wJ4Vv(V��Q[�����d�A�Hq#����Uyzl~������wf���|�ӆ��=J����Ude��|]���1x%锒��lI���n[D���	+�*�
4�S��z�����;�bއO,�{���}[a�0�f��0�6��$>|Gq�*C%���Ż��/ ��+W�Th��oW)vL� Pt��Մ�(�&O(b'��n�z���z�Y���'Q!;/
v��A����\�O��hDR�f֯D����	���}8�=�h�a�J�$�a`��/��[T�r�ۋ I�$�<��=�p��[��s�0х�h�z���Z�Hwwf  p:����pZh��`�H.�ΧC���/-T$trN�:�AP�t:�edd�3�F]��:����(�>S�
�!xV���t:��.�a$����צ�o�
���I���t:�C��2$2�E$��t;%�I%�H�C���t:�C�f���6�`BE�6���࣢�!��Ҩ��| �H����@�ImImH	.��ٰ� t:�pw�
����J*g��_$|eQC����Pl̔H W�$C���t:!�@�t:�C�[D��-�@��f ���� ��t��B�7z9�A(t:�C��儒�Iv*-�C�1_rl �t:�:�͆J�w[m���
�K�z����"�.�v��wӛ��E�d3j
�{�k��t,9K� ���q=y���:�	$��u�M�o���R��`�d������H��k��DT�=��~3#��4:�^���z��;9-ܥN�	��@�qx�_�7ǣ��!��s���c缵aW��zwB�޺\PP�2�"-J6X;ڷR�D�Ԑ3\��KA;��M���OI�-�3a�лm��:qu�s$�	���t:��P��Y(���C��-�@�n�C����TZ�L�	�[m�O+�1s�\��&�-��Nt* u�$�z��k���ݸua�[���D��fp�`�8 |�!"P��Hw�o�3 �ܫ0��+���D��pϞ#��ī�z3�=���s!�8�ݡ\���U�4�N�"=I�[���ͷ��d�V��)�9P��Z�=��{�ڪ�g��K�-Nl���]�C��!��:Ȳ&��,�y���W751��zi0|Q1�q��[+�� ;���)�3�A��1�:M?��u�� ��W�C��o�����w)�<��ȍB���P��XA�(v�T�/B.�DDA�L��"�S�}G�����b����6+�/H�JpYG�T4�"\�c$ �.h� ��D$;!�@��(&�;@�4*m=$�&�`�_AO:�v' E�
j�������m:E�Trsj�$ <W��*�HT�����5������NNNrvٜ�'t5�늪�EW]`�v�ea�U�UV�^kf��.�xg�b���^gb�]���1۞�s�,e/ٮ(��-��٭	�Wf�����]ƺy����$�s/f^B5l�ǝ�����K�F�d40 PF]o���<#�Te���\��a��� N�H!����������;���sw�ٲ��k<�0vb7C�\y����H��ٶؒR��y�m�}Ч���Uz��>�x7�k���m�۾���wR�\�(F�+�tY�	E2�)l�hK�0��n�e�sM����%���o�{���6߁_5��ܢL�}���H�Ԑqm���vba零m��6���9��bo��).����\EY�	��S�����M)̦s�`R�1^#V���e���aٿ{��4�"3�gh�廜 ��3:�����nn��D��S�y�}��$�tךI�ґ=����0�����1vuQ����Еm8�)GTFP`���w�l�����{����0y�`��~h`��m��r<��"��B\��ś��&˄%���}�SǨP�� *��@��&L�P��2v�4�eo1�c�∭[�M�a���;y��#w�7�v��7/���aO7�ys�!I�}k;wo�dZ:^����ZH�U�Y߹�f��iiKe�u��X@���"An�M�������=\�����
��SmF�٧` ;����H8w�>&TM�Ŀ����nl�!0�-��!���k����a�5d]����CMa@��b=���P��#|��ﾌG��֮���ݤR"7�Cq�փi-q�Ð�L��Zr��tk��"�:I�j@��<��i�5�����!E�3P�/��;���jȶ����C�ܭT�H�|B#�nka^��\J;i��[hza�"U���,�jE�\�����4֚W��[��j�B�ˮ44�|7�1I��!5U��C$���5n�d_���.�҈i�?�
=��8������ߞ/��zqc4���\,�1�8�XYh�tlH�$hN0�٢bѽk��>��hB�
�w���v+����@Kw�Mۍ�0�'^>�w�}�|�[ DE�h�s�b�v�&�@\�""" ����"":8۬�9�f��b���y=2��H�,��f�Fɞ�,��4�<NW�I'&�r��^;s�A;��:;h�N�Z����Iۮ�v$��P��V�����맧X�����u%(��Æ`�5�
�mFȫs�4e��͈r���v�J��Ӵ�Ԑ��
��`�����:��o�[�4��5�^��̉��H�}��N*� �������һv�m$�֚����
�����!��"�+�Y�뱦�֚�C����4�f�eU g��7�htZ�$܍U:��jC�8x;@���v"�#e�۲(㙎��8��!��j
.#�׈Ư
 �B	,n���Ց/݉]ڭ#��/��I:�6wP�>{���{+�F��a���u���T=ĥ���$ [�m"�^5��������Kt뮺v����X.�D̟�
�L$��o��Vk�Yhe�$�i@�B�w݊]�4�hi�"��(۬�XF�������5�t16>-1*&� ���l���]F�R9x��*�s�����x׏�{��!�{�C^5d!w��q��0� KU�PB4��c�dJ`�D�<F�b�R5m��4�V��{�������� ٯ4��\���4��Pcƽ�7������!�܆�����@��!�eҡYGǛ�<��	1r�f7ʙ#ƕ�,��cMa�5��!+�4�f��/u����4����~�6~O53�bܶ��-�[g���=d��@Z�eNn4��>��z-o=z������^4n���iy���-[i�ÃMa@���]����F�P�gE8�q@�XB=��kH�>!��l?8<@�y/�DA���`B=��o�'e&�ej1Q�4i@�L����Q�ٓ2��I*�!<����K�Zi�4Ցm{�J1���,��7�c��f����K<�!�o�*'�4P���q�� ֒� �� f!��ҿtf�U����5ƴ�7~_�5ZF�	k�}��HkƬ׼�}l���׉K�JCJC�+�7��<hIa~i�U�B�w�*���d���<��i�����̈�P��0�P[�0���;F�k15d"/�r*�C�
�ܗՈ�iDs�"<i^��-��[�4��SP�+�W� !�+���[@V���-���v����{�; 	YT"��yO[]\W916�5�2�siA�
�Dt3��۴ln%H�:8�w�]ڮ ��^e�%l�@�Cu-��0L#�F�P�gE8�qV�d l�s55���|�ĺ5d#1|Gn}�x��*����x��bR}�cC�l�8���H~~��=6i�N<&Y����tY��f�d�`��D�K2��6tٮa�����7���،:vAF�7��;IzΎo@�D8�*)X�w���$�#��R�kM����
�rqh>��/�F1����Z�C�jnfh�A�]�;nl�sj(N��&v�͕�]�Uݍ��9�	#rNL�������Z�Z5k�Ԏb9���aWP`�E��䞽Og��:v��Wd��~t)���,�J?��d[�p���d_��%����#�a���~��dij0���p!��!�.u�>W<�1JB�2��2��޳z���bj��`�%'�d%:��6�5���a���(JN���%	��(JO$�JB:�2G���Pn���<��)�A�D����M�R{HP�̡)
N��ԥ]��\˘�JPy&BP�X�P�����
��)z��7&k���u	BE�BRn�BP�f	BRu&BS��.��:�6�@�|@f�+��_blF(J���JR��2���B��]���y���l�z��=HP�f)HP�JRy?�:����MBS�ߞs87oHP��Ò%��);�P�'Y�P�����RjL��<��):��P���P��)HP���Y�ߜ^o�����MBP�����L�����C]u��-��6�)y}��f�V�Y�7�>�ԅ	��)
Oo ԥf/xh��5��{�����L��7��	I�䚐�.�L�^��ry[קּ!(O3�)7�MBP�f	BRwBS�������d%'~bj��0JJ@d�������Pw��y�:���u!^�^�d�'�d�!�`�r{u3��eZ�ⱺ�!,Xnqg���q�^ݕj�&R���lF0U�;�Ek5��Zސ�)<�$)|�����f�-��k\{��)
N���%	�`� ~�AdRwl��c蟞�P$P<PJ���j��d2��2R��u_{�7)A瘚��;�B�����<̥)uϴnM[�_fÒ����R�I��%y��	I˹5!M�}}���iMH�I��%ՂP��y��J��(���z�ԝI��'���	G��ya�>���Y�;��JC��UP&����G�]S&D)+q�˖R�]��P$z�}���!BRw�&�(J�C!)<���.�$({����.s�R'��!I�2R������MBS�;��_s�С(|�$(H���P�$��JR�@wϺ��9s�]l9	H^�%	I�x���<����2�u���\�a�R��A�J_5�>־ݣv���ǻ�
�P�	��.�wy���r�j��	�9)H^`�)Aܙ	B^f@	I�X:�������4�HRy&F(!�̤(JN� �%	�`��H�@w�ލÚ��P�$^�d%&����B�	{�d�rd%?~��.��hP�����
��R�I�� w�	@u����A��u��%	�%�뛳Y�{�ٜE�N�(H�)���A�J<����\����Z���)<�!(Kv	BRy� ���0J}^���é5&BP�a���H�JPwy�(Ol��);�$)�w����s���);��p��Y�S�$��{HP��R�]���I�g3�A�K�L_�}����L��>���)<��Rߖ/y��w�9!C�)C��翭l͆�j�늟��^Hd�ڠȠH��B� �bn�:oPV(s{�èJ��(JNoG��1�ߢL��]B�x�:P�~��]�5��j����l�����;�W� �@�����][1�WV��%��r�/8�N;[s�jڙH\+,�n�NI9;� ����(��8�#��(�i��=��2���j�ʺ�6y�=Ǟ ��4��0xՐ4��� #����x�5�Uf��bwd}B��	�x���wȨ��C�g�v�JB[f3|E��/q���
H  �*��9����'9Ǣu�m���B*��@�K����e74�ORst��yƙ MC鄳�i�����^�T�}�O����<kW�)}@�B���2� ��7�/֚@���-��\��f����$�(6��\5�!|�#��V}�8�pM� 2,��D̜�`
k��c� _M����ˀ�����ַ����@�i����.�U��G
�=�g߶(�C�|?ys���X��P��OP�ߣ�f�۸!v4��}B���������f�k]�ZD$�;���HP4��d
,4�!��P�]�t
t�A"��sJ��!
!��I �J ���b���"""6���r.��;v{nj�*�DDm�DE۱�,z�{�GOl1�����.0�z��͞gnְ��=^��<6�e��e�ɘ�B�b�d���ݬ��a�"�Z�C*y۝��	V�Z,��(lGj�H5���d�+v��^�	Z���\�BU��y��wZi�ҥJR�����XA���"���~}~������^���~�B�����l�^ ~>d~	�A��G�ݏZQ��l~�J�!�����9��x����ZjZ� ���i6<C o����q��TG����|䕞]�jWA��6Ǌ3(�ݷU������g�q�[���`�D�A�P�d�Bo{�y����,|(��#�J���j��
�6<j�"�Wgؠ�i�@�5�U��wdi��T|kƻ�
�{�a�#�3�~	��x���o�Ia���@�C&�
m��)�m�DDXl  �ɸ���c���@�=�4�\��r��(Q��F��_� � ����r�,�b�i���)*�|�g���럛5�Y�~L�,@[5_P+�*�}�7�q�qtYA+�XE�}@ *��?~^)c�o��\h B#H�Ps������~�'��:����h��??L�@,�|��~?���4��K����1c	~�������|B#}�/�$�����!�p��
u�O��(���ib��"�*��-�f���ߞ����Whx���(�5�/�`�R@���W�P��{��r�,A��8�� ��������2j| /��!���z���f�R��;�"����j�)Rf��vx�N�����G;h����]-.0�/ƕ�N�4���J�ʀ����:f��Y��a�b$i�k7��9>��#�i�f�����P�����"��<�UP>"���>�֑������F�«�@o�Yh{����rr/]OY�ڢf��Ps��u�4a+r���>"w��6�:��@~SGs�����=�S����FP͝��~sZ���}�s����W��jD`��e��r���z�i��P��kG�"��Th���E	C���'�<��c����O}���PR%#Gs�ߚ��[�lB��Os�����[٭i�r?H'��@�(��c��~��v���x���UGdg��f�Ai��!��h�l9�X@ү2(Ɣ�C��Z�|�ǐo�z��}���R7=��q���:�5��9���d	+��@4@���E,xP�G��:�����Ci�"_}�]�k{�0�TJ"�E� XG���W�����`��d���C�~�G��j44� d��ߚc�U�x�4��?��?�T�T9֚�"�~��9$.U�j�i��Ų�4�frFE�=�J2��v���^��Uw��5�uU�~���!�D���g��G>�N��VB�ƐCMY���X��(�4�|�˱�������e���x�@�C�C/�}j�?
l~m�m�q4{��Y��y����1�`	X!"RH�	d)H�#�ve���UU�T�rfWU�n���j��j��N^u\�WZ�Gnj;vLq�W6�AJ�q��d=�M��R�F����Tt34U
S�0�IR<���iĻ1�c��-�7��o7�0;T��z<����N�����]���3��X�&l(SeB����E��c�}��i��_Zhx�4�k�����f��5�Bȷ�ȟ�>@^��^#�U�3P���\����ZF޽yhIi/�����VG�h_���2���I�,����+qT@��jk���6���i��4Ր��8kukMYבG�V�u.��f3���jq-i�(I�Zp@Z���^[���U�Y�֙��0�OE��s$������;�˖�ꪮU��j���ScH�_y$��R ����hiwcBJ^X��i�!G�C��XF���Βƚ�4�-�N�#5*�{����F�R�ۢ�\ܣ�qa&�K����x��ɤ��*��;�Zk��6�((1%'l֑x��04ٍ�B�iM��;��a�hvYg����B�o���6�v�H�Kݰ���(:KtTQ�L�4��[kB�4EU@&���W.�6�3m���!)��h�`U ��
���H�li� {���W߱1�<j�Bȹ�ȟ�ib�@�=�����H�jȿsz2]��w|��cM� ~�����	�H���FjG�W�.�U
`*��4�!���� Y^��>0i�kMe�=�.�4���\LXR	��<C�m���l�v�"jȳ�n�_P D׈�Ͼ®Zk%P�7�9�tZ��-��|� W׿D�<@��Qn$R![�!���I��
i��f���Ր��'��j��L�C�v&!j�U���vkM[gry�f�v5fL�9��9��U�V�[kN�<���u���0�@�i@ar�H��Mf�ˌ@�8���e3Cd�[ ����5�U��<�����B>s-X��P���!���4~�֚@>��X�2�����fkq"�Q��E(��Ae"�,/Ҩ�4c��f&	AJ�+u"O\���"bkH��.�f��i�;��廬"ȧ�N�&�H���.�P�F�1yxq\� U����U�B�p�jڠ@!�h����P�43';� ���C���;�=�������>�֑�6�h*�B�����BO�ʹha�"�Bo'ͶF�4�U� �()Y��i�(L�0`����h�&�yqT
,�*�#@T�qyZ���(��D���Zuђw=�3����"""" ��Ɯq��<�[v����1���5�7aK�/��&y��WV�6�]���v�����ܧ8��m����	T�k�����;�R�Dl!���b�"gW=�Y�7k���=]��-���ɴBW%�me�ܹ7m"��OR��1J�k��E,��B��X�9"����R�r-�\�:�:�J^�Zj�D�}j��FB��ho8IՖغ�,�qW��A�+5">�N슍V��x03P�]��d�v	�vm��LK��������#�mGnSd��t����r$@ 
��]� �^�[lqI�Q5�W�ӍhUa5##H��!��2Պ�5oN�F�F�?Z�M5�S����@4��U
x�x���`*әw$�US�A�����9g�����tIǌ��1���
"����S�i�#�W�ڬ��4'���n��)���%64��C���+}�9Ƃb��=��!���rTl��A�ߨAu�J��t4���X����ei��!��˂�CY{����C�K������m3B�e�q�M��`�����
��B��6�"�P�>��A<��P�+"�}%n�f��3��V%a���T�LD����U/t�T(Kr��H׈�y"O���Ȩ�a���Mf�i�t��a�c�����4ai�1I��غ-��8-ۍ�E������5l�2�f�T �^���|ߛdi�����*
�C�#1%DX�݊Q?� �5�_�k|��
�����x�ݜ�H��P�]ȧAZO�>���ރq� ^�wI�q�!�R��y���؉�d���h^��i�����wXE�O��!)��V�G_X�p� ]��,�G}��
�5�D�Y���B�7�9��Yé�=s���m��(�-C|������4�[	�����BN�*塆���� ��39��Cw��0A��i��I}h(�E�S����{��}��B�a�
%T �@��X����v�ݜ`�i� �v�#RX��]��h؍4-"j��s&�W� l׍]��$�ax�Y�|�5�VjG�$VR��k��A�j1�K\��\�l�e�uj1�Z2�U���<��ZO?��6�V�eo�f�5�66�
DFj֚>����E]�����CH��!uȟ�S�0��Wj�P�2dQ!̬45�k^a�@F,a�`��u�X�X���łR ,R��;w���+tV�j��*�UUmU�=0bv��S���:�A�l� ]-��vƣ�z�8�X���X�]-�Q�m8�D��c�c�7B�ɸcq6�|�Y�f�f��=�� ��D<P7�~_ �-V��Q��dq��1Lp�vL	�DB��,�x���@��"�P�:�W"�"��s!��5����a�$�r2-���Y� �+F�!R4��B��5�3a�3��87J&
s�7;"�u��f��4Г�i\�0�R!4���#H��+0"a$�vڭ7&e�e��a�Tm5d#�G�:�A��E�޼�xq�:�aSAȸ��=���Z( |E{�ap����_i�*&J%{r�E�Y���J�P�ZhE�&H����*j���m���� Q�!d[���.�&���n�0�L��7/E�무5�D�uYz�-ڧx0���c�P�(P$�˸	�f���m�F
JzB4y�q�	mPN5�S�^��Ef��w"�;CaǛ��֑�
O�or���^�̩P/X��7wd2$[e&Q	H�,E&#�P����G������(�ݏ[�4����EH���U@�;���ykƁ�a�A���v���qu�r����2SA�m,9��n���.aX���cO7�[T¨�SUf��(�Վ�VfP�*�W�ZRv�˖}&����s8�����$2ID��~;���l8�q��{f�חf����7��5@�D 
��n�}�Uzf�;>�����H%����kq�]k-�Y�� *�J���f���i�|��͙I��]<}�ɗ\Lͤ��.q�gR�n���K�oV��+)B���X�!\����s�
�嚥�tPMI�ve�[/��nu�|u>L�_a0�mѽ�zݮ4�"�/�gn�P��n0�����a�ͤSyq;�/Dn�i���m��C�/p�;D/6mڂ���3w��N�	2�E��s�=��)��,���v_u�&�CEU
X���2�U{ٯk��~.re�80K �-�sL�+Y	�T����~��y�� *v��O9?AC 
�t��I�4��{�䕣g�B�{�A�je��ъ��}�~f�iDNәf�Vsb2�-�oL�DD�DE��dŴ��ӻQn�N��]��7c��Z%� �q��2�L��u	C���u5�$�6mpp��.����VNLN�̅[����.��< �@M�D@d֩z�{���[r{IZ�u�<㫍1��sD�#:6Pnv���A�QV���7�~G�@��0J� ` @L�DĀ�-[��#Mqj�|�����Qc!�XEq����d� ��þ���M�)��Z��iۿn�E�녃s���C-��BiQ��v�L����&�h2\��w��˓=6�Hm�n�L(�)$ۼ�\{]���{���~|���l���sC)�U+7��=����@b�%�+ՠ��t�Ws��$�.��N��nwuʒuU@�����]�Fo�{g�!{������a�^ʃ�o��o'컷ˉ�HH8���76҉@�K��� (^\χ�/|
���ۙ"���f������uk�ٺG��!��Ű�bN�Iy�o���¨K�oo���6�����+��AC���}ڏ�c��
4�:^z�з�ӤTz���*�W�������/���nl�.��{�~�,|��V�]A6��*�.s��N㞤A�6x�Y���a2F�%��� ��|��ǘ �����q�PM$y�6�v�nc������T���3��ҌO^��p��u��n���c�Μb�� zoW3��wq�nh���'A��u��ؽ���ۏ���m�K��I���$ ,D i"�f���-4����e�4��
4*���}�/&'s�f��/D��q���j"$.�[su���Ju@�L��u�g5^�]�S[��T�����q���ߪ��v!������BR;���m�!�ݙ�l�8���-�����y�>��f�����F�����Fĕ.,�̒�۱<:�hV�,�F,9t��d�&������K��ȓP��/�
�RIșa�j���l�J��013��Ҍl��
�ۿg�;���@��#g5^�O��Ͻ!T�Y�5�9��I�bbG4nu(� E��8bBD�Ih��X�f	!�.s@��E�sH�@��f�k#P��0{�u���o{���USQ�Ί-�2�
��F�6輅wC��x�:�j�6��Vsv<B�^��c���ѣ�;A#�[D)��ۦ��|���~:3煕y�a�im�rg\v�;�8�v'�h����L�Z�l*�h��qm9n%�	��d�(P*ͺN�,��{���K��u{[!�h�4&�@ӗ���Vn�u����6�	A0��֬���HS�\��U@c ��w��w��:�n��_'��G6�H�C�Iܳٺ.�%S��j������sw~�����:�m�Z�k{�~s��wQ����n��2���st��$Yc76b}�=��n��9�3o�qn�[�B�p��)��m)��LS�6�sE����`���4;7�`���檫r͹3|ys��m�+ם���"�R[{7v���S&m�-{�ͼ�P��=��P��e�e/�Z4���[0�!o9�w7N�M���� ![q��q.��\���P ����\ۗ�֜������36�ft��R߽��~���QF��y�0����t�73\܈��~9�T6���[
�� ����?]����ڛ�<�A1ņ�Ef�՛�%(�$���7���V��~�:9���UB��n��9Hwfm�>Έ��*������bH@�>�3XE� ��l��I5�m�E��k{���nL����E�
)!e��B�׍m��UTO�j:$��HZm�$� d�`�yy�ɼx�)���g��f�bL�(¶�ç;k�l���wF7�7m�7f�F�|F��@e8�y?nI�I�|ih+Ngt���"]�Ee% *$��
�-�O\W�Tx�(r�S
�V���ڳ=���Ԕ��b�)���Dj8N��1Û{���a�EUS͖���=����KJn��7ݠ���G�p��5]3��є�e5z�v��vI5L۾s��7w:��ő�(�� ����L���341*�3��6$	,D"R$b�9 �E!f�5$���#(I@�NS�sO>{V��5�k[�DFiw-��/O7���.��$@ Ekv�����90����In8��6�s��gn���mة�kg1�K\΍PX�\s	-��Tv������X��r�C��U��r�<��a�h�k%���+�l�oG@�f�J�9�ڍv���,V��3�PVj��ؠA�-A�1��R���)E4����)uB�2�P�*��'��g{6�/�����x�\�뽽	&AL�$��m���>���gG6Z"��e>����ܭ�f�������i�a�fv�7K&�6m�G��ŁB�:�f���9ƃ�X�ُM��W��ͻ���=�_|�b|��}����pf#u�L����28 ����y帯4��T Zҽ�ٗ3n�̕����.���H6Sm0�^�����fm���_c	lY��	
vk��oܷt�F�`l��^��/5��tPכ�
��;s��� EY�2��Zsv��W�
y��{�Ao7�^o�d�J�;K�n$��"�G�f��9�{f���9�/I"�$�"KI 3H�h]aν�C����P��>R{������`Ev,���ٹ���L�r�3��-)�m���vba�[� ��ّ�bb(�=V�7k=���8�cZ\p�$"�`�f�ٱ�Nx�Į����ԡ,&�){���jF�1���O�z�v�n�n�	��>�P}3���Q擩|2H+��-�nY�� ��BHQF�N0�h4�
8�R#qle�HY-�y�����سqv#��3v�=��Wv{د�7{�'D@TRi��^ަa���*sw-�Zsw��B���g�B�nl��塼�
������=�����@ͨ�[���F�Sm��o73tپ���-	}�=���ُ��I��^_DWf︦y�
QB��μ����H%�ٶ����a�R��<�=�/�2����3�	�Mh�i&%�%�ac6�c��'5������u٪��P��<.�ڏlD��`�و����������y�]LR��ɺ��HiO`��f����P�%�����y_����^w��M��bNoP�]��C2�}��-����� �~�?���3�*�*���X�
��=� ���>�*� U�����ɛ�~��bJ��4���[:�0A�/����Z��oa��4���k#�ZC	��7(��DU��
�B�Z]�g{ِiN�~p��k�Yo/��xS���@�� 3וv��m���6G�Md�� �[j��~U^;������N����,jy���C�K�O����c8�A	�bI-�T��ϔ`��Bf��,n�8ƟH��u���i��0=���zxx������T9���}@�����~hJ�@H�*dn�����y&�'.@zr�BO`�d��B �v~�GG��--�;?�a|��s�������F�9��U�օ��GЄ��0w;�z�{"������#��rjOR���S��o�9)1� L������[P�Z�j�����l��i����y�����pb�lr*bՆ4�����ug�<`oq��:Vh�b7VjU�5�
�B�$��
���*��J!"� ��J�
��B�@�J��H2*�*��
B�@�B���
0�P���!�@
N�E�x���u�:��<�ȭjX�;r�n�<+r��l��A�9H�*L��p%56M��7�i���s��ß�B���U�[G�O��5w�F:w��\Q�����	�X:#��/;XӱݐC��DUDҜ��q���D�mL����v:CTچEg�I��c����#ؗ��ᄋ%||�J�	���SvGg���`t���v�� 7��&'����<�Z���T�ᯪ��o"�`*��BH`e����_Z�l�d�~\9�aٔP�vv�7ȁ � �T	N�T�&��!�˦Kh�wC2E��j� >�ʗFL, �=�Cڛ��p`����!��4$�<�4�o�h�2�*��!{���
��!�K�e9��l����n������ ��������W���Z_�,����FE��%4>!`PT	)Y%�O6��(�����w�r;�}ۻq�O�U����@��uu�>?}�_����?��Կ
�o�m�z��������wt�w�<���l �>j+�D������W��v�+MѨ���q��)�A �E�:��zB�@T
���2^ص~�>S�Ln�l��o�cӘs��g�l�'y�8I��>3DwI��){Q���I�b����h�A����PN[P���.VJi�v7h`
�""�=)�_bI@ ��y��bE︖I���7#!��iR��n��q�g����5C���A+��ϝ9X�*�/������?00�"��z�^�aS�kQ5ܕ�����{؟�ӻ;���q#��r�v��	��+L�7�2���2���r��}	�����`�)�wBm?�]��BCH� 