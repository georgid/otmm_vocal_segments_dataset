BZh91AY&SY=� X߀Py����������`�|��ሺ>z���/v:+e��[�m�c����>�p c���|����V-!J���S	 CB�4FPz��2    OIRz�@  h� 5<ʪLL�       S�$#B��Q�zz��d h  4�$�d�'�Sj{I$�4y&��D���jzj�"i=4O!��56Ҙ!�4P�k9�C��+eD� �P~kAl(�~,$����{�! �� ���p��I~!\�U�Hȇ��$@(��xw|<;��z����A����O��{��܍���wy{���&殶��[�k5�0`�9a�͝�;��n7v��6cY�Q{��&��ܨ������Tf<˫̌���8��n�����hhћW{y�ws1W���̼�����5�#u����f����lR���4h���ܬG2��;��R{5�f�탧wwwv�u�������qwn�Q��ݽ�իwvssp����**�ݍ7;�:��+n*'�=�Uۼ��"������9O-�P���>R���|M�y�ʢ-�������*�aj�TN�	�r*��̮Cq_��0C3�s��t�X"�
a��t	����E։21b��&V�6�T�2�#SU#4YM�P]#w4���:�6Aq2�0��:�VBz�j�θ��U6��l��J�)U`�SW1K"#T�T��,Qm�N�^�r��Y*ԙ��x���X�a�7y�f�a�M6��&�nnh$�lMm\,h���n3lv�6]��5!�fu�r�]�]���+��9f�.��t�ց"ae�\�c� ���s��}�M}��&'^��M�Ig����L<'e�ެ�'�σ}��O';4q�;K��5%���v-L�]JK��M,������!L�	w�X�kYI���	��n�z-ɔ�]k� �tqm���d///Z��HPF�����͓[q��
9Ǜ�S)����\��*�f�1I@�F��U�wUQUUUEUQUDUD�UU^��}���x��|(EiJ�EE��PZ��iZJ)H�J%(TAh*��J#UE�l��^^I��������X5X5X5 �V,H Ab�J�b�bā
��`@���X�X�^+X��V*�UQ�������Ȗ��%�^a��#{5��6p�Gs���FZ2������)ʗQ!��$cRLҶ�Ⱥ�dĉ��#E<��û�2�T^%�RO�W��i��f-e�a{�W� $"I���z>�o��g�����]��xj~���HH��BEz��������Ӧ�3lo=듈�cQ�D�Nġm1�@��߀�(6�D�!�.�G��2���ηN�)0�Ṁ�+�̘fdQ�l�z�B�%`=x����p��$
#���ت��B37:��І�W~ؽw  v��q$�h�˩@
$�'��Ǚ� � ;�۽��E�3�=�.uю�^�䊡ھ���b�d����2�6Pmfާ���g*��ox�[���FYoR��_�s�[�i��͍kcc(�[�����o\���:o}���~�C����k{��r��/�L�χ9�ᎃ_�MY����f]�������ǡiΥ���K�7��a�6oK)�ħj��O����7z�� ���������|��r�ƺy��*gd9�	��N�&bM�e�� �yxb�͍~�$����tf�f���]Q=���;�U7J����Trn6��`v3)�q��p]p	A�l
�φ� ���G;��f�i�j� KmL��q��c-;ebI�i�]���C���6G��j���,2�0A��Cl8/�G{��AL�=��*��ɸ�~p�� DY�$�#��DVBqz��]�N�e��#��3/���q6x�9���k�F�����nw��(�;ލdz�`v܆m�fp���?��*�%��w���P)�x0�Q�A��{���8��׬��Yl�6��b��o��}�j��t8��ۙEp�eA�����片���o��������T�L����"�Kg�{�7S�dv����7:��h��у��t3)Le��+�k��p�b9/zs5�����\��J�nvW��@�.�An�����Đ�!���R�l��Y���ݶ�;*��r�T��T%(�\�����8]|e}��2exK>!��:�������ԯ��kX��{Zme��c6��Wh;�C�z!�Uķ�!ӊ��z��AJ�S��e�iؗw�vص��4�oN�s�G6GZW��u�-7[-�Û�XNF��^���p�f"���|�wh֟�S!3��Jm����c|m���+@���{��v7*��<|vN�J��9��f��A�ݾZ������&��R���ʀ�������e	���:�CPK�9@��Q��!ap4u/wU����U�ɓ����������!*X�!!b����ॾ��$^�!�4�}�E) ������$�	VqD�X��d�eX�X�]��C7Ь��sy��'��h��s�x(|�:E�bY�ř�y A�V���L�
��}��LѪy��,x�r�Lj��sl�����b��T�Xw.��KY�̡ڊ��O�T�})��W9Pjxf�:"��Ȫ��t�c}�v<�����/����Ο�^��Z�B�H]J��U�7�Z�У�-8`���JV{IǱ��\�=��H����I�W���hMCWr�ܗk�u���S����%��I$u�1��&a�5��bK]G+4��C1�]h]��IPo5���A�2�J�?��j=M�=q�Yf�Q�4FV�q�7~던3=�t�t�0؎rE�9Ȗ�3���|-M޸�c�u�\tJ���9df-ow�t��g����.+�������o�i��� tj�6{^ÂG	��؉b�c�/�=u5�Sn�
y�Zoy��л�8�湜�ZZZ��R��VR[��fff9}�1}�^u���f�m��.���b	#
	.K��xպ�dg�yə&h�+W >�d�o�V9�\�=\X9��S�=���W���z��N�F<��=YnS|O���V����*`,ӡ#��x�]j�=��H;a�q_��^jN{��s�!j�ecڴ\��vA���Y�����<�Ĺ�n
^�P{"��QF���,�,�i�O"E0R��D�Z���.t�oVF62��N%�p��
�Ѫ�i2$�hȰ s-֠��t�)��Ƀ!�DWmr�%�X��@>����&��s=�>[�롾�_(��K�y�7�X{��爸yy�Hv��̿J=�4IC�z�xR�bR�ҟ^�at�K�����óZm:6ڦd��\�7c�����k�a���~�'�m��5�w��^��X*jKԕ�h҂\�ԅ����3m�5����%��]���vu�݁ؽPt������(��z>s�n����dQ=�:+R�Z�X��9�n��0�6.TI������+�u ��1a
"��x��.���}D	�AqK/PÖ n���s/����©Z���5{cW�f�zҐ���R��]��ɼgݷC--� r�x��g��,�k"Ϯ1B�� ��}����繜�FH�f�K�Q�kw!-s~z�Z��!�`J�BY�h@Q.�XN�&�
�h��R͢}S�]G���1��g�w]7ى@��^��^u.���t��^]�Y�2�]1s��@[�;7寠ڵ�3�sڂH�������f8A��8-�DV���r-��ʼ�q,�C}P���wȽ��Fy��o�%��n�Q�]_���%���30Ќ�BI$$�B��˩�y-�Z0���_�*݊�l�\�P�,R��c,A����
	Q����"��� ԰��$T"A3�cj��(�.)1Ԃ��"H�QKB�1�B*��L��Z`)l*4�T�?:�� H�)z�X�R���
2+!X�)Z�5��lA���(���P"���#j�V�s�g��o�M��(#"�H��ng��*h�W�%�&K�f�Evt���D;@�Ec����K�C��X��ח/��P�D�C�!�
3�׳۔P/.q"�����<H���=L94l <*������������I$���I$�eE�z�}Σ^ߧ�F�w��E�y!m\�e��1٢(�X61�5���D8`��~~^��g?�toR���%������!�S���t���<�<�Ѐ/8ҲSݰ
�9�3o�A��/�cAy��ď@j�0W�@ w���
�6�%� �"G�x�`�.oh�κ�e數WϷ�@�f��P��P��G+��/�v�nA�ZbC:�_���6z�L���o����ޢ�����2���.�K~�''�:'�Kd��h ��������D���(U-(#H�IJT�DB�@D �j��@U@Z+�IHҴ�"*%
��$� ��
�$�����a���Kп}B^��iCؑ4�n��2���)��@$��RDP	k��j�`e���\C7?l!6&Ff��b%ߦe��c?�ǌ�lwYh�XX�-4��{�P(�f�:����#}՗R��˯�L|�)�ؿ��T:�B��=�=��ptϣ�n�5G5z����y^|���Ù���Mp@$ �D���k3��p��5j4����9Wi@)�:"�-���/�{_p�(���1}�Ɓá;�LJ$@�,����U��
�HB%夔h����� ��;(U������P�j�w��*+��U��� �4�9>�\�Էr��ʥ�Bj+�QJ��1�� -.B6;}~�'f�c$� ��0@���Npw�O�|~�Z�����7�z�:V�����ë�i s;��Ry�S�n���i�x[��ރe�e��Мi�?�Un3�o������s���.�]!����0�Q�XP�jGѼ���*B�%%9C��̻\��zr�?�q)���C�(�^��e�"�P�:�P����k��m%�֘7�(Kn��0���tMy� �Įt*�E�YM�Ɏ�oR�_7r�(a�J���� zU���o����x�H��u�8t�|�k~y�qq�����x��T�����6����)���8X