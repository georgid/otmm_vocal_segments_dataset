BZh91AY&SY ��3 8;߀py���������`#� z� 87`�î� �� ݀  �   v�`  %� h .P�� Q?��ꪨ  � M   O
T���4m��A�L  05?M*�=F� �0@  �db	OH�H���4d   �  �H�LC��!�O��h�#L�1h"H�&���HSM5=� �6MM��i�;�� �h �� ��a_��!g�PIT,(*��3�ŽI%ĸ"h�A}�(�"��)��>�g���q��z'��ϫ�:�un��������ѻ�����wwwwsN�������ݭ�{������3ˡi�hX�J�)t��`��fqC��&����#4�$ ck� ��:e1D-�M�&��(�-�膐�-6�9Y�KD/��, �82�X`7��;R]:�D��i���D�h�^с�i�кh��-�w���c�1ش@�V��]9a0�4��uh�DJ-������k-�Vd�"jZWDF���N����S E!e���2�q�YtZp�ٺ.�c��-+�(]7i no{Qe�a3���i����N��"&E���h�)`�Z��v����R���3~y��ǀ���;��Kr�Fw��n p!�Bz:$Җe�70���9	s*�[d���T� �ny.I�k�n�i��VU�+I�k2Y���aƯE-��ȡf-ɬ���J��18�^$q��]�:�!H-@B@�C8�bU�d*=ж/vKe5t�*�x`��"���j�J�4�]�8�B�]���۝�5U��3XF��\`��en�����q�R����1�B��^�T��I�Jj*\O���̮�,�)x�Y��L�+�}
{,bH6�r��F�@��RS�P�+m��^����ۊL#�ov�x��kZpDe�{5L�k#ec�Lkq���PPԥ:E�f&L����)(���Zl\*��g��Ǘ�=��f�lT�ڔ/�v��su�M!a�qi��\�ɑ[�ml�ܚ�X7Q��Q�&�4�P�ڢ�2q�b�J��rL\�R��.تT�4~l�A>(��R���5Jm���Ѹ!aa� s#�lJ�5��k����]b-�Bfۭ	W��&&���i]��m/�Sbj�v	��q�Q��oO�O��$��W���|���ݒjjQ�FLj�4��{l�;�i;�{!㝰��Wi��o��eb�R�����͚n�,tn��hR�f�&�BR��6ԅ�kʷl:�keZ:�hs&[b�443f"p*��٬Ԍ��̹0ke�A�2�{�vl��؊!���?J���l����������|0h`�����븡k���R�'
c�zpc!x��/�W�������/np:��)� TTL�^��g�2��*��A���5F����A�*f�~}�O R�޳+���t���41JڥFwCt�v�we��Y��&M��L*S�=���5�qD\�lL�"�$��\�����f)`��E���e�ie���l3���D�	��b���)Qm4�M���k1�jLhk�+(�,
02[�d�޼g�mv��v�](�@/�������o�}YT9̴�k�ǧk.*cK�/K��b*a�N<�ެ�Ȑ�T�ěu:[/gC�(�x՝#iC���[XD0��^8Q&vMz��q���UՆ�y��P��B�v+tdP7saL5c!���"�����v��c['T!J6��X��W�EE\����9&\^�H��*+2I�"݌��i�K��e��k"�#d���9�S8rf��4C!�����Ý��VX3�W�"�#:�$A��=�h��P���Ƚ;U��瞇v���0EUUPl�+P��bTo-�79�IS3p�_|m2���P��*�L�i/�g�L\�h9��1������|'���O9ˣ�5��t������T��h}[���Gr��Mܞ
P��D9������Ȭ�n��O�m���������f�O����&П��Hϛ*kdb߲aF��Sl�N-�ъ�u�P2���W7W5��x%�{9���:���������=���	TO=͘�x���nn"#^�lk��������7}��&1P> a�3��>��u�#u����D,����c�Ʋ;fbg��Lhԧ���Ō%�'bC��s��v���^��
�!��^�F.���T��p=�pf���Jѫ�2��ʹs�~a���#��H����<�RMA�_��ᬹ�p5eD]T7��ھ7���d�
�r���2-��b�#�:Tፅ�[���DAQ��<���S.Ы�|
!�QZ=�v�Ѿ�<��r^�
�Z���Z6�4�t��\�ˁ������|�H[1��[�W�xH&ԟb��/Y���T��b�8e������
�9���q�Qj/s:,YkD�1�`+7s��b������똁$�>�E�;�/�Fz��oR�/�WUeh�3��&�Q��y��G�ż�����^�js/^h�,�h�f��쮉�0��vTf�K����SE3WEՋ�8�k lsh-����ou��ŕ��hF��W<  9/�����bn��k�Z*��H�ZsOt뀹ބ�2ݕV�o#\m�ħ�����/�  @�/�����:=���L2�ی�JtM}^F\:���>��C���9��V�(gDLD�D�S�h�z�6���N�<x#p=
	�&&F�+&4��u�f*���.Hv|;%����{������{1e��|�p����n>Α�d��S�W�$}@��g�c�"u�YB��&/�1!�*U�FVӈ�@���dm
W�=.���h{�^�&� 3����"YN�+3v!�a�JЂ,��*]�CR��� �^i]AB�bD�7\2kD����y�2�K��<������/.Tܸ���{�TY���J���q�{���#=�pV�� �~���l�RI����3js#��0�M��i֒������1F���B$��sN��X]������+$#�\�g��!|u�k���8�*��Hϵ�%�I�h���2e��G(��nlR�;���&��Vb&��"5�w'\��u3h�O�����TY܃���!s�����8A�s�a��$�$?xډ混��݌�o��w+�y?�=�5֫��Y�5SĞS���0Ḉ�#i����,��z�fQ23ǩs9�Y9>��Pes�S0f//��燍&�A�6.�o0�e�����ll��y���s�w�F��#��r���m��XWd�ؤ�N�Z�G��F=�׼�/(��_Ev�WC7u'�R�wV/�A���/�a޸���2L(7��V�Rέ�U_�H�~(z�Y�gW�ʢ �ƍ;u���R��/R��1���_25�\�Cؼ�8ƌ�rB�_v�l����*�>�Xl�V]��v��F����#]��/z�S9�B�y#EBۻ�ʭ�ꩫ�,�!N�7�����.���j���3��U���?X��o�h��Y&]^��;o\��2s+#&27���ڜP�M�3��i�b7<�f�ۀ!C�őH�;�uu0;%�À��DtI1�U�OuTp�e�-��� ���C^�?�j��f�ըa_׷U�
@�B�0��L\�E����I��E��N��Eyj��I��C���|Z0�Ѡ��]��ٷ����D4a#$1d�FQUTh��Q�U��8�]���.W�-�FV<ټG*7�]&��:E�h��2�ڋ!H� %��Ļ0��MZ�A�K0�h�X�
����aR��L3����D��G3�9Ɲ�B���vk:�䍡%�ʸ��*A�t̰��4�٨z��_l#�r�{q5	!�Y>r�ہr9�\�D�����{�6'.h��DN�M���u~ ����Ή	0�,(���4`�C�9pzk$U����T�3z�m#l��7�uDU�/;1�ɵy�/�l�xa��	$�Q��PPPEDJZ�^h1뢹}�Z�e�K�2����Ր���֍}q"s�����y
&�(�#&�2����<.�z���1�r-*����>�Z��[�}�}�HS��j�4-=k�N�k��r�^s� ����B'C��h�"^���3�5��܄�;�<Ù����<T,5�j�d��Ě¶�n��#(���m������4�`�+�C�h�^��o_� }�BI�>���x�'�Q�5^��:�g��Ю�޴�s��M6��U�9�[1�.��w��	�]��(nج�TtL��a����2E��MI�{3zl����9�A�����n*'�BV�[<��|
-r�^ˠi[���jkA��s���q�v�9�J#h�U;�z�N�a<�����؎ɣ1�a{$��W���8��U���A���!�Ug"�w�o�u��t��K��8��F��A�3�k��v&�׎�e�|j���&U���P/A�a
�'�9BΜ8�N��ׄn�c�]Zx���D~,~"����b�ٛ^�nT��8���'�U#z�8MtY�;b��j���D���ˎ3��ɒ�X��͇�W����*� z�\�$\��^z��TI�����%����XԮo02 �vl0Gtйe4	�'��4�ӡ$�	 ��e#� 0�,����{T�]���RЧf�P���h�#:wD�����W>O#z�,u�л*{�b1f=#���T�ɾt6H/c=��R�+���k��Æ��V��n*��n:��hy���p����L����	�!�{8���]�۔:2��o�#��b"�Ψ\�s�Ԋb���J�"����Y~1*�Ô�Z6�b�}�5�(/�:���֪���6��ΚY�op�ygj ��N2vRhŠY�4��i�gL�#$'��W=� �okbX\#'fhZbи�Qͼu�;IҺ��k����~�q��tB��o`![!���
8�-=��  ��g�ʃ��&��i�ΖEY���0s8�\UiY��o�����n������K(��r0���Y���	Zۈ���hV�9[]�f��$�(�
Kѭ��;n1Ț��}y�? <8
����vu���>Д](���g>�H�'���mT�n��|~�$�ƳL}*�}~��xdM�_}��u���Z�^�<��7�|9�4=��KH�K�TUUX*�G� C�����x�6x� ����lK���a��J�.��\ɴ�U@h�XU ��jxk�l� �D)RD!�(H�3T���B��%0�D �E�"�P�_B�X�b@$P!��H�+�VF�A�(��B!"���.@!�� �ALA%��������Z��G(�T�P
BE	dI	T�YP(����H9�~q�p;��i,PP��?|<��$�D�M�Z7Z쯷L{���x5bv��&{)竷��G�X��;��i���ǚg]��n�0�j���o����ԧ�<��5���=V2q��5�)�Ja��� �� !|x)!bC`�as�+�[�Z3c���{��"�d [��[���PU� =|��<�?Wϸ��k�^���W�
g�>���p�!B���Ff���H���������2�c� v�WWl��|�\-��������8OTo�B�D@��-(R"��� �B @��BQ���E� �͡@HQ�Y3%g/z/��x}f�Ř�|�����D6TP$T
�TE@�P$T	T	o��᧓����v���#��m�dye�H%�1D����z��S-���Y9I%��L#����2fo̖���A@t��2f���|�*q;�9ɜ#N��SMr�|����Nb����� D�C]�u��[�x�hi�����1g��;�^��֌�3��7A�D� qD
�䚘b������0�HC�,rېG�wtUh�P�==���20�i ST� ?��{M�h7s�6F��769-����U�2�W�v| ��1�PU��)W�;�V!(Ǜ_��uX��>�)!5X3W��R��+�cP��')#)A���p�i`�)�a�4r�`� !Iш?f<��w���6�����p��Xy^�X�SEZ��S+hq;��0;z�{��[�߳ 6oy9}�6���ۻ��PU�t���K�T��x �@�-�Pu8����� <�FW����jO;�����7($�0��>���!�Ez@;f͵�^ܡ1� PsH{n��Bw�GCM��g2-{���n����ܑN$#qL�