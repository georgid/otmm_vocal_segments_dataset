BZh91AY&SYa<�� q_�py���������`_}�xP|�>� *�    � �>;���Av݃pĂ2&S�	��ɒzi��3P#����i)I�2��@� 4S�OPh�4 ���  �H�@jm �  ���E<���zS�zdOSC� 4ڞ���m@E���M���<S���h�� ��Z�T�I����UD� �q
��F%�$��D	D*���T?l���ZO�B�	�$�F
$�bŁ��.[�}� =�j3�U��9�}�%a��,�(�B(��I-�]�q{�q��$���.��~��ǈ�!�!I��~<G��L�t��!�"�)%)$����Ǐ<G���ř��T[��ZņW($%Ev�F
�&��>�5�e�̛��7�z��06�r��=�l�'fE����p�8[5	�=:xq�H	ѹ���T�GUR��	�DSc$�Va1���"gh�E�6n-J�xz��[�G4����;STצ��\<�f6	��]A�R�(AM�m8�R&���[(
r	SIB�a�ꁄH�A
}�H��"���&�\�E"A��x���.er՘���ܐEY��hV�b'[�����ۧn�&�Ț1�j�i�:3N\����ki��w��}S���\ ��7��P0'"MizhO.h�y�}?k�">ʈ�����ws31���30�I$�I-E���I$����I$�`�p*�"�^�*ֈ�������S�y��U�d\ͨ��&��emRr�����a�UHX#rgX��tOT�7Ri���n��m,�x`Tճ}}x����A�ԇ!M�7��2�չ��<ﳓ$�{#�=ks�r"�~!=	2mÜ��߬Qk�ɇgz������a���TQ9!���C����J�ƒ�	�s�t��_VV�ڈ�6�Z����:*d�mC}|��V��K�`�W����} ��v i-�X-vE�p�N�0>��8�,�4Q�yr�as�P�jh۹#�#���� �[�K5�ݽQ�1�Q \84rFH�r�(�bg�ž<q�1>���a�_#�ѩS��C��+zv�/=2�.tZ���7;�F��<�8fϙ���B�xg��3��)���e����zZfkM�11"^+��l�ڇ����a�R\ �-�	��x� �p\��GC��훪 G8�E�lG\�e�����{<A�ͷ��.%�_!��I���h��Y.�Äe�!��
w�`���1��	�����#E���ľK���gn����
��O��峺���(`ڠ��L�;���;>N�SA�r7�0����_A��82c�PZ��D�RU��|��v
��s���x I�PC���+���"�S�>y��+�z�<��u�_6���[�W=���,@ @,X����y��5v��r+&�,ν�5��h3��;�Pb��-yڭ������f.���q�	�1в^�^���}T*�?�]�;#*U���˦����;��ٚ�������Oj2�z�B˧���r9	���p^�QB;�m���쎆�񫴆H6N�X�|_)��BK�O�*�{�k<�h�>����*��-^�
��`p�v���f�R��9Ψ>1e��O0�T�Pyj�F�@��4�����FH�J�k���ŕ^���E���F�$[0���J����<��;��=�p���:�Ղ�K��{�+ͯ<P��O�0���{���/�4E	7��M�EHY��b8�Q�I���`�u�];��!����̈�ȰE����7�ݜ"ܧ�6�<��x@����|�߆�A�"K���S�"��7�w��z�N;�gp���lTa����K�)�x߽O�W��%]�ö������Ov�I����p�Q�:bk�['�5�Gt :�������ʗ�>��wm,8�x��`"p�[�.Y�i����]	=� �kΗ}���u���W�L�T-�dz��wT�jw�?i�Ľ��� ��e��c*�_ ]al�*�N>��=fzC�.���B�_n#�t?�.|9���=�{=.vsV=��=(�b��QUd`�'���Px y�>UT�o�hѰ�a8�h���%�ao;88GP�."�*.��UQ���L�#&�0B�+�Vd�$
I#$�(���QEUQb��a"�@4�bJ6	:kd����/���3"2M��pKJ�iQD��\4�d�˄5e	48j��%\��4GV��`�����ʆ�@���6�ha�(Q',�;��@X���BmRsf��Lu
h�|�Z�x�v�~{�΢;ɺM�8����?�n�L)B.x�z��C���X���*��'4�U���T�v�>H��H�*��_݆"Gp�y�~���p�:�$o	o0�\��A�����=i�Ϊ����Mĺ��l��=i�(�y�\�I��d$�L�_��x�K=��<���H'�&sĦh��j���~���C�LuCܪZP�Z$K�	��Ŋ1X�X�ňŀ��QX
)*��PX1�"ȱC�IPY�Ě�=����"�����*���R>��Y���.
���a-��RD@�H�E�x��8繀�o6��O4wF�����%LjUO�E;OcIeFԖޙEe�0 ,��&�sJ�b���̓p�f��G�>H����*��M~�>\�F�����8��PA��N9N���}���pUGC�
������؉찮��<:s�,dKd��	�U���F �;��Q!s���áU+�	�q
�(�3)T	�CH"��l�-��Eh$l��� ���_�V
3,�(?�-�,��t�d��(���!�)�`?1� �X�+q��X"�b�:v+ש��"���>��u��s��8���x0$��,��d+H.`��y�su��%P��S�a�5�yU��i=�,ey�<e�q�������'A����ߖ�YJ������@��o�o�Lo��m�45�,�j����6�}�$��3[�2 $Je-�E�ً�W���A�������}��� \��[`T6�0)�o!]ȃ�gc��PvQ3 _	�6�H��s�\�O���:y&�V�I��]��BA��^�