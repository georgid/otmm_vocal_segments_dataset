BZh91AY&SYM�`�U_�pp���f� ����al����u@`* )   H�$ � �( �|         z� ��()@   ��@
H�JPU PUP��@

 J�TR�T�       `P�P   �R��ҙ>�\Y֞{�^�vR��(�N���}<�l�\N�o�(	nR�zt��|֋��j�W9�V����{ml��w���ݖƷ��W�w��W< w�m�yu�cW��OJ��X�TZ�qژB�T� �P @w8�ܽi��h>jr��wO,�k�=�ʼx 7B���Z��W}��y��A9����> =��#9���[[^Z�����}�{���W�x ;ԫ��W���ֽ�z�Z�Z�^8Mԫ�Թ5��ͩ^�&�x�   @  
P�q�P>}��[�wKŏ{t�Һr�K� k]�U�}i^�u}�95_N\�_8��V/\�;��}�_N]*|�� y�N�׭+�R����r�J���X��N���e�n�2j��<  � c$=�)��}�)�Z���n-J����J�<T��}���ԫ��K� �]�uKu�� F��VMR�����}595T�J4��(*�����eqg�O��W�!��  �@  31T�)bԧv����Η��Ҟq@�䫹��w7#qiS&�x� �Jd�.��� �-+�ũO8 .�.�w�.3]i�nU�{�ʜp s�]�ʦM}iɥ���7J}�*    T�'�S�JT� 2h    ��	T��F�L��10�=Cj4"x�U*�=J���d bd hh ��U)&�z� �h  �@ ��MM�)U10 �0& �� JTjyI�542jhh�i�f��#�?'��ߊ_����~��=�O~`B@ _�
� A � � ��\�� O����l�( ��X�� _���
� o���  �����A���?�7	K�BP��?��a����S�Oc���t�V��t�^m��e��gܡ����v{ў�L�Ƽ���y˧Ѽ��v��N���Dsk�2��u]u1�8[TJ����PDɎ�b��-�^÷�e���ى>`�ڪT1���
:C)Z0�Q��VLɇ}x5w���+�[~��e>�5mR��x^����Ch�U9���/K16�#�4T���s�»��z����g��c
 ��1T��^*>��������^��]��[��ǎ]�n�r��e1��E
��sFQ�FT�52��aJ=1����Q��N"ڃ�mswu�o��K���	)Bw	�'�^&I���Wi���� 2�")����r%��zmkLyݎA��������Pg0�2��U��tK�"�TVK�X�Æá��,da/#5iJ5R�-l/Y*�PS�&�q���i�I�k��i���ʪ�T]sV��9/y3����s�Yu�����^-�R���P�yD|s��e��t��T�s/��]�
���(��{���|�#�k	Ɗ!wY��������x�3o{����Np�(�Wy�q��N,��tQ�Wy*w�vI}�0YQ\�̾����V�2��*R\�{ί;ߙl�5<\��(J��9;M�������U��a�c��t��Q=fo��{��$1�c�ִ�A�d%m���5A���2d�:�i��"w:�!)���2�,��X'!(���9!���r���NI��hh�2;8��h�*!��1F(�Mp�4�#��;<vd�h�����G16��0��W�h�u}�qZ�f1b�鴩�%�]���.�+��j��+�w�k4�N��a�p��'O4��+	zs��U�1��,��X�W�F��N�^j����-0�k�bt�t'(oM��E�T5P�xYhlk����	���<��(M�P���'P��Bd%	BP�&Bd%	JP�%	��	���Z�7t���A�m�xh�Z���_C��=��<�7�Ǐ]�uR�P�^�c���0��^��G0T���;{^.����w-1�%�2����d|8��7�F+�ǃf��Y��
5�j)��!��lCі��D�l�0�s�Q���^�2���N1T~�ќ��<�h�����6-}�[͘`��=t!�P[���S؎1�}��𵧎�,4#J��Dh+ZX#�MBV��N�C���dC�PHk�㓥�J��Gl��4Op���	�By���Bw��O$�d%��12�`m���ɽHf䓹��P��N�I��F���c��{�.OM��z]�r3��
l�p�9��x{x�q�.��^�����h^	@a�"�-�ܥa����<�1�DҵMb4�0�´���A^%Z��o�w����#��+z��[:�ePB�^�Tg@��kl����<�F�K����:��h*��FS4�QuLL��CW�8UQ�28�	��8��
*�ilCaA.<�k��^����*!��ukw볘� �����aAQ*�ʳNl�N�1T@�7 �8Z�P�|�}v3�4}4���5E��J1�k�O��3ˉ��g�r��wг�s.��Le�%���;\
h*�a���I���U{h%��2�e��d�yW�_�2�u���p�,�S�*2���%Pގq�9GW���U�oN�ՙL�x��o��t��h�7L)��ASVZ%Ev^��Ѣ�k5L��]��%iU�tp-�RŬ:��0��D�L��=�a�J6���ee��糙\�<�4B;3iΘ��ݎ��Z�D��o��Mgz{��-:�(���һλ�o;͆��:b��8�F"�t��3K����e��C�[�h��?�9���E�ڢYV^l�u�]W3й�����9�r���C�T�o���%	�`�%:\���(J��2y�Ȝ8Q˓�O>B��(�"��|�Oy�nCH���Z�Ej��Q}�ft��g��7]���w�q��y�wJ4-����;5��FA��'����qq���(����U�:�3��0�pd���ӗ�=�4d�xT��R~�
5�P�G��M���%)BP�#�G������FQ���UJ�)>w�qGwܦn�����ax�"�bi�h`qh�k�8>N��i7�8t�v��t��p��){r�S0��ň�n�J5IS��z�-��B�h�M�Ƚ��mZjK.�V3���j�[TL��g��Yct�-ڳ�'����}��r��-�YamS-�oI��㌨Z�4�Q��F<�`:r�Va��hղ��o�+�:�Y�w�_�8X 8��[U�^9&���p���]кAT�I��gK�ǹ�[�t�x��4�2�ml�*8��6iSQ�g7����sN�l[5:�-[a� :�����C��s�]Cv@U/,��0{�\���r��=���7	BP��P������4��AZ3Y(sB�u��6x��.�c;Y�-`��d3q��`Q�Pva�c8�2�Ӗ�Eǅ%�@Ի��Np��=O�f���>�tcE2�����M�
85R�y�k�c�(���Q"�3Kn�����r��W.0�v��:n��}���2��Ge>u�Ow��n��|�uV��%ڋ���.����t��V:/"ф��)D6jLc�qu��ȸ�e��u���hè�C�r2u�۰ltVJ��㳦9�5p�/9�g)�9g%V�U��1��c
b;)Y�yG%f]�T`Z���R�ʙ�Z��YW�n��cuq�i��U�h�Ud���w sk��
�m*E��yk���Ѻ��*eT���"�YK��V5�=%�1ǚn��K�{3`��V���B)�y�lDh�23FJ�r�{�]�9É��8�R:O��M�\��K�U�}����蘱f��h-b�Cb٫F�5�K�I��A�	I��'!2d'Y�P���' �|����3QjѰ�n41��b	K��	@a���d%8�E��	w��c�a4�V�����1��;�۽W!�a�TH�H��u�S�cn���]gL���ܲ����:̢'nX�E��e�����,�v�u-�є�#�wu�5P���nЌTɌ� �-wk:���]Y�j�� �!��lCb�@��3p�}4�Tv�T ��f�a���
-��f]˧�uw���ݪ���]h)p-氬�U��F���gl�q�����N��	��v:��	BP�	Br�JR��):j<cM2EI���P`�&'E�l��|�Z'*�aI�V�
��
�Nܸ������x�,te��7]�UY��_�i��I�2٣&a8�[v��{m��jS�L��;��(J!(MJP�	I�۩12qrL
��%ݏ�ڠm�:51���,��[��݉�J��2����(J��J��(L��(J!(J��(J��(J��J��(J$P4P�%	@ua�	BW`Y�BR�a���JeKL�,`QL)�����n���3B���emov�P$�q��vKU/e�s�̐1��H���[�+r��2ƫ�z55]}�zᴨ���B�����p3NwF!�J��:lC`QT��B�8-��o
;��R}�y����F!�%	BP��	BP�%	Bd%	Bu)BP���(J��(JS!2��2��&�(JR��(JP���M�n��7	BP�	BP�&BnR��%	Bd%	Bj��2�ް���eM(�����l8J�q�g�#����&��T�Pū��Y�<��z`j�Z5�b�z��,�K�X�YŸ�Y���J�,5_;�)�-����g[Dt���o9ӧ] ��^;*�Ù�O�i��F*u@��Dh8ꈛ�o����;*碾5���׹�qԹyX0��EAc%����v����)��q�j����m�h�\ì.Ѯe�DB5@����D2y�l���P/;�
3'�S����ղ�T鱘�E a�a�Q�ɜ�ԙ���Q�+4��B���ƈ���+9�1f�i�U��(3���nꕉ�lu6<ʭ�#���s�oi��n�����kٹ&g6���0������X��6�"�R˿f���+��;�펶V5ԩ�lCb(J��J��(��ty�u�k�}�V���œLx���c�5];F�U�V��l].��e(؆�i4`C�&��1��
����[N��4�LNfG8�t��HfI���:2�N��%���ۨJ����%�a	c����y��_��s~�vl��    �       mh                           ��  � �|      �       	 6��                                                                                  |��                                                                                                 �                                                                             ��                                                                   R�����>    8��   �` l:�BBI-��Sm��@m� m�m���m�p[@�$	 $�-�ЖPp {M�:�Z�V� HH�  -�  �kXӉ6� -� ڲ�`  $�K.��+s�̭HpJ�A�;U w[@    ���FP.-m'�q��E�(�l����@V������!��q|�R��R�ʻ*f`*����9���H p$�܎����` ^I[n���\ 4�l�צ@/Z�l�r���X�W4j,�b��Q�N%��m�[u*ҭtd)���x�
NM'�=[���&Z����9	�2��cF®�NV�H ��k\��&�WU3i�5 r�P�!��1!Ut�e[�n�*���m�fy{k�n�C�n�m+��{�v1�jK�����C�%��LU��� $r��gK�_�Ŵ^��Á�U��Ѣ�������&�YoS��j�^\Ӟ��[�b���6�ݪ�T�gD�֥ʺ���8{qT\P!uD��0�tݰ`�^�ҹT�.��Wg�C�����]�f�u�r�헭 e�iتM�:E�m�j�]�&�3e3�-v��LTu+��;]*�uT�UN���l�@m: +�U�S%V��P.ю�U��;폻�we���A�,��[��$����w  �H-��e��n�k�Ĝ���b�ŲW$ 	m�o4[&r� �:��	���������( ��� ,�ڐ�8��'a$���9�ɠ�66ڶ�hr��#�X˦�k +�,��Qns�:� d :  d   m�3�   9��     '     �l    
P[rA��  A�    �M� (0 8��  ��� �p� �� ��N� �  d  m(-�1 p ���� )@A��: d �� 2 R���r���       '    ��    9��p�R���� )@A����� �p �@
P`8[@ ��     �           i�-'8�����mm��	����T�B�Ġ�m�S�❕�7g( Ռ������NӶ�6��&�D��v��E��j8%�v�����&F�m� i6 -�Z���6���	������L٦��X�ۄ��qf��p6ݒ  m� ���Q��`     k��T ڮ��V����Y"1� [Kh��l  $��͖��t������/5m�A�T���@nlҪ���m���Bz����à�ڪ�*���]�v��UPlA�J��[� V� ���[�m��v��Eg�
s���&-�bѺH!�3����ۍ�S �:0��g8I����+���3��A�[UUrZm�9J-�������!U�.�J��v��*���[;  �RP���G.��`����巒�v��v��xC�LTɹ�kl��l�J��mB`$a�;.ߗ_}�@,T���<�b��}�]��[@m ��v̀���|���&�ܬl+��KUJ�Ö��U����
U�Q��W`Ht�[m�Kh���pd���dQ���;�@�֮Z��8l�8
�ȸ������Y\�R��v���/GaVhO�||�|+@Xn4���[E���6��
�clT��r�yj����Uˍ�r"��U���qu =�`�꥚�n�5���i� ��H��i��ŧN��Y-	�@k�j۩��viW�UZ�UM�E���v3D�À�����ۻwm���,WA�p�J�Uj�4;J؈ߤ��Y�USʁT�xnv"g������d�j����55J�9�i��<�����U r��v�H��J�8�%$[��kf�]5\�; C�9�`I͖�����m���U��U;	xv�駕�gu�.�;���I[��ڹ��82U���Q�ֹzr�pqj�h`�F5<�ܨlr]T�q�=ny-�J�t,媮�b�m�a�j�&AvG�6׉UV��x�p[�v���1�ʎV�͕�8��5+$�t��[�t�;i ���&U�dl���T���U�+�L�2Kn�hՕkmHuU ��E�5[),�����Z��]����Uv�|�x�V��;�m�m�L��&nӲ
�u��!����$��c�	�K�)U&�	7k� -��n޻hw��i�Mۀ[��ą�4������@w`���L�WV(Cce%ѪW���uÝ��V��'K�)[Um����)�^8;	ݺ�q�g2�*���R�і�ߘ���%z��É�m��5�pgd%Z��VۋÊ���:��T�wVӂ�j�&��JM��s�7�ʺc5UTj�Wv��KC���l-�<{l��W��=�X�Vx�xg��vj�m����U�̼n�9rg���I�Y#�����'L���5����� 5�P ��Z����t�l��$�����4Y-+�s�� Y��������,��-�2�6G6ۀm��;shÇ�    �vk�6�sc#Ֆ	Z�jڎj � h��lWV����p  �:޹� �`��im� ��@�  � m  �mK)WK��H��-��F� � ���Vm�v��8-�6�i6      m��k�Z�5R�F�l�.љ^` 'ϟ>>   HH$�  H���p���8$m 8�kn  �Hm[ 6� ��T���R��@(@ � �      � H���� 8���&���k�� 6ҵU@PAdL�r�uP�     m�m��a����kZ�m�m� p ٥� �m�`�����m1,���>mU/&Gd��^j��m��,�J��  ����� ��6�s��!!"�m�v m�$���l�2ut��,�l9�l�6�0����͛`[\[RH�z܆�HHm�j%�%�m�'J4����p6�K0��I5�፶ @xcYU��m�o!^��M�!��H�o-(�jZ����\6XX�C�wBem�ڽUWV��rKuK$�mX�$���ri��+��t�v�t ��Z�Հ�&���:@=%͕h ^y嶧��\heGggj�6���ɱ�K�UUT'�K���}W�G��S���,�UZ����[�.���@5�I��v�4UvqJp4	�T���qm��	Щ�Y`8mׇ���
� ���/X®ƭ�������'�J�-���[����#����q�1#�m��t��Қ���]�:��}�v�e��i��:v�6U�S˶F' �u�`p�m[mYe^��wq�Yi�\Ē-ce��A�mK�$��v��h��}}�|�|�;�-�(+�E�l*��v���c;d�p��Π �� ķ� ����l�'+�Hk�6�l5���*�4��*�T�k".� �Km�֒m����S$�~��ԁ�O��5U@�WT�M�d�	n�]��\^�T�D�zM#�9m	l�u��H���m�k$sr[@H�M�S$u�&ڶs:S�.ٔ�O���EO��݈���ޗ���(�/�?�������O��
�����@�W�EE
== 0�h�
`�(�
' N���Uv�?�@>
�EH���i"���)����(�&` bT��`HH	a$!`dbb� Id`�Yad��
��!`���&�%&X�B��j$h� ��I% i�!I]��ڊ.��G�A^�� M�N��(�f��`*$� �� &�f&�(V�����( �	Iba�&Y	hRa��v�Ђ��o�Ъb���0��� 1S	 �zE�T8m�P4!ꠞ�TpD�B!�N�S�<UC�Cb���&(8�i�Q t!�@ CJ��l ����P}A��i���
YF�)��D!lS����J�v��J�@<<zv�. ؂)�xiVU�"� �ࡊ�g9� v��x!��b�@=Pk�}v��?����A@ ?���������?�s��X�bP)d*AfAE���a�`%���ZA�@�A�A�A���(J��"��(J��!�(J!(J��(J��(H��(J��(J��"��(JB���(H��(J��(J��"��(J��(J��J��(J��(J!(J�(J!(J��(J��(H��(J��(J��"��(J��(J��J��(J��(J!(J��(J��(H��((hhhhhh��(J�J��)D$�ZJ����c  m�    lm%l  m�   6�            5�      	         H  ��              l             m�m�
���s��*� ��n`C`��5R�����<bI�ȵ[\q�'m[�\Y��j�IP6�6���+�2<����2�n�3�q�l����F�Q�ȫ�嘽+D��Ku���h�<$�m��m�1�s�Y�{d������^�,��Tc��O)�������I�3�H�wgf6��ٍ��1-m 	�E ͮ ,�����m'@R���8p 	� -���qm �J-��[@  5��eX�u2C����#v֎Y�c�9�@uY%�Wl�l�P �N�{\� ;��&��]�e�D\�Qc��8�Fv��G�mҳ�8�g���+a�2���a�7v�����Ī�\�P�� ��1�E���n=��@B�;���u�Y�f933��qs�l�m�����d�6�XT���@ڣk��]�wǳ�;���;ʻo�΃�	�����6�6.��N������D"�۞� nI�9�+Sҍ��62�m\	����\\���Юz�u�Wnn\퇉�I�y3\�z�vtƹ�ѓ����/���٘����-��U[�.5,[� sM���ev�[�LQ3�����#�rM�vU�@ xsf[.[c�������ʝ�]
�f��S�������_[����ŶH�7n��G<��e�L:�4r��

۞��N3�S\�3��6p��rgs�E��Ѫz{uP�d6�tr�7[,��UAt�̦�X��Z�'���\�qE�e�a�(3�Rի�����@%��(f�랹6��D���f�ٲַ�P6
���e� ?�TP�� �	���|���9~���l۳l   8 �m�  m� "����\���v�Y�k�n#�30	z��n�`��غe���8%�Q��]�7�.+�%��l�Kb�u���˛�O�g�L��D�����vi&e��:S���V�uZ;s�ЦS��8�E*��Zٱb�ew2���t��<�b��;qs�qr1�߽�{������*��Cr�;nrxS�2����_p�;���m�r4!*��{7;]��@-_�u�>Y�}=�� EB'��C����]��UG@��U�3�|$L��"�9�cr.�������c��gk�^<��>��
�d�2F��t/j���%���)�}��;�ɺ�lDdq9@��;]��.��ޕ�@������ci4�rI E�.��s�v���d���p�Mð��b�1)&j�]�B�7�)+�^<��>�Ұ�^�>�fv�/y�a�%*���|�l��IQ����|ｆ6��غ���$��AG)���t/���3�=��Γ�����ꙥv�(��'@��;]��@��Jày}�}=�� EB'��C��*�=��g�U�3���� �UUF
Ƃ���c7rX��WHl-�����S���ڰM�Dޑ3Us�>�m�6~�]>K��1V��|��P�q�#RB�����/���@�~��>��
�_{ ���Q�r们m�=�1����c�)�����tǙ(�
��B$�����s�?;Nz�G@߫T��.�@��7�#C�Q$�Q���>�Ұ���@��;]��@/�F<i4��@������ʳi�@sd�gD��crr%qg4��a�#UV�	�R����oժz|�c�b�S�>�n�ꙥq�P:��Ɠ��_ٝ��x���}��a�=��.���u�"���r!�]j����p����r"ej�t���@ό�u�s�&��]�+��~x��v�� �&4� J��V6_��P� �'R5%C�{�L:��@�~��/�Jà�m���%Z%;eM�;v��-ZnM��ձyl�sz8�4p��j�L���Lվ�~~�������O@϶�~�G@J��.�&�B%$:����:��à_ޘt^�x�4: I)Sb�����7�t�m�:�j���#�(�FԂu��0������~��:/bO$d��(q���3v��>k��>J�~�G@�ۿ [xp8  $ $ �      +j�zݦ#\��B��=���/���NT�H��kv8�����Đ��E�zJ,����Ei烑ёnۥ�N��rt���+v���K��@�6��,���Z��:^�M��ç3Ε�g��o;[9iӅl���.ͳ�y=]��vtW)�<ܖ2j�w6�M�����'n���ߞ��A���
Ʈ:�ֿ�����1\������w+�ѻ�	�g[DU�IȈ�`}�4��L+�{�L:������p*$� �&���h����Dȵ[:�[:J�]>�aC�l�mH㐮��0��L:��>�~��:���(�t�JR�%�ݝ7m%j��������:y�J$B�B%$:��}��t��N�~�à]*>�i4��I��bg�V�UI�XΓu�A=�N��Z�����7�%v����ki��O�o����g@=�d��L:��} ���G"�]U�.J���������&�bVaDL�2���H�N�$0 0e��� ����:����/ޘt_bO$d�P�4���L:��}��@=�d��βQTj�q(��-bU�3v���W�3v���D��¢NT)0nE�/ޘt��N�~�àZ���=���n6�IU%*��
n��mڷ-�D6�wY��S�=�@���ƫa�6N6�q�t��N�~�àZ���/ޘt/{ ��ӥ)Jd�rN�������������n꾀���$B�7 ��@����Z����W9WʧT����=�0����Ht@����}׽����t���f>�_��#�G"Qʌr&������@����Z����D�MUU \�:�y�����F�-������ӓG<�V�#�
�Wl�;7#_m�?��t��t��O��I�@m>�(�U��J8tǘ��{@=�d��L:|f�����Q0NE�2wUtwU�ݴtT���� � �'R7$} ����_�0���V7Ą"�rv�1���}n�\�*ʔ����@�y��Z�������m�?]��܂UUW������qZ�-�����G����'k�M��f�j�vM��"RC�^<��-{���{'@�za�1{�#���)Sd�t[�����n�:*Jz�j�����J9Q�D�} ����_�0��1t^�>���I䌒�ƕ')�'C�$�s�Ϟ6�������{���
�{6t�޲Q�	ECq(��/b�;�����n�: �������p  p� ��    *��-�ݺ�,�A�v7sl@Y��n]�ۓ�e��Z�v�&5�p�mt��f��L�K֙�jݷ\����v��f��@kݮ�7=v���<�nm��lc<X���3�����W3L����wӞ��Ď5=vt�:,���v1�m��n���:q��qw��{V;r������ki���m�:�o.�krK:<��^�����X���Β�t9W��vˉm���e����?i�@7u_@��G@�IO@ϫPpt�R7$} �������$}�4�k�]׽��y{�n�)JS$#�tݴtT����] ��}m%t��B%$:�����>Y���{'@�za�1{�#���Q6]\���] ߵ_@��G@�Z��o�������nx��F�㞣��;��iR�qaq�l�ԝ�\�f���Q�D�} ����/ޘt��]׽��b�)䌒��eSNN�~�ü� H�鞬m��Lm��m��βQ�	ECq(��/�t^�>�{�d��L:|f������aUW='uW@7�W�3v��1V��|?`P'Jq�#rG�}���@�~��-{������&��I$�s�{����cѵ&�1Q׭�+�Q��:5�g�7.��AG�JR�����@�~��-{��ｓ�g�d���&�rI���:*�='uW@7�W�3v��UUčY�c���$)Sdqt�f�m��m��'Eqcuht�V���K��X��&ʰl�l33�'4����M��@]BD赫0�9��6XZuF��F��J3�sֲ�fb��m�[������0�L�ф3����%�V�2�;�Y	j�j���u,.��,Ѡ���#-e��M��0�fj8�p�(�����l�再IHWBַ�*�����18��4j`a&h�Ɋ6$�F����9�(h8tc�P��0���$&$�D��QCDC��-Oy��@Zf�]h�j����e%QJ� ��$:�4`Hh�t#��f%�=�l��,9�X��&!6�����1���a,p+.�:۵��3\������ v�P�E@z�iS�v��!"��v�8����F��3���O��Vzn���+��"��R�٪GnD�Yq˺��Z)��)��]��5���rN���\��rL�����ԝCM�M�����M����O�����21�&Kɍ�M�M���֊b��h���4k4S4r{�L��rL�=�=�\��rL�$�==��6Ͱ �ۤ��]�e���כ���9_n9n��ܹW�nJuڷX#��;�=I��'o߹�:�$�rN��k�ԙ)I�����)w)Jy���w���(9[�t_��Q'9��;\��H�{�LHm!�w��}�!��{��┥'^����)O<���kef�ڕWr]�Ć�G}]��Z�H�>)JRu�����R��=��qJR��ﾷW.Be\eۼ��-i�s޿�)JRu�}��R��=��qJC�P�10
�G��=^���9_y��!&�T$s��Ch�w�Z��k��֐��ﾀ�~�Nr����ci4�rI E��Y���1���n�ϧ,gVt�dշdD�0-0d��o{�5�7�Ҕ�y�k�R����{���JS�}���˒�����ܮY�Ps�{7�F7���M��r���9�ﾂ֐�G=�Hm����JS��ߵ�)JO����{�\�
�#�d��֐�G=�Hm����JS��ߵ�)JN��=�Cԥ<��޲Q!PJ*�I;�Ps���n�z��;�}�\R�����ߴ=JR�ٛ���+>3���'8���:=JR����)JQ�	������)O>��8�)I׿{��JS�M��{�ӽ:{��{�~o�`96��  �� ��     ��@{q;\��%e��:�4y��xV�9��n�p���9XY�
�Dq�����T�&�}[S=�c%v� �H!z������M��w����x�J�MFݺ�ZSӎq$v�Ē�Y8z�X�z��m��O[�"�br3��fA��5�!k���R���IתPG���Yq��w����w{޵��9�A�����Z�=�/FԚF�6�mL��f��^[�W'iR�H�	Ҕ�Hܑ�9A�Pr��=����JS�}���):��~��)�|�5����(9Y�͂�6�JQ�!yy�Z�H�<Hm!�o���-i�y�k�R��{�{���JS����@��P�RC��9Aʼ���,��9]��Hm�w�AkHm#�����Ps���ǱćJ:$�*l�v�b�'���k�R��{�{���JS�'��Hm!�o���-i�?��]�\����T���6����6�'�w��┥'~���JS��߻��{�'{���t����@Wv�K��<$nrxi���;79���r�`{[s�4y�r�0ňs	��ZCi��ՉR��~��R��y�k�R��{�{��g9A�V�oY(��
7R.�JRu�����?�i��0"����,����)�}��┥'_g�~��)Jw��8��Q3�����
"s�Ls��9�r��>�JRy�y���)N�׿g�)/77��9�r����t�16�|R�����ߴ=JR���~�)JRo������9]��Hm�}���rF�ʸ˷y��Z�H�g��Hm!�o������9]��Hm�{�Ak�(9�=��M8ܒH 0M��]��s�v��u����a���V�{ۙC�Vj�Vk7F���oy�)JN���=JR�����6�z��6���}X��9A��}W�ߵ��$:Q�$)Sdr��R�g�~� � ����}�}�Cԥ)���qJR�����R��������Q�Hԧ�8��Ps�����\���H�g��HmbI(���1��_���R��<��qJR��~�5����8V�j-sW7�hz��ʋ	���qJR��߾���R��<��qJ��d�}���r�r���ۿ��D�J(N$�]�
R�����R��y�k�R������Z�H�g��Hm!�oݯ��r�U5UT`n"C�=3w%���%t�b�����Nڷ,X��Vڱ-�ho8vZ����H�{�LHm!�{��}�!��z{�┥'_}���)O<���kef��*�仹��6�z��6��O}�R������ԥ)�{��┥#����W.H�YrQwu���!��z{�qJR�����R��y�k�R���^�u�9�r�즠�&�T$��┥'_}���)N��~��)=�<��R�*����8�)I{�����GQHS��'k�s��|�7\R�����ߴ=JR���~�)JW*�۽�Y�Ps���F�i4��I$�('�{]��Vn�jc�&���Z�Uֱg�{\��ah�6$ڡ3�]���{�'����=�Cԥ)ߺ��┥'_y���&�������Ch��?�r�0ňs#˼�֐�G==�bCi�~��`��R����)JR{�{�����Ò��}���[�l�qf����qJR���~���R��=��qJ�d�{�}�Cԥ)����qJR���}��kt[�m�Q�wx-i�r��$6��=�����JS�u���(O��'����ԥ-f �t�17$}�(9�Vyg�hz��;�^��R����~��ԥ<��f���+����Od��$�N ���	 	 ��     ��A�:�kD��z]��֮��-��3�tf�6���n��	�r���Q����\ş[i�	K�]p�뱇J����`*,�5ٺdx�F���.M��.�dʥ�m������]�ۆ^�ڈ� 5�6�c��ڶ���K��&Qŵx3�ː��׮:s@��}����#;|��+UZ!8�#��ĝ�pE��+��tlVӹm�<�n�;��%f�J�ׅ�>|�����Ox�����R����~��ԥ)�{����Pr��3]r�r���ǻ)�p*n��bCi�~��`��6�������)=�=��R��~�߳�R��}�}w�\.��	�൤6������JR{�{���?�$d��k���)�+�߿~�r�r���}�7 "0���6�z��6��O}X��):����)Jw�����)I��^��r�0ň����AkHm#����"������ԥ)�{��┥'��f���9_kX���i9$�IJAՎ���nwifL3�@���D@�/'6��'�Bq%"�9A�Pr�ww��8��9^��Hm�{�AkHm#���w���(9[�-n9�&���JS��ߵ�<U��	8��6��+��(�,�	,�+���������)Ok���)JN�w{\����+�hP'Jq�#rG�%)I��hz��;�^��R�����ZCi�{��6�{���\�#ue�E��^d���9��Hm����!��W��Ć�G�]��ZҠ�+q��j�
d��y�r������kHm#��}1!����W}���r�ǚ��Ps���=��i9$�Ia;/g�sf���,n{s����td+�vMwn����R�;<OEnyt�w�7��{��?~��)JR{�y���)N�׿g��{���Y�Ps�o�F�A��I����)JO}�=�C�~d2Sϵ��┥'�}��ԥ)�{��┥'���O�����22VG�y�!��z{�qJR�����R|Tz]��=��┥'}����R���~歖��۩uU.�!��ѿ}�Z�H�{�k�R����{���JS�u���)H�o�`��D��6�k�s��|�>��(��$��{��r������Ć�F����kHm#�O���K��UQ��Ì�Flv��rK�d�o!�H�zn�.� qMƫd����)j~��o{�G�]��Z�H�g��Hm!�o���-i�r���Hm�}���rF�˒�����-i�{��V$6��7���R��y��k�R����{���JS�^즠*P)�&�]�(9�U�����JS��ߵ�)JN��=�Cԥ)�j�9A�Pr�s�:RJR)���)@��{���)Iߙ�hz��=�^��R��ő����i�"� �I�d��߾��)O(�f�����$�7y�r������ZChG�=�bCi�y��kHr�[���Ps����m&��I$�	��ם������U['[U��Kv�M眫)�BU�'��2\���#%dyw�Z�H�g��Hm!�o=��-i�r����R��3�~��)J}��sV�f�yj����o8�)I�~���S��ߵ�)JN��=�Cԥ)���ഥ'�y��j�CRq����r�r������	�����-i�{��V$6��7����,�(9����4�1:S�G�>�	�����-i�{��V$6��7������9_{��6�w���[�)�f��7��7�hz��=�^��R��� Iߟ�~��)Jy����)JRy�y���)N��yCz���f��[3d5���L�܈��[��bƩ���e�I��*�X'R�̸�z���`��F!�,����C��U���ԫYn�n����Q
[���*��t�v�4�[K#�Ȥ�\�H'�G,�rTN��iQ:��`4<���HA`�Y�ְp�[�H^`9��"$d�鉌ì��A�da8fbY����1L�5pq��0x�}/l�����la�q����a�):4�!���,B�X[h9�X�Ř���Iw��61Yy)�i�o#��a���ԀOJv�9�Cp� �f�-<�N�TmԪzں ����6!���^z���-e��CYE��Kݧ^�;���~w~5��p  �`     ��  �v�  �       ��   ��      �        �                                ؀��}�X�(Jf�
Zڪ�^z-`6�^�($��R�n{V�jG�#.nB�Z�J`v�����:�s�����{5�g^H�us<C��Os�ez6dCV'Jm��6�k�q-��G#�m�+�v�=���xƌ�,�<��&�ku˩1#F���Xk���W��\�@�F���yv���}o��}�TKV�hmp��8 �,����e� ����d �� �a������ 8���  Z�kt%����g�VX�.oj���:��de�ed�ҁ�]�����b�ѶC�F�uu)�m<�nؼ��vse{z�wOc�����z��!��[��5�u�s�s���uM��&u�Z�+�Eiu]b�W�������Z�q���M���cp�V�-u�J����q�N;�+�5@W,�a�mn8�sŏ]�����L��v�랗�km�r�k�a��\����l�se��Z�ct��ͷ=<�s��g`��mŲJ��P�n a�К�㬊����ܝ���� �ݬ��O1�:3�$9�1����H���YՕq���y��B�Z��k,k�,�P8;\��/�������в�Tnz42ά��e �v�fê�غ�8�ٮ�s-�,Ut����5���#L��t��� W�� -0�WJɂ[mLV�)J�ݱ��q,֬��㰍�m^L�s�uD�-�����{���{�ܼk#�-��V���u�u�n��0ȶ�����b��r1��M�t��F�qL'�����&���/H��v��|�}���9����������o7�6o7���<TC��	� =CG�(= z��~V#A$h$�@�]�N�.��꨻���  	 	 m     P&�'fѣ���r��ٺ�v)�O!�;��h�?���;�
�gb%`��b��UE��H�i砶�f��zHwR��g8��릋\�{G`nѳی�h0n9�8θ�#��f�Zㇴc�7\�\e��ki���KW�mKʬ֓�=�]׺�\5%�hr�=�]�N�s[v<��{���{�Gk����U��i���H�vB�76-&�0�u۲�׶�q��Z�-��[s�Z?�{��R?y��R��y��k�R��y�{��֐�G����Ci���>��®쫶Y%U�ZCi�����G{]��R���{��)JRu��}��R�Q��i�$�$M��r����{��hz��=���qJ�����R�H�}�$6��>���\���#%f�o|��)H���┥']����)N��~��i<�<��R���{�4@�aR����y�r��{���,�r���Hm�w�AkHm#����r����{05썸�m�$�R��"���7E�.�rޞ�gv0]�P��nj���z��ݤ�9���on��o{��JS��ߵ�)JO<�}�Cԥ)���R��y��r�g9A�W�=ѥ)�Ҝj8ԑ����Ry�{���bt;d�`0K0# ��$�	����F�i ���~�<6p�Y��&886bf(�d5�ɒa�����hM�B=�}����r�<�>��w���H$߬�*�B�.�b��/���~:jo0�@}-:�y�k�7즠*P)�'$:UFjo0��]�`�[:iS�:RJR)��幯�}癮��dӠ_�v����i4��I$"�K`��<s�t��p�/R�K��<uG9cu�n�;�F�I>�� �dD�7@��7^ �[:ڛ�Dr#����?W@�f��#/����S]ggz��M;U@}�o0��]��`��.
�.Ku%�m�����+�}1���B������ ]kz���uW�}��*��3�-P(i����a�������@�=������PG""u7ށ�SeL�Q58�q�#�/{@�s����~�۰>[�����li4��I$����7��y��mI�L5����;���p�x��F�g�i�Yƨr�j���z��M:�7n��ju�G"?A�T߫ �z��Bj�"����:jo0�Dr#�s�&ϟ��y������=��?(2�	����k�p)%)���_���y�k��Ds������'�f -N��ɘ���ռ��浽r�(��0AeT�DȤ���X����3Sy�<�9|�sx��$"�J�_��\���[O��*WYMu�����<��?Ur�,)�I߿~����?}�\��5�k�I����ߡ�m���-��\�aڹ�9���n��q�c'-�:+.U�n���v�v�.	�&j�f�� �Zu�>�Iע �`����_~�U��s�Y�7E���Y��z�����~�? K!W��~��~������D�9��"D����)�Ҝj8ԑ�ǻ��皺�7n��nk��f�A���#U!.w� �s�i9����>��t<DG'U7�`~����� M���t�n݁�#����tT߫ [I�@��;��8�6�� � � ~��    [ZԒs��.�ɥP{��:ܽ����^Qڞú��%��tW%T���檭�j�@V�P��T��1�	���J%c���]�N��x^w�����:s��J;{X��psn8�q����Q6����8d8�y�����n���:5���N6���u=��qι��2]��V��\�c����U�A�3��<�{\2vG��s�3q�:wd˺�L
���WL[*W���g���>�I� ����Ȉ���ـ��� �9)FDIq���5��� Z����`KN��(�wFw��*{۾� -N�jo0�9���I����	S~���E��ArE�5pM]�#�����{��g���7i'X9U�ɧ@�yc�MIvɧ]v�u�-V΁����n�E][���2�al�����E�u۩#�q�0.C�e�5v�����c?}�����"f��n�N����3[yȎF���@��6
��"�޻=�N�s�9��"#{�^c�e�]v�u��C�J���?�5���ַF�������~���Ӯ����DD�9�Dr)�������������)$pjK�>��t�I� �[:�p� �#���?~�v���rT��dD�7@���ߵ�@?�P%eIS�~��}��~�幯�}�^��JI$�I"�ʦ��C�F�'���{Vslw:�l\�n{�����$E��R��k��v{&����u�]����~$V@�	W+1��v������DS�8&��/���u�@p��0� ��s���]���V �[:ݕD�����&fS�w���}�6�]���t���~V	FE�����o�ʼ����uW�=ѥ)��S$Q)#�*�TW9_�W�Dr8DD^��~������wa��^�������8 r�$�;��W�{��U�	R@���߿s�<�o��1{3e�f�km��m�$�#vx��Í,s�v��ţ�$�}���q�<f���	H�s��k7F��\�Wvt����>��t:��j�:�c{#JI�Q�幯��XO�2���������W�o�r������`'�HIMW�,��k�J2"H���~[���X�t�ݻ幯�o���"/�
��S]}RvX@���!��>��~�W������>��r��S1%KARL_61J4�3	%IRLHD),�C�pP�T^	�"B�f�~�o������j�[DS�8&��/wv��澁�36X�t�Z��&��I$�$�$��s��7rX��W1��ַa�k��X��V��w��bXH �o:՝f�kqfkUU_~g����N����G<@p� AH�,�!���~몽����JSD�H�RG�1{ٲ��I�?������Uw�{������*�!����s�73ATp@�HS�[�{,N�tz�`N�]N�w�5M�T�3Z6�y�o[��_��I!D�
�,�w��ߺ�3߿k�{�y�����LS3�
B�,����:�ۭ����$�I(�R]����)�N��[:6�`�aF��00�#�0��° �A����rL�hI���~'����#�l  � m�    �������KzZ��c��,�"vr/�M�lNn��s�G�sd!de���	�]T�S"�1gՊ��	m�-��#1�u�=�F�$���q^�Mø77�S-]Je��֞��e�zw-���u�u�̾|jn9�(u�r�)ۊ��gɦ��s.�V�s:�;�a�LÞ� �UUT�y�(�Z��3��t�&mn'u��BRQ
m�F��Cn,�W�p������X�D�BC��γ5��T��tJ����ş���`}�t�ͻ����74��"/�
��S]}Rs}Uߞ���$�"jIB( #�G �Dp�r(7��~�K���
V�xp�L��Ȓ����h��싂b�����:����ө�@R�w�}����%̈́U���k[�]W�S�$D)ȧ����\��~�������w��� �H��a�`	Tן�����U~����k7HM�"�I@ř�,��N�{��`|������[m��nI$"���L�S���v�"�gM��uչm�7M�8�n�����$��!� �wm�r�7,�d���{��N�tm��>�N����q��j*MԨB(�:���ʤ;|����b�)D0�a�[Z�M�,�bF�E�#4Y��Y�#4!��tkX�P�U� �0q�� �Ӛb�((J�>=�O�C$+��yך�]�}�}Uߞ��?�X$�s�?~�o�)$jIDd��,�Ϡ)I;��9��Χ~:���� ���������oz�kz�"�		N�r\��x�~:6�`~�s�����~����"�B�X���'e���iР�"���~����=���W��f��kZ�M'$�I"J8�H*�������� ���!rv�����6�N-�x��w]�*P�	�ۅ���߿]���k��3�Ŕ(�;��~��~����"�IE(�#����_yUU��W+� �Gs�s��r߽x�~:ͷ�xy�Ԥ&�L���>��3vXw���������H�\�:JU�1Ը�a4�f�*�XPI��v^�r�����w����w��:`2u�Hd� u����0ѭ$H"�λ�R ����HF��g�9��X�:�l��5��|�;��b;mh�Y�|�ml#ldlw�}f�lSL�KDy�q����.�u�ѭ8��D��47$t��EPq�nt���b� �Z2L�kF�kA69��QX����D�X�+��� F��2 ���Xf��f+���*zT^�Qx"�=�H'�E}V~E���@>T?� 	�@������{�]�o�ϠfflGT�9%����y���r�?~�����<��r���*�.}����}U��~��Y�0�ո�.˫��|�y�}:�t)7xڟg�'������[��͋��&�ٲ�7K���%n�V����k�t���ߞ����۽�&!�L�&�I�q�U�ܫ��軼���]JM���g��G9��E�Y(�	-W������P��rT����M��1{7e����x�������+��b@~ �I�&2� UU���6�HB�k���ҋ��� ���@��� �u:�
u7xi�Q���e��5�ֵ�����ID�9;��f �?O@S����G#��8 �����=�<m��W��.��]�sWWy�-���r=r!�����~:�7��Dr�D׮�ꮪ���{=;��3bMط-�JDb�o!�䋖k72ꙛ��/��W�qt��jRD�BF���K��׀|ճ�|�y�-��%��Tn�J��$���`}�4�+�����f �?O@S�����*l"i'
��C�}��vy殇*�_��՛���=�g�n{�:RHԒ��n� [I�@����5l�DG8}����蜃U!*:%9M8���vX5l�ko0����sb#�G9Í0$��@H{��ff���{�f��    6�      �f��݉��,�:�v�W`�&���p�Whۍla����D�ܵ]��Ut��Kh��p��5��������4p]v�XD���$�n��S�������-��u�X1���ʫt�^ݸe.4��l��N\�Zt�$)=� ���dK�'ڻi3�(�S1v��u�aw{�a6�j��	��ם������Uu��M���rz�l�9�+�C'��{�����ko����C����w�}����s�d�����7w�y(l�Dt	�ۇ@�ۻvr��i9�:��歝�s�����~��J%�r���ǿ�@��n��ɧ@�ۻvxy�9@�%24�]s���?z���m� ������ت7T�9%�N��ɧ@+���[}��s�6u7x�;���� �ڜĹ���a+X���4OiwM��nwa,�A�aڤ����b|�}����s�6u'|���π�;��=������$�I(�).��<����*�
9���r"�R������3[y�+��۩��I���]�ٛ,��t��r&~^�� j���6���uÏ9kY��o[����©�_�Gߺ�V�߿f����u^ ���\E�[�Y�浭ܫ�>����Ͼ�=���׀|ճ�%��]��U]U�UN�Ǣ���������u��c�ND�tf�g��*RJH8�%�r����͞�����>j��G9�s�9��f�{�(Q��9@��n����ʻ��몽�^��Ф�9^���GT�9%�w���ퟎ�~�y�c����"*��s�2V�xt��M��f������{�@�Q ;����`S���I��V΀�UNd���G�`g�j�Ur���U�r����9M��|��@�m����ku��;_:������z�y��E����s�Yѧ%t��-�ctvv���:��歝5��Ȉ�G��� �����_~�U������n��ǜ�S=��_o ��g@�m� ������}��D��(�}�߸쵫t[���UY�>^�� [I�@�ԝ�54��,�8�%�r���s�ʯ��G���
S~�歝�G"�J@�x
o��������kef�xQe�M]�@�ԝ��G9��Do�|t����`g�j��,FƓI�$�H���%4ܼ�z6��k[uɸ���h�Dn8e���pA%HS�_g{,�&���� [I�y�D��9�)�^ �^���R����C�_�v���]gRw�|ճ���s���#�{���¢n�E�r���@��3e���Ӡ_�6��ۭ7�"#�S�Ӌ�UU�U����5���Nzlu�/��w�iuv9�`}�4�s���/?g�5O��7kS����6�M�ݒ8Xc� � �      ���5�u�ޒn���v��k���ORԩ9��㎈b�1�Rw�ꚶ��F�U:%��ے�v�,g��9&�AE�v}�׫���=��D���6���vqq�j�s�GG*3Uc��wҸ�f�����7+���7�]�nڍ�k��+�՝v�F�k�m���!'AU+m���m�m�*��v8��w�vr݃����rW�ˮ�Ol0��[o�y�0�������܈�C|��@��[�#���M9J9vy殁�?f��V΁�6�s��F�~�jb	r.���;�ɧ@��v���]��ةGT�9#�����s��A�}��>�{ـ-���r9��i���w�5�(�'7�@��v��D~�5oӀ%I����tM��FZ�� Ǉ���,��<{ s!��l���Ν=��e�r��:��d�DE��~~ �����Z�`5l�"9 gͼ���H�9)GD�)�@���]�9��<���׷���o���n��皺�[!�]�z6�R�vۑ�>m�����G��~���?~�37���(���n���=v�:�#���[:z�'	��&��&�� [I�@ݭN���t��� ��ڛ��NI$�EM�A�����h�K�[ngn.�s�*!����[A������u��SR�ڈeIr+1��vۓN�n��皺�ٱR�$�PrG}�k ��gb"#�'��{0��z�$݁�3i��GR����C�_�v�/|׿g/�XM�bXab��LIA Q�;?%�ߟ|�~����q�pt��E��m'=v�u�|ճ�f�� �d�F�Ȉ��4�����`W9Q��>��>^�� [I�@K`t��f�U��/	��1EkKlH��>���CYTq*ND��H@��y��mu.��`}���3[y�-���A*oՀ7�����n�8�p��ݻ<�W@ݤ�`5l�9�n���	��&��&�� [I�@ݤ�`5l����3��)�Hc�ʒ$�]�9��UʉJ��`�~:ko0"#�Ü��>q!BY^߶���w�]r�7vZ�w&�{X�[:�""&#���~���{��y�k�f�ۍ�ܒH	�\ic�)����GQ�a&3�i��ݞ3��v[�ڕ(�RqSq�t��݁�y��{�3]���Ӡ{Mǭ��R5U*8��m'=�9�L�S~�|��@�m� o�d�F�Ȉ��4�����`}�l�Ds�ko0����	�a����&��]s���ri�/ۻvy殅s���5�����@6�p��o0܎s�[��	S~�歝�����d$<����QC٠
�XXfPc�Z+ZHdHbB"d��h���>����u�~���  5�     t� p -6   6�            l      	         -�                                8� ���{`t�L�'9RV�%e8�0��u�UT:��mg��j����=��ѧ�m�Vsh0n��료�.8n: �umۃ���)�%aƲI�x�n��ډ�%�v�>����%t�v��pn;��}�83��\�A��O72tYul�[k�#�\�<G]�kl�l�#8ش�,�`�UST��������8�� ��� Ԏ8)@A��� ��[P����p-�� �f�f�j�힍he.g��p�+TU����؆R�T���#mZ$��ݶ���[��Q��O�������)MmNG���x�k�e3��&�cj,��`�	�u�N�"���t�x�)��o:vۂz�nt�u��7/Ⴭ�cu�:�ӭ�𓗞|V;s(\n����7NWOo\�Jer�e��;���{q\��k.Ѯ�+w]
��I.9�r<2��4�rgv�.�-.�l��p�q���Z�b�/�H��݌�62lv�`J���m�lq\j��;����
vW��rz6��zf� ��6;D�S���sm[g'Z*��z�ЭV�v���Ʈn��5U@���5�v����BV8]�VQ!j�j�N'�jt*�v�@@T�;\'Gi]�n�n��V�J���8�.怩$[d��$N�鹋b�Ci�$����fҜQi.��p��ܽ���lR	{���ޮ���GF�NE�P��v�5�k�b[%���8��(h#�E��zu���+nvwRi�\���'�m�kG=��˫6k{��ox
��>z|�$�HȀ��! 
���%�ݒ96��  �� ��     T�kizԽ[��]�:�(���t�y�n��n��m�{:���r��PvG]o`z@4ډSx�yy��g��yV����1cq�u�6��c�92��q6�%���I�IE읽�L�*l�tްa�m`	�-(g`�	���vgZ;Y�\���[���g�}u����ݙ2	���8+�R��3w%�j��u+l8��N��&u�Xi�(�B��M9J9���^j����`o�i�W �n����Ԥ6�j,���������t��`i}Y� ��M��}�]q2B��ܛy� �w�f�� {I�@ݤ�`Rf�ta�ѳ5�5��{�_�@!_�ן?���?:�������tcTꬨJF���G�`o�j����`o�i�/ۻv�ѯZM'$�I$��*�R �\��b�njW4x+y��ty_K���H������$��rR��RSN.��<�v�&�5���NzBN�l2��;UU��k|�U}��竂�$X��������#�T�X��!��I�0	�����F�i��w�n����Ս��{�Ma���@l�aMƛ�@�n����9n�N������. ���Ӕ��`o�j����`o�i�/ۻv�y�5)���Hӑty�:�"#��[:ko0�����	��e���Iù��k�`۵��:nn�j��L�N�n.�5Q��r��4���?�=V΁����'=�9�7i'X�ͦ�R�JN*r9�~�ۿ�?c�ˠf=����dӠ{Mǭ�Ҏ7#U*H��|�W@��f��W��W*RIA0b�$C�Z40�	�5]pԅ�����o���m�g�c�H��J:%IM8����R̶�X��5��r!�'=Bq���Q]��}K�u��t�wn��<��=���`~�l_�_�I��I$��GQ����������ɡ�<����Ӕ�v�&�t����(�7��?�˰�s�7kS�s��l��t\UDRi�Q˰7�5ty�5��t�wn��\�#�Ԥ1����9@J��`U��gͼ��s�5jw1��UG#w����+}�N�n��?�=�c ������rko��|J�ʥJN*r9�n��皺�����M:��*��Q��4�NI$�I*5����ba���4���u��tjR��]�]ۊ�{7}\��;[���B��s���]�N����3��`����b��GD�)�@��ٮ��Po�i�/�ݻ|�W@�񛱺��Q]Ci�.��`=V΁�&� {I�@�kS�$����l)��p�r���7n�����>��k�7�4���d�U�R�Sw��N��Z�`U��gɼ�4��D0B^�d�!J@Iӽ/ϻ��� �  �� m�     ڱ}tλ3a��=�m��@J�ls�{�ݺB"�s���^�	m�#=���A�E*�1g�*�#.D�97\a�n�c��zG)s
�u�lR�u�h7���R�98a;UӭF�̄�M(o�x�񚘲P\!k�v5t"�v;<��X�<��ٷ>(��f��F�%tv����h"R�1%(������J�+UTCۇ�xY�Y���:i�2��<��w7Nm��%�y�.5Y��sj��� �M�����3��~�D��o��7����7R�I�����V�� gɼ��u�>��� r���R�JN*r9�f�����}�%����7�4�g�6�I��O�9�?j�����U���Dr'��� ���8ێ�)GD�(n>���3fǪ��3u���u�5�n�f�Z�T���׭������Uu��k��5G��ȹ�Y�2&�P�F�[}Eu6�Wc���-�5���N���;�O���,m��%ʒ�6��{��!|�H���y�GJ������x�l�u:%�n"�ܧ�W�_@��3e��s��g�ߎ����`JL�n(��(��l����t֞`u:��f����T)��w���dӠȎz9ϗ���=)����;�?rw�?^�[��{S���-��b�n��<[�;�����c�䛒ێ'��������u�6~I� �[:K��F���	r�^�}�Uʢ��܎T�W������������]7R��RP�}�ٛ,�M:~���>���	7Hb�vCÁI9�9��f��u�7v7R�y�6�]�vX9�W���:���`u:�z9�T����w�E��7n���`r�\����<�����dӠfeb[$���m�$��J�ű���:��u��˘e�ܑ�{znJd�U�R��`j�k�^��`o�i�/ۻv�y��2J	wu�6u'y舉�#�'����{0>�}ٙ�58���
jE}��7�4����"" �u�6u'x��T�R�JN*r9�~�۰7�5t/{�^��HG.����o}�I��p�iI�n]��y���Ux�f�}�N�~�۰=����i9$�HQ]�늻s�=GO��ii�sd��y�z���ѱ$q�R��RSN.���͖�&�57�����]6?]�E�Of�{SW=��� �[;����Rk��ـ~����/fl�33{�����n4�:jo0:�t�Rw�=V΀�S�Q8���Sn]�\�+W�_@��͖�&����`n�JB$��R:���:���G#�9�y>��'�f�ٯ�{��I9$�$��nIRI$�   �    m�[V�j�M��p��/m�(5��i�3�m�&^�qv�,0*a��ClTj�Ӡ��tN���iٻ9Z��ܸ�@��V��&a4��&�e�������u���P�ݰ5۞�Tl] 
u��ƣg�f1a8��ګv��r�<��/pÍ��r��B3��i$Imٯ�T�{�"jA���<��)��z6��k[unzlvv�k�kǚ�f�%�MԨSR+��e��ɧ@�f������ٛ,Y�M@�J:��TԒN�����s�<��=)���o׀S�������J4���"�]��ٯ�|�'x �;������]U]AVM�pU]t9��ԝ���f�� kٯ�{0͑2[]Q.�i���e�}��@�M� �S����N��S.��YZ����#Y^�F��Mq�t���7+��"l�0.������޶]vț��}7S�N�]'���;�w�Gc�܎�;�J����w�L� �����N�kw�3u<� Sn�JB$��R6�}�y���͝��۰1{5��f����T)������ɉ�?_@�'���u�3�I��3i��GR���rI�/�ͻ�_@��f� �sg@�n��N7$�h���2t<����X��:ˆ�g�X�r{=�W�|��Nx�2P�ߛo��']>��`�;���`����(��%��/癮�>���/�ͻ�_x��6D�o�F��8�\���������|tT��-K{d��d
F���d��3��1��ɀL`ȡ"I�b�b�"���6���("�1��aPd�ٕ��3z0��o}Xk5���'��fay��:��[fP��PP�X:�sj��I���kE���j�h55M�0�H.��rK"%�2�̂�q����p�hΎ��=N3��X8ebRP!	�-C���J�8��C0R1��э�d I��a�h�����0� (�%O�`!`Q�U=E�J>�!� z � �IW��}�'��U�3k[�$��	��
��*�
������ �S���RN�5��o���D�6N"9M9v/f��<�v��΁~�m�fk�i4�����[&M�w�-��2�v�8.�ny�z�],y����1��1J�������n����O"0:�tZ�7Ԩ1H����ۛ;��Ifo�5f�}�y��Y�M@�J:��TӒ�f�y�)���>��`�;�f7�1ҍ'"U$NK�1{5���l������$! h9]�����ٱ��t:$(�%��/癮���6t��n�����3�Q�\n%$�IUyk�4�$nrp�OW%`�6�>�
l�d��!�9"d�֣]cO�u�ۛ:n���N�}I:�O�dQp����_��vr��_@��f� �sg@�Of�Q8���SN]��S���RN��L����$��jm�P"J)�#nG��UUTs��=���=�����`
u:��2*n$*��n`����k >i�@�9�'��~���z�ߵ�[Tؑ3C@R!H$�B)�R���u���y��~��@s�1��À �      ������+Bc���IN��c��o9=s�/\k��Y����+T���檭�eY25�V�s<1����;�&������V{6�<�hS^'��r��mgV�ݴm����X�u�g�fu�7u���`ls���;[�ۨ�1�hħY�\�`SVu<��^��kgf7g{����{��_�~*���VշdDs�icʝ��	�u�g�W]�טݞ3���M�*QԤ⦜�`�ݻ�_@��f�������tۺ���F��*�*��N�]>��`�;���`�v8ێ�D�������5�ۛ:�ٷ`b�k�g��%���(���_k >i�@��� S��@ϩ-vfoj'R���Crt��n�����/癮�>���/uj64�N@֒�X����;�Kv��I˭��}mF:��ͅP��N�q���l�J9Q9v/f�@ϩ'X�N��s����~�����$��R6�}�y��+�U����!I"(���~��o�}��������/=�1u*5JEY}�`��f�y�)��gԓ�W�hq�GQ:i�'@�{6�^�}�y��ۛ:�c{#(�r)�����N�]�m���y���ٷ`g����rI$�D���I�!W4F{���ĵx�w3zɞ������ag�D�������5�ܚt��o�W9�Y����7��Z�u�q>��`ճ�f�y�)��gԓ�noj'R���6��/�ͻ�_E�93�էX�l�u:.�U7W5y�)��gԓ�Z�t�N��SaNP"J)�#m��/癮�֭�7S�N�]܈�&�AꪦYZ��9�˷&Y��6�mU��3��ד2���Z���V��F�fq���v��_|��/;��3u<��u�3�I� �S��R��t�r��۰1{u���k�=�4����t�IȕI���n�}I:�5�g@��� ��q�萢T�9C�r�}������Uמ{�]W`~�ŒH$��
�@������U�~^��L���gX��v�殁~�m������5�݉%�m'$�I"D�.:�u��nwc��g��[&��K�G��Q�o6��ʅ'R�!�6�`}��������3�I��r9����z�~��QquqsW��n�}I:�5�s�3u<���#4z�t&�i&����`{)z99��`
}�W@ũ�]Q*R's�v�殁~�m������5���M@�J:%8�F���c�N�]>��`�9���9*��ET*J���vےI J��$�  � �`     �	�D(;JZ�4g��I��\�WB��8v�oWhBFX
����uQzJ6����R[dI.��m��wV��q�[s	Q�Ѱ��ۡ�\����H�U���;�!�����緭�9r�f^箫n��qg\��w�l��w+�S��K���p��:�ɹu�fm	���s[��Ͳ�^U���Rn�2M\�]զfn��pul�n)Z��QD�H��X�����5�ܚt��n�7����t:$(�%G�3�I��[:n���n��E�&K}q���q>��`{ri�/�ͻ=Ȉ�r���m7���ز	��
��UeM\�=�s�?$�� �{��3�I��y��o���D�'R�G*'.������$� �I�@��� �N&��UZ��P���i�3ln�[��˛������ә++i^z��U��c6��*��oϩ'X�Nzn���n�-L*�V]�U�^�d��~���$:	�DDE���y�})���$� s��LN*�Ҕ����f݁�ۯ�_�3]��ɧ@��odc���T�9.�S��@ϩ'X�l���`����t:$(�%G�/癮���Ӡ_��v/n����m&��I$�%P�vϭ�[[��ۆ�둛�r�X/�D�t�xz��ld�&K}q:�j�O�u�ܚt��� �[���V�X��A5RW*���:}�� �[���V�X�l��f�Q8	ԪQʉ˰1{u��^����x,xd��0�������X��bD�O9�p�9�DWo��t���56슸8⑶�����`{ri�/�ͻ�_@��h85I8b�;��5�g@��� S��@ϩ'X��[�� �=.p�v�G�Ů�ت�@��H;lV���,�ru���yf����� �[���RN�j��I�����r%RD��_W9\�H�i�V ���@ϵ<����T�AP\(�����_�ٮ���Ӡ_�ͻ�_@��3dL���u��8�\�=�l�����n�9�G+���XM��Bu(�n��m��������nM:fV%�Hۍ�ܒH�cda&���Sặn+X�Q�i�D�[-�狮Ux��Ԍ���N(�˰1{u���5�ܚt�ٷ`f�
r�8��U]t��:�5�g@ϵ<��u�/����I�����]��ɧ@��<�b&T����ju�9�캊�	�Jq�q�t�ٷ`b�����k�=�4���i�4
"8�Hܗ`b����ju�kV΁�jy�荍��ba�c��TE	�T�Ad��a�U�݀A,4�Lɬmۆ�$�E�k�a�$�|Z�Q��+:32fjvfZ�̓�maZ:gi#�P4��8 �wł dهIo3f�t���� (��n.��D�����`��R9��˦2�*-o�������� �     t� p -׮   m�            -�      H        �                                �  ���Y{�K�Z�V�g�V|;&Ҳ��;�����Z�r�<��Q�pv,�KR��s��^�h�:�;/��*y��wnÞ'����J����Ftۚ#vu^�W�t�W��T���`m�����������&;.�"Xh&ݏa�vյ��s�j68[��vJ�)M����n����h�� l�e(-�����[�À-�k�� 2 R�� [E�,Js�m ���S��ytA�^�#�۞x�y��kZAtB�7@@me�ȅ+d��7ul��@u�����Y����<�փ�t&��7�Qj�i:W�6uɹ��7d�ݜ���z�4�sEή� <�E����P�lb������,v�����%�4���sGnCN��Qۍ%��Rt�4m�\��p����٨{<�gW��:;{:wm�{:�$d��7�D�=-����mA���*s���RK����V�g��"�ۋ>���n����Ū�=��8��;�0k�nn;)I��P�ےku����Hh�LQ>��:sy��ڷJc��-��g�E��,`�-�HMU]V,�
���t��*��m!��CaV%r���^�iV6� b�U7 ��Z�p�Vp۶��1h6�l�=�o!l�0n\`3�:�-�c��#Hh�n�U�Tς�O�.ݹ4)��b���1Þ��]�짜sr�]%ظ�����{��t��u�����z����Vݧ@�YNwoG�]����jC��'vA�-��^�ڲ���xm�ո�����[������w���-�HV�C< �@�w2UT��[xp8  $ $ �      l�ݵg]�d�u�z�D�hʹ]s���9�;Gkfض��2,[r�K�b	$�+"�&�K��Mp�j�����4�:�u+��uj�%Gn�mq�+����+���m���\��њ���)c��q�Pd��-N�ێ	V�������q�u#��ѣt����[E�R��'A 8 8~�o���v��ok��1�Q��s�U��nz$��gs�3��6Ӻ�N�T��{]av\M]׀�Z�`ճ�g�<��u�{�l���\N�ڧ�v�#:|��N�]6�:��#O݋(N�C�pmà}���`b������`{ri�>�٬��2����Ix�n�mju�k��g�<�����!�N)n>�~~�v�殁fm������FƓI�$�H��=���n��!�K�Rx�qlp���{^5ƴn<�[9�j�p ґ���=�5t�3n�����/�ٮ����GMF�d�wu���}��X���T��emP�!,�a*B&b����#��S��@�Z�`�9�%N)��Q�RF��_@���]��y��_�ͻ �n�Q��@#%).�}Z�`�9�����n�ۦl���\N�ڧ�v�殁{6�^�}�~�v��ײ6�nI$��O�F��b7;=WkYn�s����6d�0n #�ԕ
�@�J��N.�{6�:�t��:�5�s��tXU�WS�9Dr�^�}�~�v�殁{6���JjRQ⑶����n��ϵ����?
_��B%#�I���V~���٣Q5I8iIU�����s��o��>����n����o�`~Y��4P����ܒ.�jy�)��gթ�������uS(ĵmI��­
�<�ǲ2KdD���lj���M�5��l�鎩k��:�t��:�5�s�>�� �$mGC	 �����_�ٮ�r�UT��O��>����n�ۢwsE�v�j;U1W5ھ������jy��92�{Ϡ}������(N�m*n8�7���m����{��}5�$��G7�\����/ٚ�S)ʜQ�#�`)��{���i��z���gڞ`/����A���5���f��� �iZ �\N����z�i���ح�q�ט����gթ������jy�)��oٛ�')�޻��W@��<��u�3��� s��u$up����]��m��������k�]s1�7������v/n���V�X�Nz�G"~��� y{�wT����FJRG�-{3e��y��_�����*�>�$�A��8�N6,aa`��=��}�  	 	 m      -�m�xH��[O��lm���p;&�-��NӖ�t�v��Fcr�w�� UE��H���Z�z���J�u�3�9�	YL�q���[n��Vc"�']-��\���#h�i�������U�������}"�eG[U��� 8����s�-ԞB�Ҹ���̲�`�
�����{ܝ�e����4�.М��F�'Q@����X��[�^���Z�j�=��٫���{��3Ry�6�d�N���j6J�i�6��/ٛv�n�N�� I[;�""&O5�QaW�*��7W�� o���:��%l��ͻ<<Қ���8�$����� I[:jO0����Nʲf%:����{�`fdӠ_�6��ݝ׳6Xۡ���q�$�DP�DCK�۱�4�T����է	�!u��c:x���4P�����$:�3n�>���-{3e���N������@�Q�RF�������1�z1���$bX�-�bNj"��1�&�������R`:h� Z(%f�F-ٲ�L��LV�3X%V��Cna�gb}��߾�X��N�~�۰�쑵�R.n��d�N�����3�oـ�ߧ@��3dL���u��8���32i�3Ry�6�d�N����E�7CMA��~�۰�vt^��`fdӠ^�j64�NI$�EIH)�vd�nwb��Ga���gYE��l�������1ʜQ�#�`n�������ɧ@�fm���Ԥ6�L��''@�ԝ�	+g@�I� |۾��I��*IԨ4�v���3&����gG �n�8a���P�R��o׍�W>����k����S�IL��!����Uq}����~��t^��`fdӠn���F%G#��� ��}'Rw�jV΁��������[��W{A��u�A��c�r�J:݆�اx3ٶ�7�J*�X�m[���]��I��[:jO=�s������7��\l�j�]NvX���&����w�2u*����@�1��p��ͻ �7g@��͖�&�s۬�9�9S�8G.�>M�@�ԝ��9�(����r"�V���iMJCh��H�rt^��`j��f�� >M�@I8�UUWUuTMΜ�i6�B['B��g��&h;Ie���7:h���Vl]d)�~���m�~�9��<��w�2u'xΧe�R(Q�T��r.�~�۰�vt^��`{j���i20*7H��`&�d�N��9��<���A8�A (��rt^��`f<��/ٛv��΁��f��-ƣK��f���%I�@�I� |۾���;�>��wݰrms�  �m      -�d��l�Ȝ��ș�ٷ;gS��Ѽxn�0�t=��W]��'�~�A���!�U[{j�A
����J��.3ȹJ�l�q�<E�Ӹ��c�x}����{7Ly]���wm7����v���1�ѯ8� ۛvژ��܁G��n(C��Hl������qY�z���zfݝ�\�r���u�=��{��P�5UT����_�}��8{#���%�Q{R�N�`p.�Ԓ�[�˭�vrY�{��f |۾���;���5���9�9S�9Dr��ݝ׳6X�5t�f݁�iMJCt�8�Ħ��N�� J������ ��}���pJ�u*R+}�e���W@�fm�ۻ:�fl�<���r�2ꮮ�f�� >m�@�ԝ�	Rs�I��=??~�u� 96NK��RT���(θ��2b��.��k�:��V��t�*7H��`n�������y��_�6�}�\��	FI#��Z�N�����Eت������ |۾���RG���d��.��]NvX�O@�I� |۾���;���XU���N.�~�۰�vt^��`f<��7=��C�C�8��G.�>�w�2u'xT��Ԟ`.;��������ԼIAZ���Ӷ���^����g4�;I�O*��\j�Np�s�5���u'xT��Ԟ`ͻ�䝕bT��Pb�[�{,ǚ��3n�>���-{3e���=�o�(4P��L��"�f���vt�W9��*|@U��e�0��1a��015�{ph���q�2 ,��f���ٌ:�1*��;��a#q#̀�ܰB�R�N�B�p%]����a8X�e�a�ŒFFl]�:6bkb�J���٢�E�3X�Ze�ĳ�"G0(����9�`�a��b��&6�-�k�� :E<^��]"�ڂ�B)� �1�O�~S�6+�C�VU�r��W9�'wr��=��7w�d`"TN:�I.�>���-{3e���W@�fm��^�'$IDI#��Zԝ�	Rs�3Ry�6�&�:������vϭv�=nG�3U�4���n�0{Y�268/1�m�1!󹏆��	Rs�3Ry�6�d�N��{P��:tƠӋ�_�6��ݝ׳6X�5t�n�QNU9O�9E�� |۾���;���f�� ^h�c�)�N$��׳6X�5t�f݂�r�/�vt�3`��$�E�M��w��*Nz���ɿ}��޾�kٛ,2���i9$�I$�I8E�נ
�Xe�ف�=�̒<�5���8(��h(4P��L��"��ͻ廯�Z�f�1殁����#�q�j]�����9�L�Jo׀7O��3Ry`�z��T ���>�kٛ,�9��<�>��t�Dꮬɫ�iu���s���<��/ٛv�7_@��͖�7���@�N��qt�c��M�@�ԝ��9��3S�U�H��   � �`     �U��$9��/���-��e4v�ݧ�kkBvK%ٸx�:��N0H�mi�*���b�U.bϬ<у�k��ٞ����q�<���\�n6խ��m�#��+t���0�ݱ4%�]!;3����.�!Ǣ+U�4��W9�p�s�h��l�t�&����#y�HSZ�#��������w��R���S�#�a�cO���ⵍ��e���x�\��7s>���u{�)�z�N�� �I�@�I偞h�c�)�N	���fl�5+g@�I����?�vU�13Qq)�����dӠ_�6��n��kٛ,���(4P����C�_�6��7]'Rw�jV΀�n�h���Ԓ��n��kٛ,fM:�3n���[I��I(��B(S�c�����,��D�Ile���k���e�e�bg�⤨�(�8�}׳6X̚tԞ~�r#���W@ԇꫫ2j��g�D�ʗ������Ȅ��	��	]��o��6Su�2u'x���	������ʪ��f�� �Su�2u'x�l���d���q�(�˰��/=����7��5+g@�I� ��ʛ���R�T����Z�f�ٓN�~�۰>Y���#cI��I$Hu!A#ś���mI�5uu�v�5�(��k���z��k6Iԅ1H�����&����`|�u��9h>Y��Xַ�(I��I!�3Ry���Dɲ���Jo׀jV��+�ʤ�߷���#��Ԓ�-���N���FD.G9<��]�V΁�7��׮�qRTH��Q���~�9�/�7��w�f����DD�?z��?��N(�[T��s���dӠ_�6��n��kٛ,Է(??�7�I$���y��駃�ٰ��mh�e6���Ge�p �I�	�
l�p�>���`})��:��G"9�n�t5�QpEJ��Q�囯���������{�t�f݁�h�c�)�N	��N�� J�������m�@$�pJ�u!LR+}�e���W@�fm�-�}�z���S�<͖��l(I��nE�/ٛv�w_@��͖c�]�n��N7$��R@�:j��c�Y���Im��&�Zډ����3Zi:0!�99�]�����-{3e���W@�fm�{v:��IQ�*�'@�ԝ�	Rs�3Ry�}-��}��ܕi�G�ۧS��c�]���`|�u�^��`o�{�$�&j4��@�I����d�N�=�s��Kv����ߙ(�*�t
9Dr����;���f�� qO���n��m���  � � l    UUQ)<p>'H=s��#]s۳�ͺ;i�s�L�Ou�V��x��,%�ClE����x6ȭ$�-�K��ii-�2t�f�(���Z���͏#f�7&:�鶌;�h�l��sGi�u(7;��kG	�X��q�,�04Y�g�H�΍Ч�;Gl�Xӵ���`�<��P�w�fg2� �l���n8{;�-͵DYɖ���i��xmv�d���u��������x�NzjO0�7]7S�����HS��{�`{j��ͻ囯�Z�f��k6
$�S�G"��<�>��t�I������n�T@!�99�]�����-{3e��y��_�6�}�F⤨�R�G��:��*NzjO0��]~ޟw��h *�;r��\Frp������]S�tGgb7Z;xi����?9f�{5}�*NzjO0��]'Rr��n��I�
L8�qt�f��A$��#����߾���s�����O}]s۬�S�N:�9v�w_@�ԝ�	Rs�3Ry�-)C��I���ȫ&j�d�N��9��<�>�����hpJ�u!LR+}�e���W@�I����d�N�[UUWUj�V�ݑEM��T����f�d��	�ua�@/]b�N�&�5��6��4}��Ԟ`KN�N��G�)̀�n�b ����I.��{��{%��y��_�6�}�Q�IQԨ�����}�}U�����(�BJ�(J!	-< =C{����]廯�}��\�U��Sn�]NvXi9��<�>��t?DDDr~�߯ ���w�I�
L8�p��ͻ幯�Z�f�=�N�{孭m&��I �i)�/DK3��R݂���G�!����%4g�3�wD�6�%�S��G(�]�����2u'x�l�?RO0�&tI5J2����Z�fˉ�t��۰>[���ٴ8%I:��)�����V΁���=��D�Ͻ��Jo׀}�f�F��'�jI�~�۰>[��WY�����`��*����ʺ���Ѫ�:���Ԓ��kٛ,̚t�f݁�wZM'$�I$�s�Ug�)�1��b����Q�l7[m��Ms��=��9Q�IQ�*�'@��͖�&����`|�u���l�J��F��t��s���dӠ_�6��n��kٛ,�oj���0q6��/ٛxқ����;�5+g@k[������Q�囯�Z�f�ٓN��UU/�w�����Ҁ��J�&'%t�I��V΁����I�@��C��#�̼!�$kB�n(�6D�NCj��M6�tj�6Z�Q��!� � �V	5(bB�bD!�d&4�@N���,f"mN$�� 7Z`�ձu��F4���a8 Q�Bp�'K��9��+#I�1`�a1&*Ia��M�31
��iL�M�H��0�&B(* ��m���`F3�1�f%��Ngn�u��6�堃J�F��0���9�� 6:M�A�C���������&���6�f�3$UU�˻q;��ο��  [@     -�� ?x|I�l   �`            6�               �                       |�       � �=:[/q�תܦ�q���m��R�.x��ݎКj���׉��bt�%Z��*�R��d�m\l��sx��ts\vPv��7m3�6tǂ�7�v��Y
��i�y��	C	�mǃ�g���+�MѶ�lSl���'^`�nC��b�b�cWO����U�)�X�V^��f�y��hk��H�h 6�mp �:AJ���oR� � �p� �-�HYF� 2z�-��  ����ԚM7��Κ[���=�T��,qժ�v(�eT�(qe�%�#�q����W���s��h��E7k����]��q����r�r�u��X�#lqz6Ƙ�"]nyb�@�x�θ�Y(�㮹宓c�PE�lwnǳ��c��p�vk�cO6�G_�ۭvݧ�k���V���n7�ݽ^�k��p�a����ݭx�6����v�ݱt��0�w,Uv����Au)R�\|O��4�[X��B(u/(����l�7% Pr ޶0�׶��ݗ�,�cc1�V�� �sLd֬�������Q(8�|�s�yH�7e{<�5S���q�@V[�Ö�W��ۥZ������Т���x��ە2Khe�V(2@�a̳�+5UUUR�5U^ѡ��q������T�����m�:ډ��c��bAUC獺�[yRs�U:�8�%�������R�E��k.6ŷ9�Mk'f��́���۹��Vn�g��Rs���pF�z�	k�x���Ƶ6#.��%�x��srv��(Su�:�0l6D���V1�|�v>���ci���<��<Xد�G�� ��� ��;C�W��^[�{����1� � �     UUm��t-���:���j���֋f��Ė�E�^]���V�E� �Rn�$� �k��Gka����[��ʖ����#���{Y7����ͬ��c�����x�nӸ�b�e5��w��N]Z��[���1��h]�9ں�蝬�d
�d�۶1�Y�t��ldkt�{\^���;����{��������\���� U��N�\�	l�	��hho[�tC<��[�i��M��F��`�y������a�5'�ғ����;����n��
q�$:�3n��fk������2i�7sv5Q �Q8��^���d�N���tԞ`���9)*!�Q�#������2i�/ٛv�3_@��f�$�O�o��9=����V΁����I�@�ԝ�����ʂUU F3��^���'d~����Vo\��q8�n�	-��zۄ(*檬�>M�0�'] �I��#�_ ���t۟�2QNU8�r���JN�����V΁����Dr&F����*����f���fM:�3n��fk��f��T�d��U����[:jO0�'] �I� ř�Q��	H�RHt�f݁�����f���2i�/(�֓I�$� �[6���H�ۖ�R������ �q��\$��Q���C�*�JIv�3k��>�%l��<���Quw	QJUR>�_�7�ٓN�~�۰>Y�����=���I*���i�u��s������W^{��uz��&i�e�� XU�Mı "c* �D4�y�}޹U�~������B�u(6�:�3n��Zu�ԟp�����"�"��&�ຼ�>��ts�����~�~:�3n���ײ6�q�$�Ru8rB�ˍI,��\��L�v/'_<�W7Nm�q�W��v˱)JT)19@/ٛ�=�N�~�۰>[���٠��$��1Im��� �[:jO0��] �I� R��Gt% S�9!�/ٛv�s_@/ٛ�=�N������C��"����i�@3R}��g@��9�"�$BWn{�km��}n.��;��������jO��l��<�>�������i9$�INAҜ!+g�z���b� �s�ۜ�x��k��ם	UU߃�'���Nw�{&����`|�5�����5fk�$�8�0q���/ٛ��Ӯ�f���-V΀ַE�qN0��9v�s_@/ٛ�?r������@�7]��3D��AJR�I������ �[:jO0��]7S��*IӔ�R[}�{`g�i�/ٛv�s_@/ٛ� �c�ܒITN  @ ��       r��h͔[��;kXw7c��xa6��b�-��q+ �C�Tq������j���G3�ivvz�)㧡�w1ŭ�,8��Gpw>�{<Q)v=�'����zX�X*�Nz�Q�8M��ݮ�t� a���l�ѕ�\�gW%»q�v���%�"��W�n^�M��n ��<�^�+=������/���G���<T6	�LmД�N8䅁�n��幯�Z�'��N�tG��wu���Ye���`KN�N�� Z��5'��݃��)""J*8�}׳6X�t�f݁����>�ٲI*���sE\�j�x�l��<�>��t=���7K����I:�I�n���܎my���7���g@�(S?Clٶ	��n��IeT�V��V��[��;X7d�Vʡ�M�N�sw3�m7��Ӯ���;��g@�I� ���)NA19@��͗��*s*�<�r">�w��t�y�}-:���C�T��)��V����2i�/ٛ�{���ϟ��})�^ �'d�]U�8��3n��nk��3e��ɧ@��ݒ:&�S�8�幵�=ȏ������z$�`��M������7RȲ���x9�#b��օ�3X�qٻF�2�ӱVzmph��������w�-��bI����}�f�$�O����8���3�5t�ͻ廯�Z�͗�#����I>N&5C��@�w]�����*���UQ�
���$�D��		iP$�JF� �$J��W�<͖h�W@���%�T����N]�����-ff�<�W@��۰7�h.�R��Rbn>�k36�G9ݿN�oـ}-���9�|�����A���I�g����ѵ&������;y5�v�F"�Ǫ�b�6�����{ �?O@ē��m�@�I;�1{6IM��"�q�@��۰>[��JI� ��t�wu�5VW7WWy�}-��)'xJ��1$��3۰u%$DIEG�����wL�~:$�`8�rv���|�������i�.�;,̚t�ͻ廯�Z�͖��^��JI$�I"#��mvZ{nvl�:�԰�r�
�O"��7�@�|�Lj�n�3n��n���3e���N����J)ʩ!I�����d���	+g@ē���D�Sbn>�k36X�4���v�w_@��h5Bl��rNW{��V΁�'�қ����w�y{6IM��"�q��Qy��`})��)'x�l��Q�ȎD?W�mߠ-�8    m�     �n��e�v�텫N�ڷ/g��s����<=p���h�!bەX)햢5kb�J��,hZ����W�n��=��a�캧=�ë�#�;zl��k�=z�e�����l��b��s� 6C�
�&��*TjM<B�^����v{ˤ+���\<Q����ۿ�}�����e���86��j��c�S��ԅ��p��s���i�q�����]Oc�Մ]����@9_�W@�I;�5+g@��۰��%$4IEG��Zĝ����bI�����ɺߪ��%�ӫ�&��s��������v�7_@���,^�j&'S�P�màbI����d������5��(�*�h�$"r��n��k36X̚t�f݁��s]�ƓI�$�H�7�/=]W��,WY+�7҇�-�Xo.h�ŝ�k��p�%B�q�,�}��à_����1���i��d�S�[�{xJ���IȂLԞ`:�t^��`b�l"��E8��ɿf��z�N�� I[:i����P��T�%$���9������>Y��X�4��ͻ �n�pP����T����:��%l��<�>��t'���t���u� +i�m��]����=5ɫG�SoZ��$v�kosH�W_��o��.�5}�%l��y�}-��)f�W�Z����T8�p���v�ۮ���w�$���n��*�.�)I��廯�Z�͖}|�UX��L�L$��&!R���$I"&�kXY���h��=�%1�I�$$��Z�cF��Af�2X�-Jl��e�d�XD�aD��"�c�� �"R����58��N����Fo�c3[�Nh#Z&N�:H"Ȭf,��Γ]��[A���b��Db������#��N���S��	aeٻF���jMZ߽]�:tq�G'�4��c2du`�)8bsC��T5��`�fS"���qa��#4l��T$�	Ң��*v�'�	�T ��Q���������O IE�Ul������4\(�6MU�@�ԝ�	+g@�I����_��J@�%2���{�`fdӠ_�6��kٛ,����q�ے�DnAQEM��T����f�d���9��
-���J���#��JlQ�Ht�f����d�N����6����&䢤Q)%�-�}׳6X�4��ͻ �n�pP����r8�}֤� I[:jO0��]�:���o�:�X�S��fM:�3n��_�g+b�D ~����(J�8��߽,�kQ18��6�:jO0�7='Rw�$��܎s��~��O�A���
�&���f�v,Tl7$g�M��*���;�wJ�λswR7vW��o�ޞ�g�V��	+g�""�}���������"C�����M� ��t�<�>t���L*n�&�L�"���`fdӠg�6��ksvX�����E��jO0�7=%�� I[:Z��
�䢜Q�%�k�]���32i�3ٛv�+�\��D'�I"J�� @@ [@    *��	3cK;%���+ɂ룓��.+>�]�l��b
�:���l$�c3�� UE��H�.�Rg���D�Ji��s�6H�[�����`�M&`�z�[v�ݸt�2]t�r���m���� m��i�"�[<l����T\��|�sGOsG.,i3h�w3Xz�1ծ08N��v)���)�3��H���1\g���w덦�pny��M���3�s%G[5��h��I?�������f�� ��s�>�S����}��������32i�/ٛv��W@��͖�f��JP�màf�� ��s�2u'xJ����S�R4R�r��kٛ,̚t�f݁�3Au�b���cn.���w�$��O0�7=$��UYej��絣g
�f�'Bi�iL����\���[pi��Ϋd��]s����{xJ��1$� ��s�#��H}/w��5f��RS`��drI�y���/f���o.���g*�{ٲ��ɧ@���R:	�E8�R^`:nzJI� ��tI<���E	B��(�����3e���N�y��`}�5t��krJ��ӭ���]��� �[:$�`:nzJI������0�UU@�������q8{#���%�9��ڳ�ҀY��΄��Hp�r�T8�p�>���`}�utY����ɧ@���%��)I9v���@�ԝ�U��f�� z&ڰb���cr.�kٛ,�M:&�Qȉf�"HI;U��Ϲ����ˠ_��J@�%2���{�`-V΁����I�C�ȉ��~���ЊJlQ�I!�/ٛv��W@��͖{&�ﲌ��i9$�I#�{kf�ue��%�)ֹ͇i�I�l�Ƹ�i�1�Q�(�
�䢜Q�%�k�]%$� Z��O0kqus77�M����ws�2RN�܈���~:Ϳe�����>�ٲI)۝:�SM���e��[:$�`:NzJI� �'S�JP�mà^fm�k�]��}�}W��& �*zE;�{?���̔B*�l�$��k͞���w�-V΁�'��Nf��v�Y�ZܒΏ5��:��Z{�l���sv�zڸW���.	����-m�%$� Z��O0�'=7S
���)��W���=�N�y��`}�5t^��`b��E%6
(�G$���<�>t���I� �[:i�D�T'%�I.��9Uʥ��.����x�l��<�������77E��@�ԝ�U��f���"/�����$�������H�\�  ��m      -��z��O��������ֹw^dϳy�`���P۫���ad� �ȇ5Um�UR�ڱY��*�X��E$ֶ^��\c���1�.�����%4�n�M�ێ@������m���Ƙ��6:��X�ms���a��j �V�;8�cp:�=���-��+Z�myr�eu�������}��;~( �UPs���6Ls�t��p��S3Y1q�q���]<v��H
��<s�[�ru9ـ}������`}�5t^��`j�֢br�A�m�:jO0�'='Rw�-V΀��Q����#�`}�5t^��`g�i�/ٛv���QFNA���z�""'�M������<�>t�t��hr��mJe9�����dӠf�� ��s�2u'x������ ����efm%��Mg.���@S��dE8�힨8ti�˱�5V�m��$� ��s�2u'x�l����	��I.��<��W9�q#��6X�t�f݀g�j8�R�ME)T����:���tԞ`i��}��$��΋��m���e��r�������&���nzN�� S����.P(5C���~�۰?s��o�`|�w��7�4�fV%�Hۍ�$�I �{sY^�B{U����:7��3�T��I�FU�n+���B*�l��Dr���]׳6X�t�f݁�3D��TQ��m����bM� z�����'==���$�R��.>����dӠ}�߷_�$y�C �3�7ko����f�G`��drI���v��'= �M� I[:z��w$�4�q�R]�����{7{`fdӠ}�ݻ3t:�M'$�I(�.����x�=��z�����7
۠D�-;��
��R��"�����32i�>��݁����/�͒IN���M�;����	+g@�[y�|�9��o���=u�	�P�Mà}�ݻ�y���n���dӠnf� EB6Rr"�� ��s���p��м��1ȱ���Ch�Z[�)mT&��fִV8E���4A4A�0j&%��	�	o�[l]�Qa��h ca�ivh�;�{��3D��TQ�Tqt�M� [I�@�[y�|���Ӣ���p{e^L-���yd5��]�he����yw�䫃�U��vn�*\�W��}���9�ko0�7= �M� R��G`�##�Ⱥ��ۿ�U�H�����O�� �'=�s��=��\rLUYs3w������o�T����݀{۱��R�ME)Td�t����	Rs�>��`{���zz�?]��W�n�*�o���{�%I�@�r"9�^��[~�'����}��������?B@ ��  �/�E�������p�� ����iP$E^�D2�T ���5��T�$$�o����~?���ߏ����_�������݇����������?'��o�����?��H  �O��������$ � ����D����O�����C�����~��  �A����~��s��iY��������?��?��?����x
"���
䨓*$$���
L��*$�(�*�B�$�$�)�L���HJ�H)	!!!+,�	,HB�� @�
��"��*���@�!(�*� �@��!���#H��H
���B� J�! $!"$��2�H��*@B���B$�0��) H�(H	��$���0�
������B*@B H� J� B!
��$2#@ B�!*0��!*� B�!((@� 2�"���,� �H(�(�!*! H�B*H�B�! ��B) H� ��(H,� ��� @��" B��²�H��2)B�(@ J2� B��� H,,	B�!H� Ȳ�H`��#JB0�!"� �0� B(��#���2!�$�"��� ��2�����J1̃�0���* ��l���������A@ #������~����i������"� ��Y��������3�a?7�$ ��l�'�����hE  ��� �O�G�w�@ ?/�;�X�� O�E����Y�r��,���z6l@ /�������E  �O�}T�_��w�������P!  '�  �'���6a��)T����_���?��Q�ˠ�� :;/�I����:�����~?�"� b�~U�H ���޿ӿ��߷��������
�2�̆��@�&�����9�>��|4��T� RDT�@ *D" ���)E�
�% *���  T@�R���EJ	E	*��  @(   ��E%��(
��)A  T`    ��     f���Uf�j˛:�ŝz��>� ov���˷�����qO�(>��>��4����  ;���qڥ� �Ub�6��z�{��Ub������.��2}W�r��3ݵx  |�@ �
�(  dE�|�Ҕ���i��� � (� A@��DJ �
��0 ��   �� @�� �% Q �  �@  P" �:Q�@D�  �P  �P � @���D�������s5�ox (��Vgv�Ǳ�ny�z�F{n �J�w�+�}�O� ۟-*w;v�/@4w�L��=��eUeܷ���W� }y\vr���{�s;m�ݶ� o���  �
  	.� �ӗ|,��M{�g�w��=|}� 9��s;����]�{���Ӑ` oAfx�ru� .,�mɮ[� �Qc�I�[��99t���fz�qg}��m:��zz�  ��*  �   c`��A�����xům8 Ԗm�w��{���gk94;��Ξ�v�ww� ���������o� +w��퇼ڻ�Sɕ������ ����J��}���s�����    OPSm*R��`  ��Bf�T� ��Ǫ�B���&��T��*)�  T��%6�JU@ Ԕ� 	�._�����G�������,�MC�m��
Q
�w��DWJ���U��"��Ȉ
� ES��ѲA, ��B��2!C ��W����Mk{�g�u��x#����:�_oa��x��橬��^f'�%�Vf��3�|0��7^��7�n��M�[)��� �d1���P�^���q��~���e0tq�\c���l�{��3��k��u�����o)��q������/������!5W�{U��;^}ի�a��'��7����m�kf���e#s~]�!hKk���S̞���ak�asM��h��6�G4�-`�LM� ��x��$�����Ћ�, ��	��=a�>պ�M�*`�xs���p��)Sf�i�F�z޲����F����%>�/���2ҥ�Lߴ�0�^|$*J�ixץ�5T�]�ث7SO�#�j���V��ߐ����]�}��	���{U՛]�ԫ��MUZ��S^������N���k����.HN�{����73o�g��ë���o�}� \��6��̽�G����[��L�[i��HGY��NJ��5���LR2C|�M:��Tt0�"DF1������ Pr
EB��$�04�$4�ӦB��xW�e�F�v&� 5���y�!8�!�i h�C��Xa���y������z_#2�M��j#+��d��J��L��6Bp��0�K�s�ͅ<8�CI����d$a<�5�$��&��f��$Q�-Y,���"H���R��0l���yvaN1���A�	�ǕZԒT���k�ݵ�ʫ��9�x3F�浯>&�%��t�.j�������|�,�uo<�7ֹ��m��hÚ8��[�&3[0�L0�x�Ml���t�<���_�g���Zu��֏y$!Ѧ�����Wb��kنa�ōk���7ɘM֦�%B0���Yr����4���R��h H#B"�H�1�� j�H\5���F؄Ypu��&�|�h������@��y�c�NBB�i����w0�ǁ���T�Xh�<�������6Sֺ%�CIP�Z�~��XA�4�8W�!L���<~��c���2�h�q6���M�<|B5���H��[}&��OM��#\4kzפ�==v�������g5����u��s�|��O�Ħ)�����x�p�ձwzU�^Ym?�ϩ�Ye��p��=�k������55�S=���8fM<
�<Q�3T�g<�缵�u+H����u��o���]�;�4��	�yr~U�����j����+:��[�_5��P��i�ĦM���ݻ�S�� qR4a��hb�n��l�̜�5�^;<J��=4��=p8S�R�`��˥�j���d�Lj�������f��.�	�W����A�n�r+H��+�e�����OW��e�n�b��`B�0��8a�0��$�4l8�O�^;��+{T�߳�����m��=~����ˬ���^"���@##Z�yu���׸s�g����]��m�ҽ��K�'�|��y��-��W���y���+�`�WԢ�����=�E� �	�C5��^��L��1�i�xx{�Jm�
����P$9y&z�+��3�GF���s[���xy ��6q��޼�|��99��[�F����ס
`ku��+D0C
&&�"Q0tl�5�j\I�w\|H�A���xa.a�lk�F�>��&����u�,}cHjݛN4׏����9�=�/# �l���߇����|(��Fp������S&�7�pfsI"���y_���#�$��{�u����&��I�K�޽��!��׬��0=w�Ho��^�.�9���:n$1�1�_a��}qXU�6�_�8�O��S���<5�YW�y|�)�at�}�-3@n SI����R0
�l�����6�x��<rG����<}y0����)�D�RA WB�**�����U���-Bv���K������~��}^��9rE���oܼ��>���N�>��7���~U���T^1�޽�v����b�S~��ˍV���˼�۷�^���C�4&�<�r��Y�T��D�^�Z�K�*T��iR�E�V{k���+��2���-V�����~�\4n�===�B�,����g�����G�&U�S��~�^��hh��#�b߳���-qӶQ 05
g0�8^雼����h���3W��to|�U�W���������τ�w��x]��/O�!�U��#s��O췕�X-����+yz�ZW�W�=f��ƾ�������GZ6)$hkg�
���s�<<���H�CBĩ�D�&T B(�H�a]�4�<�d�#L��{o:�ɷ�ᧆkų�R��m�~�c[�T���.���;Α�CE	���*|��v_|*��}�#ȍ��# ������?&����<4h�����`h�a�<8o)븒g��8S^�ȁ�=B����Қ���)�F���ȕqJ�)�9O=��|��A
���S&fFCF���9�r<16�H\4�dOxzi4����P�a9�X!����6�H��W��Z��?���ʖ�/,cć��=�W�w7�P�٤�h��di��q��<w�<׼���;9b�K��y�<��<<�3[�|�_,5�׌.��jf�y5Z���{��-~����^�_޷F5��u-Ht����0i�S�[�b򦂼����5����n�
����u���2�l�!at���Ѯm����k�EH��ϯ�^�݂�}k1��~��Z�F�k�5�D��Ѕ$&Ny���"�O��3p�nÜ�Na���ϰ�h�F��J�0#B���t*�3�p�F9V4�a�P�8x
f��8xp�B���a��J��^!
a� �\`b���	��
ᆶr������d���^����.�'��44�#DҹZ���P�Y���]��>��a��R���G�A��$n�3���� S5��Þ<v�!�����^ڿ	g�[B~I�i��^W��)��"Ab�H=�׬JX."��aM&�!�(:X,`� 1,0�)�N|�_s��u{#�!Z��զٺ����r��q=+�.���k�`B��5���x��n��w��̗����1aq��Ŧ:���4��/7u�>6�$5k/^�w^��*�ϑ�t��6g��{�j��MNfϴ���/R���>�Q�$��X���W��k8��	�T��y����'�$.�l�9���_�LFS�ɞ�p�D�
�h����B!
f�L��6���ٲsk�	)���rTә�h=��!}�aW�\��<�>T+�3R����4�D��)$i � +A�H)�Ɗ�E���FA"�Coʑ����Ug/��N��}�V}X���q�M���f.��BzI�
�����j��;Fw*y��_*�I���"TZ������ք��=Yv��Ys��k��ᣁ#FK�6o=�<�x1�h�8o�rs6��-��%�ҋ-1�5����l5�&�f�w�5�+ˬ�q��E��tC��D��@*0�%��CA
M,\Tņ�����77|�˞�{
2�{�o�^��B�2��|g��M��}k1���'J�/fay�����ĩҿ�ν/U��ku���Eny�{{����z�7���s6K���k<� U��8@I
e�Q|��*Bu�N�>)�4�ɭ���, ��Xj��9sZ|��܇��WG���R�9Q�v�)A�Ժ��h2oA�0��S��|�E�M�Ԅ�0a�CR+J��0���\���[�K��XXI]1�����ĉ7������%'��XCF��K)�#���i�P�5��L5�M_0���6q��q=p|c�y�ɌOH��'1�8i�֜Bh�����y��<|#�=�4{��Es���~���~6��fj���0׋ ]��Z��=��h��}�Kf��6�{㼯�k4�^i*R���8B�75f�M2��=��2k<O6��<��cļ�c�_���j�ev�%��	]��l��j�S{8c����/��!�ʄ(۷3'<�+]&�;0Ѣ֐�RR�" 4��DnHiWi)"�b/���焆����~o���lє��~zW?=�{��7�     �     ���     m�          .t���zQ���[Kl���6h�v��]$��h���M]	�J5l�I|�d�4��۶̱��D:�l��$�Qm+EMˋh8�m#�M�y�>��;`O��U�C�봏E���@���3�{<�n�m�&��e`    m�  �| �      ���|       �                                       ��   m                                ��   �          �>  S%R����gRlq��ط[��˦�m�UJ��Z�iY�VX)�Z��`j��*�[iV�U�\a�j�3�%�m�rβ 	z[oXn�d�8   H "Z����h�����Ͱ m   [@m�!#qh�� 6�l�4�`L�-:��
�Uj@�b�m�m�����`4Pl  8���l���ٽ��f��d���l [@  �`�l	 �P���[@ 9 ,]��
%�����ʲ��a��Huٶ �$ 6�  �<D�$U��b�]UI���     ����	; ���h�ڐ ��8[m�e��K�K;jm��%Zꢍ�6������M��鶷.9�6 �m䩕�  l[��Ck�Ͷ��k�@6�e<�U)(���cWlL�,ʵ�骶kgB�U�f�$�!v��8 �K�.j�]�jn��筪��<�v ��1�lA�s��<��U���'"w�qN���q�ӷd㭢F.�ݗ��mmlԫK���L�V릐6NTdj�U��QqF�c!hw '0i� ���� Gn˦���$k}B����	 -�h�k5�v�GO��>+TF�JJ�++TpA[i3�Gi.i��nFKbIq��Ɍ�l�: �2H�mR� .I)�xh��g�`eh7�� �l(��H�6��Rʲ�-�j^UY8��m��8uK�R
�Um�����(5R(-����  ��^tm]P-�h��9ivA�t�Ѻ�,R��@P6]����UUA�Uςt�U��"�
�:=����(���_��/�k�*��UtӲ�b9&8�"�Y�6���I[���F�l,3j[u4�	ioi�Ӏ��)[kW�a�ĝvt�p[i�;D�c��κh�������:R�%�m��E��%U[Oe���y��lqA�V|��r�܄�	�Ѫt�Kumn�����i ] 󲨨�b���~|��:��j�-�X[l�2��,�*�$KU��I[�qN���8m�ٽ+m�ӧi�I`�ښ�*T$99�t-V��&7@tX�UTc+d�vM��kj�%}�h{����A<j�U�Ӡ'�����۶��"C���U����D�ͧY��H.�g5� UU�-��j�+U�'�ӱ�Ȇ{�v�[d6^�Hh��Z�a܅��j��eS$ :t )e���m�l�J��������#s�!�;x'�eZ�j�X
u���<�Õ#�ӻ��[�LqTs�ݗ.������[h퀞^W\�s�q�	�Z�-n���q��Vx�Fl�b������]A[��α��<���Ө4k�ɵTQ�ju���tK�s��M�V�q��f�Xҥ�=�(�nwX^-���*��=�O+A&���W!���ɲ�[`2�֎6{[�{p��l=��n����L�W�_2�pVS<]UU��m�g��:z��Z@VۥeK�:9]4��%�Y��b�æ4+]]�V��C�1�xU��8'/B����+j�����y�V�ZUf�g��vM�V��.�^�m{M��η6 kZ	e�Ŗ�8�6m���m�@��xm  �m�  ��� 	 �#L���  �� K(p�m��m����\n���d��kv�hh  p���j  	�h ��ݴ��-������5�vv8pkXkM����`�az�u[��  8mq��ml�����r]�1�6� �}��m�� H� p 6�  	  �L�m�     �Ɯ���5V� � ���*����Pe���u�7j��a��8h�m�M����   :d�m�8�&�6�[@��� �� m&�촛]"ޠ�u�n�k� �u��@ ��J    m-��e*�ܲ�Լ�UR�T��   H�3�m m k�    �� t�ݷkh6�#��Wp ���V�I��p�`F�ۀ� ��\��v�   m��m m�x^m4���|���v��6�          a%�pq��mW�V��  -��  �m�h6� Hp�I%��[m� �-��6�A�|8Z��i    m � [@&�p�!ڧl�     kX� �-�6�  v�g]ׅ�Ւ9si�n 0,s�-��l$6ͦ�L h 	 8:v���`��v�۶�� '8r� m��Y:��[�l� 8 X`k����:kn;m�� ���m�M@8 H۔�m�` ���z�{5�k�m� ��/5�ʹ�fiݶ  ۖ�D	��UU.�&3b�N���[z}׾�I@nհ�c��D���p�`
�*�ƌ� �2�*�J�.�U[�6��	����(�LgIS`�r�4��/�����@m����:�:�
꠮Q�n�0�[�PM�q <�f�v�cNԲh��Ύ�8p�m�I��%� ,�ݶq%����շ�N����3��ƻIR�9M�˻-���,���d ��'PqէM@l��V-κS�²6�ت��q5��Q�qm/�v.��k$n9ct��W�U�Z���mAV.Nz7�����x.�Z�A���W�O�������Y4������Q��z1gKP�hZ��н�$�|�>{�|3M�l��^6�Jݴ	���Hkq*q����ڪ�Wm�g���rE�u$�gky;N��D����aV�eV��dمv~��S��2B��4 �M$Ӕ���	2 -�o^�ȸm�-�m���z��+�E����׏o�D�|�e8i�$萑��-�V��  ⎽��� �ղ��6�m�^Z�n��J�Ҭ�� ���RNY:�$ $ m���hI�R^ZRV�u �rp�W���m��I&�m��smj�ˋ�� U�� [@ l� ��J�u�Gʡ�Öl�n��p 9&�l�o4Ѷݶ��p$��8��l9��� $Xa;k�@�_v���M�M���H�`�I:Z�sm�l RN�IJ��*��(�ÛD����:{ne+�Κ�h[n���Lv	 q��7kk)�y]�ű�������n�j��a�Ҁ����@f�����.�,�=�l#��]�a��l�utUu���u�ۊZ;Oe᮪�˃��6
�����uG�$$9$�,� $&�&�Ų�]��mJ��7e�6*���V�ڕ���Vҽ;;K���j��U������@vZ�
U�z۪ ���]�m��p-� zm�^Uj�Em�^���Y�h�we��k����2IG  [@9���  �]m[�w$V��m�
�ݶ���'
�2��T�v���l�R�uD�(��UR��zg�&�z���Z� �� �CA�,��I�:N�JIի�~>�{�66m�[\�L�q�*�/ �UvK����b�*�8r�v�i�ѵ�����k��G��e9Q'd��� .��'A���P*��0q�k��J�m�z�u��ʒ�r�n�� 5�  -M�Z�W��|��nW`�a5aU�����;b�r�[����l$��-���N��U�5m,�;!᪯[Sn�+r��S�+�Ή���b���93��UT��1Q�Z;`v&P�vA����k��M�0��H:��4��&�9m  �����������-�-6�	�V�   8[@  -� pu�Y ���md�l�[@     �g     X`M�2��8$zB [[-�` �` ��  h�>m���K�m��h2�Ā  6Z4Pl�sm�/Z�rlm 	�e���		 -��<t����N�]�WI��ԽU�V�y�h�ۯ'C����sm��ͣ�jU��v�L�ln�p�ڃpҭJ[ʚ�p��7�'�`�n�m���m�̇lv�A��WV^켄�ogw�'�ڠt��t��rީ���&�n�(m�Y%p/�_�Ŵ�ւt��6�y���T�r����gN��Pƌ��^7_�mn�,r�\��I&�5e��f����TT�J�#�*��@� ~P�J�@@4���_�)�Q߀=P8�� $G`!�W`���T��"��� *iE�	�H;\�F!#@X�1�B�!#`�"EH�
������!1c�E#Db�B �`�"c�1���"��H�d! �$�H2H�b1`@H+!$d"B0�1�HFB��bAH�F*�1#�Q��1��`��,X�B�`�@B�H(�B,�,R`E!��1$$�#	H�O�PT�pV>���X�V)6��O�G��
x(�	�D�1`A��E�$ B��da$# ��A�2E�P��V�B���A���(i�
 |lH(��OTИ (� �q �$B '��8)�)�P�C�Q�؂��@q 1dT�@� �LD�@����!�@Aډ��� ��(��(�8 h�*�+�Q���#�"�b(|@#A1$�� ���)��U���4��@
��Fx��ȃ�A��*�Q����.	j
����@CJ<@��H?(��A
D�CH������(PD<H��D@U~Q� ���Eb ����kE��m� ���u��۱��,��C���v��
�!�;MճE �h5�		 h-�    m� �  ���� ��F�uU�izt�MD4��^�����6 4��k��om��G����,��n���ޫ�����W<
�@�Ԥ�+�nS�5oUG�Ҭ��^�L�M�b��z�Ny|��n��O0��nчVkV��n:��u���;Hh�{q�����$s�pv	[��n����c��<��֝�`�c�F#n�]���
����q6m��v�F����m0�ۮ�;q�����s��A�X��7E��x3���SZ�"[6����NU�]��ݽ����;[7k���m��x� ��j������zG��(���z5v{ �<盝�nE�"k+Gm9�1�۷U�݆��5x���8�.��z��28���*��S�l╕iZ��m��`Tr�q��Q,�<ѕ�gӡs �j[�U.x�
�n��檨���5-�m�q1�$�½�*�WO��fPxW�mR��I���P��⪮UH�BiגIm���k6�����Q�T6G4�.Y���C�rɸH��q�����3���$j���6�yܪϮΠwd:,ܦ��_E�p�{g7�v���0�E��f�n�4�칷������M���7Xɂ�ѶV��'��p�֘5\�h*���y����q�{.U����窤�[	��	���Ev�8�õ���c�ؗ'ls�q5�n�
��m�x�ַ����K�7Xuێ�E��q H����Uض��Vvv�=��R둛��n��Z����ۮT񒺢�Q�v��%^�W���)l���BB�C9v�hk\VN!7T�=[RuC�;�ؙ����@BJLpUJ]7dс�\� e���,W3�����3'E��I�R�s|�{]�������.�@�tE6��*�z("�1��qQҏ�k3y�:��Q'"Fn�o3d�..i{/���Q��ɷ9I��b��Gv+M��w1��X5'Bn8׵rb�t>�:��7<�۵�8�Y�x������x]��'d�3u�![+���u�vc2t����[�������V�]���.ޤ7S�\�vz���۬�.�ɸ�e�m�:��n6�����n�ڷ1�[r6�[���a�76���0ڌ�4M�Ie�nI�,�d�K��v�d��7rl��#�4bп�,i-rG�=z��֬��X6K��EEv���]�G&��u��>����u�����]����UU��� {m��u���s@���6y1��UZ�l��ޗ�n�ŀ{zb�-tJ��nc�%"jI�{��=oLX����L��TS)۴�œ����ey�-�I��h1kpT�p2`Jꂚb�Idm��c�D��=��, ��x��x޴FR�;������`{^,B�S
!$�Cn��޶h�]�բ㢉�ō���� }�� >�w��DDB��}� ����;wec�6�6��M ���옰�1`엀�T�G�h�N�www�nɋ ݓ n�x�,�>�	a<�� M�dI��ōݓp��\�9�ŞѸp�X���F������{��V���Z�7zb��/ =�^�����ș�X�c�M��޶h޶h�w4{��{�%cq�j�s3w57w�y��<����P�T/�>�w4�Y�}zPDMF�Ȗ9&���:BJw�|�o�`����٠_t¡��O蜎9$���s@7d�Ϥ�gLX���i��u�6�ݤ������u=�����ݎu�m��W(�,�]<f㖖�������x�IX옰L7���Ͱ���@�u�@�빠{��hz٠�ƮI��A�E$�@�� ��ŇBI)��u��u�^�3Cs9�c��{��hz٠{��܂���D�R���ٹ^��D�"ǓM����@>�/ ����#�X�t��n�Z����gm��h�yOg����Y��fBO�870�$�MI4�h�w4w]� �[4�q5o �$jG�{��h�[4�Z��T<x)���$��{��h�l�>]k�=�w4V�ʔO��nI��[4�Z�z����s@�A��ǌ�m�m'$�˺���%����7ذ�n�$�u�������ԝ�G�h���T��Vʶ�WGcr���WU9Q��k:K��#]Ow��u���Vn�@G���V�S�c���wK+u�U#��6���7d�vs�� B��3�~u�����89]ӹάB']��g�Rr�WRG:;7[��9�Eu9��m&�n<v�s*.�բ=�t��<]����Xz�xq�n��h\�0=�h蒌+�W������w������d���Q�rl��.ɥUmϐ�����nD��c�I�L��0�L������=�1`엀y�J�5o&�bT+���UTլ�o~���S!��xͿ���[��}z����cɎbI9��%���`�b�=�b�$�m��aN&���uz�n��[����@��.!��m�19NV�&,�&, ݒ�}Ұuӏ���k���ܲ�݇�]hѳh�ǩ;�)�U��_d��!%��ze�`�LX�%��J�6tŀzSd�AW!UwTU���w����c�"*UQ���@i�cHF������I����=:b�=Ę�L7����UQm���hW��=��hqn�{��{����a�#�=�n��$ŀ�^�t�V�n%B�*�T�Z�>ѼXD���Հ{���������x�#���4� u�s�p�u��I��[0Z*�%�.g �Ծ�T�U���� oIx�Ұ�1`qn�}bq�na�I8��h�����5�b�<��X�n��x�4�i��7#iǠ{���>���?d$�M}׀l������H��]�mɚ�[������z���բ�#�qr693@;����Xq&,XoDS����ݞ����s;��Y�ǃ��3�s���j�m����	21�1��FӒM��z�x��o%�N�V sj���V�4�q���hqn�W�z��X������ʷO�uk �b�*��@�^�{�����7�8bHNf�W�z����w4؆��%��<�o[��n�M��ԏ@�^�{����h{���O�co�W]:����b��l���V͹�v:7V}�@��L�	u�7c"J�nNFӏ@�빠}Ż�^��+���aP���9NI��YM�uz���բ�#�qr67�uz����;f�!��TU7UUuu��DD�s��;_b�>��0:%��_V ~�5�`9�d�8��YM�uz�����YIbj2Q��%�5� H	m;z��V9#�
��y,�cؗ��!�9ݓ����w<|ށ�q�u�t��ؠ�N��ۇup�'hƇi��qo ���IAò�x�\����l/m%�u�\-�v���S��G�n�]Ǝb]����>���P�;pXy��Y�5�u��l֎�ι�g��fG�r�Gn���g<�Y�њI�3.�ڦ��u`@�!�ԛ-�̚�Ѷ�k�3���y����j���]��F�M�&+��Q��Lx<I�?���k��3�����*�W�y^�@�빠}��{#�,p��&���]g�"!Dɳϫ �}� ��)�wtB�<�@���m8�+���w4���^�����Sn��������@�?OƁW����z�px�Ȝ�'$��K���\�Xޘ�	\݇�ۗjޮy���ݢ�׳�i�4g^���R=e��`�64��vY\��{Ұs�`zb�<�\0L5�E*(UE��U]]`��Y䒅�QP�B���X�]� s�u��*]�51B&H�@�빠}�e4
���]��b�cW	����5�ә�yt�`�J�5�J�&ɋ �H�d��A��
C@����uz����l���-r6�H���I1x�^�*9�����m�8�����nl�79�ob4�a$ BN6�z.���w4��M����X"'�dr6�x�1`R\0��`��g����4r)R.�sWusUv�.w� �}�7>}���Q�M�!3C����!�Q�K+)"��`@ @��(F�������Զ��Y-Hל���� 2Bnz��!3N������څ��t"�`�O4hJJ�d c���[e�Q)��\h�n�[p�f\3L�5VɁ*�&�iu�VT��%
Z����B���)sX�:�@��:R#�ۣMo�&sT�-	i��2����4K.�qw�� @ā-�%Yt1Ѵ3EmIYU����1�i�L�5�n�SZY�&�U������8n�؆h�тZkV댸��B��,�.h4H���"C�@��8y�$�Z��$$a�J@�ޛ��@�BIX���KJ���a� �g�ͺ�o��XĄc�$�(x $E8��@ؚD�O����Ъ>z����Q
,��v�{^,�
�k�x���Wuz/uz�]��)�{z�c�1�En8�^�Xޘ�-�=�X��D�ˊ�3ͫ����z]�:'�βtĵ��އ"�䋚�գ����J~m��?�q`[.�t�?%�^�m�t�^�mƪU?ȵG�T��:�X�o�d���n>��I%���J���f6��~���#�X�Xݡ��׼��~�1�����y��銱�ߖ���6ٵī����E�N3RIy���䒫��Ԓ_x�㜶��� �	���"�,b�v �x�����9�v�o����V<i�#����䒫��Ԓ_z߳�J���I%��[�%���cx6�K�7�]g�1*ٹ1��L���q����^s�:Q��v�<��Y��� }�o�;�m�]2�m���W����m�s�*��{����O��7#c�>�$��Ԓ[[ҽ�ۏ�*��{��^�m�貊��1��m��$�����IU�q�I��O/y��t�1�ۚ��e���v����n>��m�y{�n>�F��_�$���j�1�ѵ��s�[��s���E�}��m��w9�m�=�y7m��y�H!!�!��)"�>�nw��d�F���$�\�T��U/-[J��'+�61ض]l'\[7��V���0ld��l�=��G]�n�����v�q�m�g��5�p���[&��vf�W���/r�HS�Gg�k`%:�0�+��Ξ�f^��F�[�Uz��I�v�,vA:i6@`;�������z�y��`��B�n6GvN�3p���gc��;�㳦�;1%��A��{������/������-#&ټ�����iѝ�w���ק@O16ՉFKV�#�P��$)�Ir������W��%_]f���i��${�W"�Ńj6�f����W��%W]ǢI{��o�%_]f��]�`��mC#��#�6ܮ�F6�ݏ!�6�}1V6��ޕ��%z@�6 �q7#5$��]���qɊ������y��t�1��ɔ\�Á�,���>�$���$��3�_~�^�7��~�1�ߴ�y�ܟ7��W	;�J\���6:�ܬ�5�*ܾ�8�a"EîYv�����HVn�m���W��r��1�ߴ�y��1�I%}�N�X�m�����IWn�o��(J����Q�@�����
@���P!V$�YHT�"D�f�n���g9m����ݶ_3Ͼ�s�����^�FGY�S+�V�m����6ܩ1V���W��q۸�$/�n'�N$�
C~B��~�߽F6���߫�m���X�o�L���G>��$m��q��K�ֿ�m��±�ߴ�y��I�cm�Z��,y{<���3��	��2>�u��c�[t���<ɗ��5'$��fN�-f�n��ێ\+m�c�{ͷ*L�m�m��J�px�#$�&�����q�}�(J����(ə�u����3.]��$����O�d�Q`�m����%]�Ͷ��y���]�m���~�k零��-��$���\[�f(�M8�5%����^���[oouٛ���>��s�ނ~߿��� ���w��KԔ�~ �
��~���mʓ(��}[%{͇���}������9.ێk p���;(sA�u���:�n.ٻ<�uY.�;Җk���$��[O�I*��jI.~���IUe�����H����`�R|�U۬Ԓ\�W��%U�z�K�i��$s�YI"@�m�ӌԒ\�W�m�R�<m��!�6�rb�m����!Ơ�P��4�ߒJ�(�$��VC�m�Re��_�|��Ε�6ܕapx�"9M�=I%�U��䒮ܣm�N��6�u#�m���&�m�ϏN�%ͻ=�3�U�c���[<i� ���/f�&�dؖ����l��������Q����J��n:��6��G���oU\[��3q��q��K�����6�nw�7m�ϧw��[o���ɾ������{�h���W���� ���� ���>�z�U]O������}_}32)����P�H�������䒯���m�g���巨�gs_v����z\�h��
`Ф>�$��Ԓ^w���ێ�:��~�d=����lȪ�wMXT���I:.��L�J�8��'��:�ip����#u�{>׻\ۓ�zA��۶��Wa��\�Λ�lE��������w73�C�h�s����*�	��`�n�Wjuq��EY	��#��mq<� qǵ9�]s�5V�P�{('vk�[ͬnݜ�3�P���k�U�`�۞8��<d�����%�v�����zH����'ns=���v~|p���8�ĄM�+HΆ��k^/.���KM�k<6�I��j6*x���VU�� ��~����G�SԒ_qv�|�U��jI%��q��y"�$i���%SꞤ�����䒯��RI/^��Jٓ.6<��#��Ԓ_qv�|�U��j_����m��O�����? ���~��u�6Z\���nWL�m��/�m�룬m��&C�K�î-��6����f��^�o�m�룬m��&C�m�]2�m���~�t���8�7>�m�&�WI��k
�4��K�r�s6D��槮j�-��'�$�O�z�K�.��J���I$�zϾI#��p���21�Ԓ_t�NpzD�E�$F1�1"��aE�BAc#@* U��HD���(
0`�`�@���*���w��RI+��}�IT���$��o�CF��Ф>�$��ԒK׬���%�u��S��hq²<M�#M��s4׬�*�^���j�-빠�`���ǎ,q����ڴ�;V���s@=z��`�-l����<g]:۔����M�k�19��'�4����p��7D�X�ccɈ�r8&��;̵��w4׬�>�ՠ^n��@�U]�J���x��D�o>��]Ӏr�Z���n-��1����� ��xΛ��	dD�I����o _gc�'&A8�y�M��ZyT� �� 6t� ]����Gõ`�f�� �*np��6������>�ՠp�����$���RF����v�r1�cni���eq��L�kK��;,e9�!�H�bG���s@=z���Z{�@=N+�blAm�ۙ��f��v���^���s@;��E���ɠ}]�@�2נwu��^�@�recS&% �pM��7�7X�X��<���F$����VDX$y�>��I9�ٟ@�@Qr!�@�빠��@�WG��K�7B\Cj��t��&ܽ6����=c4{v�4RZC��a,��n���>v�)��c���MI��[4����f��빠�Ȝ�q�Ȣ�xε�I��]׀=}� =�� j�"-Q��X&�U� �R^�����^��}V���*ka"�2B!I�Wx��� ����>u�p:guw^�{�O�E��i�nf���^��!%�g~� 6�~�}� �R���c���S	Ow@4B;4�o\�˺�&a���wWf����iw!ؐ`�b�bƙ��ܑ�.4f�\�BB1��g7�S	r]�֝l��8���%L֘bJ�w�a.1/��	$	��F����.q�K�)v�1��r�h`ؚ�&	���zټ4��|�IsD��XS5��X�����\4����&��4�ݢ����Z	i��L8xx���"&�HIvB��)�Vа֎Blƙ����!D�V4 F
��hX%0��H���������[���0ơ$f�r���t�nS	SQ�u���l�)R�E������RL�t�.F�C`E�$�	B2h7���JksI����1�e1e�.��.�\�҆�9�!	W����wv�!�}��o�-���  ��7h�w����f���rݐ�vӵ(�  m�m�	 -���      �  ��m�� P,�Y�s����:��v�����R�m�7�~|U۪�b����K9G9��Nk$�L���lmuA�ՙ�f啩I4p��x�I�=<�En��q�����%Xv�ݠשĔ�s�i��u���z��x��ۮ� �\v���q�O �f��
Ǒ�n��Ke{"�f9jG�{>�$y�NU��ݖ���;J!F�p m�i��s��1Ė�Nm���=q�t�����=��g���a�65���qpI�!�9^xα�<9KnWq�8�����s��Vێ:�.�\�;=,K8���=%�#,����n�v��W K�W,��Ȧk�n89�
;	M�>ݽ�a�`,v*C���Ož*�|$��Rzv������U�W,�#!ʲ��J�U����+UX.�ێ��T���\h�u�icb��-�eZ�*UP�m��RͣQ�C�����i����[���&���,�P�Z�P8	;t���ڂuU�um��p������"��6���;N��L�讋��Y#�޼�G7m�g���3�ʭ��C\���{C�[��DN����I��97Lʴ��H�ְ�E��뮮�nۮU��峻W�:��XC�	=��&�����]h)�|aq�t��[� qͳ.Fq���jԵq�vS	���\F8�`Ckztl�]izp�Ѣn�G='!�L��s0j���D�����+������)��l�hz��hfT����&�1$�:���x$l ��yTݖڻ`ҵ��ze��H�]�Iv��1��V�Pk��6<=�;�|7awfw^@��s�"�[�Uw9�ڶ����Y�5P�Z�p*<�[��U�^���m0�s:������\�=�����J�9}Yӱh�9��|n�R;=b��{����w{�p�TG�h�T(�(�PM�D�*�<Cb*�u��䄏6]�k&�j�Wf�e[x�܍��;��n�]3��Q�g��)��J�m���w^mM�15���uy��m�sg�Wc&�8~����-ֶЎ󵪭el�N�[lj���(��mq<�ێg�F*�u��2��ֺ:��	����5��x�1H��n����(�v�t���ey�8��c]��n��V,C9N�����*��U��wwn����>�Z��n��d�� �^h^�7K9Ă�՟h�K��}���o�7�匑ӞwLJ��m��ߧ̓�M��׋������9�#����̃��9�{�l�ؑz���9w��@���@>��Dɉ�@�sŀz|�a�>�}8��� ��6����������X;[�X��N {�٠w��h��6�#q$���:�8)�]��_b�=>n�M���8,����gb���X9h�K/
�u�5�n�
q���*0ݑ.z����.��� n�/ �� ײV�]��<��*�v�U���-/��I� �YXBPd#FA �d(X�,A*5�ɡ:s��{���'�뽻ND�,K����iȟ�0���������L��+
������K��>��6��bX�'�k�ݧ"X�%�}��u��Kı<����r%��{��>���c$q;;�%g��{�K���}۴�Kı/���bX�'�}�ND�,���ͧ#���ow߷�o�3��l4|�~o%�b_};�m9ı,O>��6��bX�'��{�ND�,Kϵ�nӒ���$.a��4%"�]�6�R���=��מ��Ϯ{%l���^���V=�тZ۱�.����p�kiȖ%�by����Kı=�{��r%�bX�}��v��2%�b_�?~�ӑ,K���Oߎd�������Z6��bX�'��{�N@lK���}۴�Kı/���bX�'�}�ND�,x�����'�C��)�����{��'�k�ݧ"X�%�}��u��K�U��z
��
` �$r&�k��8m9ı,O��߳iȖ%�bS��'I��.�[n���K�lK�{��"X�%���w�ӑ,K��=�siȖ%��6'�}�&���t��+�UvL�ͪ�� �����pI/�}�Nı,KϾ�6��bX�%����iȖ%�bw�;���%�#F�O�â9܇:�1+GgL�i�������+{59�Ge۴��捧"X�%��{��ӑ,K���ͧ"X�%�}��u��Kı^o�Y����$)���*nT�
�WY���r%�bX�{�y��[ı/���bX�'���6��bX�'��{�NEı>�]'rf�j˭Me�s5��Kı/���bX�'���6��c�"�C"dN�߿fӑ,K����ͧ"X�%�|�s;�	u%Փ5��m9ĳ�*�E2'����iȖ%�bw>��6��bX�'���m9İ4�cꆄL@t �b\��u��Kı<=���035s53Yn�m9ı,O���6��bX�(�{�siȖ%�b_{��m9ı,O;�xm9ı����1�x��\��<ڹm�������e�p�hJ*郷C�e*D��vjNJ�պ�Z˭fӑ,K��=�siȖ%�b_{��m9ı,O{�xlyı,O���6��bX�%;��t�j2�P����m9ı,K�~;�� "X�%��~��"X�%��{��ӑ,K��=�si�
ؖ%���Nܹ�SQ�kRK���ӑ,K���w�ӑ,K��=�siȖ%�b}�����Kı/���bX�%����kT�1����\��iȖ%��b)�;��~ͧ"X�%����ٴ�Kı/���bX�X�����K=���~����8��tĬ��~oqı>�����KİV�ߎ�iȖ%�b}���ӑ,K��=�siȖ%�b~?~�m��ճ)���5u�$�.� $�����Λ�����p����cs��)]����gtm��kz{21\�Hv�<�6ɮNC=���n��Y�`öĩyf(j����;�;2x���mt�mH�Qj�}�ݸݚ�'
�9��L�$n���¹�gy�0gl�=� n���읳A�1�cZ.�Q��y6u㭣Y�wϛ_5�\[�;F��n�'F�ㇲ��ѻ�\A�,��N���b��Z痌��IҮ����`
�U��g��Kı/���r%�bX�w���Kı>�{���O"dK��~��6��bX�%����ڐ�D�0�kD�k[ND�,K���6����bX�g��m9ı,O���m9ı,Os�ͧ"X�%����t�I������ˬѴ�Kı>�{��r%�bX�g{��r%��F
"}��~ͧ"X�%��߿p�r%�b]�?��/�;L@ORS�������6'���6��bX�'�ߎ�ӑ,K��{�ND�,T�>�{��r%�bX����1�%֡3Z�m9ı,Os�ͧ"X�%����6��bX�'��{�ND�,K���6��c������c��KܝKN�.v�D�*������1��L�F�R���(ߝ��t#�4Ff�$�Y�Y��%�bX�����"X�%��{��ӑ,K��;���9ı,Os�ͧ"X�%�~�}:���bQ�n�����{��7�����v��UR�"8Ȗ%���{�ND�,K���siȖ%�bw�w�ӑ?�"DȖ'�v��i��)��Y����m9ı,O����iȖ%�b{���m9��"�S"dO߻��ӑ,K��}��m9ı,N������j�Y�����{��7�������r%�bX�����Kı>�{��r%�` X�����r%�bX���3���f�f��.ͧ"X�%����ND�,KW���ͧ"X�%����ͧ"X�%��{���r%�c���|{q�
�'��X�r�6�����Q��ac
:.y��ͤ��r�s����.�f�je֍�"X�%��{��ӑ,K��w��ӑ,K��=��lyı,N����r%�bX���3���.�j[�5���m9ı,N�~�m9�@��,O����m9ı,O߻��ӑ,K��=�siȖ%�d)zÑV D݈RU��B��$)!H��{�ND�,K���6��c���E_��dN�y�6��bX�'���ٴ�Kı<��.sQ�	�Ԓ�hֳiȖ%�Ƞ�Q�����߿�6��bX�'s��ٴ�Kı;�����K��A��|~��ND�.��~����hyS�Q�n�����{�K���ͧ"X�%������ٴ�%�bX�g��ٴ�Kı;߻�iȖ%�b|z}gy�[�a��f���� F,墷%�뱋��V{���m7gb��9/��y~�l��:bV~{�7���{���w��ӑ,K��=;��r%�bX�����Kı=�{��r%�bX�����뙂��g��{��7��=�N�6�����:���'����ND�,K�����r%�bX�����r'�Tr&D�/��f~Ԇ��h�kZ&�m9ı,O߻��ӑ,K��=�siȖ%�bw;�siȖ%�b_};�m9ı,O���2L�e�[��Z6��bX�Eȟk�߳iȖ%�b~����ND�,K����iȖ%����HE��db�$��d"�H�V�JB�F+��#	H�,���E6(!�O�����6��bX�%���2��YX؞����{��7��������9ı,K�{��"X�%����ND�,K���ͧ"X�%�ﺓ��f.ɴa����Ń<��{S�
�Ѷɍ��ҽ��[�3vy[�{���������E�lV�Y�kY��%�bX��ߵ��Kı;߻�iȖ%�b{�������&D�,O����iȖ%�b{�O�.sZ���jIu�5�m9ı,N����r�G"dK�����r%�bX���fӑ,Kľ�}�m9�A�"ŝou��������)W�Q�n����bX�'�����r%�bX�����r%�bX��O���"X�%����6��bX�'�}{��52Rh����3Y��K�O� �L��_�~ͧ"X�%�~���m9ı,N����K��D$r'�����r%�bX���ݿ�ffj�����7���{����ӑ,K��{�ND�,K���ͧ"X�%���{�ND�,K
���"JB�K	BD�U!
6�F�X�H� �B��4�����֦�r�ΒD��6킂����y�Dd��Bv6rqǎ�,��s��&���=kǧY
f�a����62�w��m������A�l�:N�hS��`�m�niJ
Pz��P���&�2F�sYNH����=&r�r6I�x;�Nn^�-sv�r�:�����<�m/M�n�����[��y�\�Îug�n�I�)M��gc�e��p� �{@
�ǧm-ͻ=�#qæy|�M����i��ї�g/k�O����V ę���jCZ&)�֦֍��,K������"X�%��{��ӑ,K��w��ӑ,K������r%�bX�?}��I�Lչ�u2�Fӑ,K��=�si�� ��&�j%���߿�iȖ%�bw���ND�,K���6����(A	�2{��?߿�?��lOJS������,O����iȖ%�b{��xm9ı,N����r%�bX�g��m9ı,K��I�Z	��j�Z�fӑ,K?�
�� �5�?zm9ı,O����ND�,K���ͧ"X���R�������r%�bX�w��r�5��MkT�asFӑ,K��{�ND�,K���ͧ"X�%���{�ND�,K�O��i�����w��߻��c�Ϛ�L��8fgi�&�<�Om=�GPt��I��ŝ=�����w�{�w�_/��(�,�*������{��'���ٴ�Kı;��siȖ%�b{��xm9ı,N����Kı=�����ɩ�����3Y��Kı;��si�_�2��t%�`8�%�`Vd�L�)���f�@`a�r�
G �b�-��B�2�.fB�p�2� �eė�	c�6�`��	�� ��� ,���&�{�iȖ%�b~���ND�,K���ͧ"���\��,O����L���-?=ߛ�oq���}����6��bX�'{���r%���"dOs��fӑ,K����~ͧ"X�%�|�nwR�0�Lֵ0ִm9ı � ����߼6��bX�'���ٴ�Kı;��siȖ%���"}�g��"X�%����/c�5nj�L�Ѵ�Kı<ϻ��r%�bX�@H�?k��ٴ�%�bX�}���ӑ,K��{�ND�,K쓿������S�*���=�92q֔�P�\�ݝ���<^D�a칩�U�lOJZͧ"X�%���{�ND�,K߾;�iȖ%�bw�����L�bX���߳iȖ%�b^��?�&[��!f��ͧ"X�%�����U?1��,O߿~��Kı=�߿fӑ,K��w�ͧ"X�%����s��d&��K&�iȖ%�bw���"X�%��w�ͧ"X�|�i0��/��6��n��춐$n9r��ə��M7�eM1�.
`g��W�4Z-(��35�#<BbK�JϜzBT�l<<=��e֒\�K��B�L�<'Z4#	sI.F��A��a �V�5��
�i��mOX	�{�RasF�\�K���)���e�4��sL�ŗhA p߿$$�\N��HF�HJ\�0�t����e�s�u&3
]o�2�"Xa=���4m"'R=��$$ֵ��ֳ>t�.36���ˋ3b��Q��2RP��e�ƥ�	&5����KA��j���GC�eTSGh�T�6�����������h1��T��1�>��~��Kı?}���iȖ%�b_����ճ2a��˚��Ѵ�K��H�~��6��bX�'����m9ı,O����"X�(�ȟ�~���Kı;ޟ?���������{��7���{�ND�,K�;�iȖ%�b}���ӑ,K��;��ӑ,K�����~����䞒�N��u�N��1��1Qs'u�tb��e��1ɬ�K��Q��\����fF��i���oq���������ND�,K���6��bX�'���6��@D�!�MD�,O����6��bX�%�����Hf��E3Y�Z5�iȖ%�b{���ӑ,K��;��ӑ,K��>�siȖ%�b}��xm9G�ș����/c�5nj�2]h�r%�bX���߳iȖ%�b}�w���Kı>��6��bX�'��xm9ı,K��2�5�����]a��f�iȖ%�!�H����ٴ�Kı;ޟ�m9ı,O{���r%�`z�� #G$Os��m9ı,K�~�z]2L���,�ֳiȖ%�b}��xm9ı,Q?R#�߿xm<�bX�'�����r%�bX�g��m9ı,O�?ݿ���]��y�%u��zN�5�I utۛ<��3���.����{���ۿ>]�G�5�K&�i�Kı;����iȖ%�by��siȖ%�b}�w���Kı>��6��bX�%��;�[3&�̹���6��bX�%��/䉑2%����ٴ�Kı;�ߎND�,K���6��bX�'��w�nM\��Zj��\ֶ��bX�'��{�ND�,K����"X��`c�2'߿~��Kı/~����7���{��������jsSP��ND�,K����"X�%��{�ND�,K���[ND�,?D0ȝ�~ͧ"X�%�}�۟�I��f�f�Eֵ&ӑ,K�����"X�%�~�{��"X�%��}��ӑ,K����K��Kı >��a(�
B{��֦���0�c��n�v�i0I���2H��7KR�O<�Ś�$q���Ɛz��s������S���s���N:����7�'��g)q�Oe��������}1��:Fw�n�,�r]��yD��xҋv����ܜ�];��<�n(,�p�ݮ6RH��v�æf��q��f��Zێ.V!�y�ׂ�^{ ۧ�3����R�g4p��/���=�w|�7���6T���K��|��݊�zs�%(�!�՚��L֩��&��a���k�p�!�eԹ���u���Kı/�߿���Kı>ϻ��r%�bX�w]�v��bX�'���6��bX�%�ݙz�B���,��w���oq��_����9O���,N�����r%�bX�~��ND�,K���[ND�"��5Q,K�����]0�5uHY��fӑ,K�������9ı,O{�xm9ı,K�{�m9ı,O���6��bX�'�|v��kT���BYu�.ӑ,K[���ND�,K���[ND�,K���ͧ"X�%��uޗo~oq����~�;~�1+w��Kı/�w��r%�bX ������Kı=���9ı,O{�xm9ı,N�e���d��5�]K�sI'\a�<6��f�]:����q�p�7W[n�\�7P�ه�tA-|�~oq������{�ND�,K���3iȖ%�b{߻�h�"X�%�}���ӑ,K7�������jsSP���~oq���b{�w�m9
#� �D+�Qڨ�Gl�bX�~��ND�,K����ӑ,K��=�siȟ���DȖ'��]��$���.�j��ӑ,K���p�r%�bX�߻�m9��C"dN�߿fӑ,K�����r%�bX�?}�L��3X\��d�h�r%�d�*ȟw��&��	���ٱ$D�߾4��H��{߻�i�����}�߹?V��^����%�bX�g��m9ı,?$A����=�bX�'����6��bX�%���[ND�,K�>�'u1�z���������h�^p.���g�W)�\pnu���l乧%������O�����bX�w��ND�,K�}�ND�,K��{���@��&D�,O���ٴ�Kı=�����kT!��%�᭧"X�%�߾��"X�%�}���ӑ,K��{��ӑ,K�����Ӑ@��"dK���~֭�s33WWZ��Ѵ�Kı/���[ND�,K��{�ND����B�"{�w�m9ı,N��xm9ı,O�����jkW	2j��fk[ND�,O�AL��_~��ND�,K����m9ı,N��xm9ı,K����oq�߿���멨Jj����x�,K���3iȖ%�`��b�������%�bX������"X�%����ͧ"X�%�ߤ���nX&)8�<v�ޱ�n��^�\m7�7.�3n�|��u���5�f�\�Wg��{��,N����r%�bX�߻�m9ı,N�~�l?��*?�E}���%�����fӑ,K����r�e)�5K���5�6��bX�%���[ND�,K�߻�ND�,K�����r%�bX����� �@AY��,K�ߩ3��]Rjə��.���"X�%��?w�m9ı,Os�3iȖ%�bw�w�ӑ,K��>�siȖ%�b_��e�t�2�ꐳZ�fӑ,KP�����r%�bX�����Kı=ϻ��r%�`hȐ F)��D�$DT�b���߻�ND�,K�~칙�j�3Z��WZ���Kı;߻�iȖ%�b '��{�ND�,K�߻�ND�,K�����r%�bX�}'d���Ƒ�����y�u�s7\Qt\I�g���3��g nJ��Bv�6^WNe[�'"X�%��}��ӑ,K��w��ӑ,K��>��6��y"X�'����iȖ%�bw��ܲ����̺����fӑ,K��w��ӑ,K��>��6��bX�'{�xm9ı,Os��6������dL�b~�_��:sXi������7���{�����ND�,K���6��bX�'��{�ND�,K�߻�ND�,K����&h�Fu��Z���K���dO߻��iȖ%�b}���6��bX�%�~�bX�'��ݙ��Kı=~���R�ɨ\���Ѵ�Kı=ϻ��r%�bX����������,K��;��6��bX�'{�xm9ı,LAC�ݽ�m�&I�W5��$�v�n F�N�}'���p�5�3�$D;P.̈́�Ƀw;M��Ӽq��m�ֽdb�p:��<�v���<v�r�U.���;�q �j[t�jUU��.��!E��\���'�$������L��y�_ ����Ǝ۳�c����q跆���S����l�lg�����&0ػ*ⅶWN��,��{XΑ��ԍ�\s��ʕ\��=�8N�!���۴#��V㴘�uH�r�ٳ�4��W.��'�,KĿ�w����bX�'��ݙ��Kı;߻�h#Ȗ%�b_~�u��Kı/�}2�ӄ�uuH]]f���Kı=Ͼ�ͧ"X�%����ND�,K��{��"X�%�{߻�� ؖ%���s���jIlֵ.ӑ,K��~��"X�%�}���ӑ,KĽ���ӑ,K���}�v��bX�%��;A�E+2��=ߛ�oq������93�����"X�%�~��m9ı,O~�ݗiȖ%��@&D����6��bX�'~���)��ui2���35�ND�,K��w[ND�,K�����r%�bX�����Kı=ϻ��r%�bX��O��%0�2I��ɭ]a�	�8a�`���ilF��z��d���l$�WOK��1,�CU�������ow����fӑ,K���w�ӑ,K��>�sb	Ȗ%�b^���iȖ%�b_;۝�$���.�]kS6��bX�'~��6��U�"�vРx�mș��s�ͧ"X�%�{���ӑ,K��>��6��bX�'��ܽ�\�5���5�6��bX�'��{�ND�,K���[ND��C"dO���3iȖ%�b~�p�r%�bX����;2kP��fa��Zͧ"X�%�{�{��"X�%��}�fm9ı,N��xm9İA,Os��6��bX�%��^�q�5uH][�kiȖ%�b{�}ٛND�,K�}�ND�,K��{��"X�%�{�{��"X�%���Bo���.��WZ�ֹ�;�YȞ�:3ȝ��#��s��N�kWeF����5Џ�;�klY�����{��7���xm9ı,K���bX�%��bX�'��ݙ��Kĳ�~�;��¹V敻��{��7��}���ӑTlKĽ���ӑ,K��=��6��bX�'~��6��bX�'��{8S5���L�պ�ֶ��bX�%��bX�'����m9�f�*�J��k���e��!���J���J��#V%�T�	IB��a(�����XYP���e	vx�P�9�s�6��bX�%�}y����$.��깚�.n�j��5�kiȖ%�b{��fӑ,K���w�ӑ,Kľ���iȖ%�bOou�/�RB���Ϧ��a7ASvfkY�ND�,K�}�ND�,KT����iȖ%�b^���iȖ%�b{��fӑ,KĽ���/m��:A�'\3���v����G[-m�yu��V]���r�y��1��n�����x�,K���bX�%��bX�'����lAD�,K�}�Noq����}��;?���;9ҕ|�r%�bX�����r%�bX�������Kı;����Kı/�w��r"bX�%��^�p�5�XB��k[ND�,K�u��m9ı,N��xm9ı,K���bX�%��bX�'��v��f�S3D�浬ͧ"X�~Qb�9�{��iȖ%�b^���m9ı,K�{�m9İ>_  �
iR'�k}�߻�{��7������ߥ&ni[���bX�%���[ND�,K� ED3�߿ki�Kı>�]����Kı;����Kı<~>��ԭ͞[�+rv�6�>V[��V�����u��`{]��o]͞H!��Ÿ͠��{�7�ı,K�{�m9ı,O}�}˴�Kı;����Kı/�w��r<oq���~�oݿX��`j�����ı,O~�}�i�
�%�bw��iȖ%�b_~�u��Kı/}�u�w���oq�����m�V��%QI��Kı;����Kı/��u��Kı/}�u��Kı>���.ӑ,K�������ɓP���3Y�iȖ%����3�߿kiȖ%�b_�~���"X�%���o�v��bX(��߾��"X�%�{��gff��\�5�u�m9ı,K�{�m9ı,? {��~��yı,O���ND�,K���[ND�,K�<>X�1K�����QT��+b��F��Ė��#"F�"��>�7�.K�! M��	C$#p�2) ��{�L#��d8��I$ad �a�٧͙.0��dI ����}�oo��m  U�g�u����t�r8Y�r�]iv.C���9�� h � �       �  �  p  �zz��u�^�;K�U݆�Џkt�Y`�[n��YUƚVVb�A*�r� =b����IгZXib՛[ȫR���i6��^��*�jk��ayv`hM��v�gbl��;)pvl��z�5��Q�E����wn;A ���{�gS�kb��S�Aw	��ֺ�IH^�d9��"-�s���F�s�뇒���<ڇ�$�qρ��\��<
H�;�즠��͎p5�%�'=�����Yz|�Y���GH�oi�q�����6-i��\�܊=��/[��%���ɸ���r�;B9 �k�Y{-�x�õ��,�N�۞8}v��k/�t�ŋ�%�<a�2v�$�m�jj�U	�p��-�����W�V��ȉ`;i��������/T��Y����Z��4-\�H;��AT�Ij��NԭW�T��V2�F�s$��U�������U����1u]����I�ѷPC��Ymv�r۪΋l��݃�Vԛ��m�s�{h%;cve�r�ͺ����g�kA���cv�c4��AY��C�L�`�K�uɎ7M�&�qd�M�y�#;�j�8��61��zQ��S����v���evR�Vz���7v�gu�e�q�s�;=�I�HkyTӜu�!vDݐ.�c�S���`���s��6���'/^"�l�r�N�qF79l5!l��1��U2�m���:�K��s�ꓓk��^;tRZ�J��G��ԧ4�;�{c��.{�x7��vX���e�q��� �.^ɱ�&��J�k���rv�-��=7qnӻ����=rJ�X�f[.DUm1��
�9��)MT=��j�����`(�]Ur�0)������1�S"v�.��Cq�lvQ�Z�de�q�k��֛I����"���!�����U�Q�:�Ox��'�D3;�������i9���ma5O-UR�m*瀸�m�J[	�l꧎P�wm�T����1Ƚe���z��.���5�6�Gy��ɸݱ2���a�=��%uαnnU^<c�q���Z�UO5��sn!����U��M҃x�X�i�A���6��M�pэ�g���c�5��Ԛ���sL9��#)�;V���x�t����؛����j�d��=��;�tV������'myk:F��wc��i��v���j��^}�'�U��D�,K�����r%�bX�����r%�bX����؂�bX�%��bX�'��N����34IL��]�"X�%�߾��"X�%�~�{��"X�%�{�{��"X�%����r�9�"DD2&D�/��?k5�%��s4f��4m9ı,K�߿kiȖ%�b_��u��Kı>���]�"X�%��~��"X�%��{{8S5�ɨ\�չ��m9ĳ�$"g~��[ND�,K�����9ı,O{�xm9ı,K�~�g���{��oݿX��p-f���{��%����۴�Kı=����Kı/{�u��Kı/����r%�bX�ϙzR��r�)�,5sFk(VF�3hm�ٞMe����[/�/!rF̟=���ɬ�E�]T�7eڻ2�)!I
H[ϼ6��bX�%�~�bX�%���[ND�,K��o�iȖ%�b|���{�ɓP���ɬѴ�Kı/����r�%�Q�2YW��5`@#X"�cR�R��0�(V$��B)!�E6)� .DȖ%��[ND�,K���fӑ,K���w�ӑ,KĽ��g��wt%?=ߛ�oq�����bX�'���fӑ,���w�ӑ,K��;�siȖ%�b^������[�!un���"X�%������r%�bX�����r%�bX�g~�m9ı,K���bX�'��N���XL�S,֦ӑ,K���w�ӑ,K�P�;�siȖ%�b_��u��Kı>����ND��oq��}����e����L�r�����+�2���A�ۘ�Wm�������Q5�틖fk&��4m9ı,O��w6��bX�%���[ND�,K�{�۰@�
HRD�{�X>�1MU%�MYsUUu��/ ���=�b�9Ε�n�qD�ncM�9$�;�*��n��~=>�Y(��%`4��b �L4J�0#W��'D�˾���O~��ܒ}jvmI#�-�b�~��hy�`���?%���p���E5���nE&h��@=�@�YZ�>�����`&�biF%&Fړ.�n��xN�횎5�t{%qƹ����<�Gf���#F�jG�u�4����[��DD/��u`�T�ڒUM�t�6�����<�&,���w������J"����T⛕"*�����_������/uzy�o@�:ՂqT����n�`t$����g_V��uX(P�TDD$�7� ~�f)���8D�q�^����ށ����=-��?DD$�Q"UTjf�]�zu�=��!*^y5+F��ۺ��ҩl�|��?�{ٓ\�\Q4ۘ�r5$~���z�����/uz���L�C������>�x��BS&�wV��� �����	U�k!�Ȝ�L�<���kޕ�sގ�l��H�PUWb�J�������Jv��`u������<��@:��S�,n
<19X=�� �I� �$�_t���P��+�(B�JP��l���w���r�Vw\�����v��Z��ve�V����k����Q˻8(۳�mz�n�L��F;�E�l��{R�]��9���m���9�]�u��Br�v��#���7X0����]�璶N�A��+9[8�:�Wg>�=�nݰ[Ge
[c(���v:�p��:lu��<qͰuζ��I���Z�k���s���GM�v���t��C.������'� '�b���*B ������o�˵T���F��:Nڶ�-�7-Bh%q��r�5�3�,e6y.#��vҮ���b�=-��=;�����z�O@�����N`��dJ9�����!B�6[�����o ���Rɍ�x�"Q7���^���Sӿ���� Vנ{�9��lm&�m@����sX���m��Q
'i�� ������ɑ�5$q���������wW�l�Հl�\����%M\c�1_d����J\/bg:�:���n����7��6ĢYN�$����.��^ꞁ�[��Ճ��(S2��ֳrI�����;U��.$.Q
%ξ��7{�`��`�*K?����M����}m����(P�v{���׀}婪�WR�V�d�'�}m��<��@;������U�-Bs���ȣs4+k�9$����ξ��>m��6t�g\��͍Y����ٻ[�F��Nl�<v9.=�7i���\�7Q��Қ8�,�wK�9�GX���rJ�;z���ɪ��u5vM]���sY�(Q�"!%To�߱`w���w�ni�+����*nk ��� ��u��!/%B!#��!� E$ ��K�D(0w�xOwM`�vL�ET�һ���X�%;\���׀lP�)�w|���T��Wb�J�������w�~J"�ί��wb�<�J�5pbnʢ��-ں���|^8�p��39�.��څ6@h�7�e*�"朄��x�#Ŋ(��
�?=�n��^�wu����܍�N`<�EXͼY�����(�����X�߯ �ީ�e�N`$�6�E��y^� 7u��L���`��X��1Sɍ�x�"Q9�wu���M���7%T|"�Q�)�޾�y�wt�ȣM�di�'$���4�P���/��o� 7u� ט[MN��4O�<��9�3d����q���2�Q��Eۅ9Gu�\�!��Y��+���� �w]`ۮ�G���V��ɞ�MJ�U*�����n��ID~I%T��������^, ײ�\�Uq"�mFӓ@>�@���hw]��mz�\h��m�H�b��h~���]����6Oذ=�������*x��"��IT��� �u��?%�Qo����~�Mػ��9z�vA�#Ƚ�����vj�U��]@����e��g�=ڝ�n�]����ݰcv��s�׮����5�Xˣl&�Ƒ�����.�)�[��u�^뉯MW�`�`��'p�J��@��B3�����;���3�գ��#�:-n�N83�k��3�F�@ݤǌ\����i��Q�R��<p�>9]�Z޲a��gf���/wp�l�Wm#@I�<�kun����.��#��,frI�f.�l7m��ҷuV�>�����O�V�� �ʛ��&��9�����7����	~P��uߧ ��ذ�����E�,#24�#�h�t���u��>^����h�L�28���H�fB�-�|�N�V y�x����/�X%V	��7�6���|�k�I/ ղb�;�ŀN�n*U���s�]5�mӷ\W��m��;WK;tg��.��v�������W���r7�㤄g�m���׀y=x���`>n�wUH�̚���]K�krO��f�D�(u�XηX���D%2n��T��nb����߷4^����@�^��,�('?�<m�$I����IG�J*���x �~�x�׋ �o3@��M���J��I���T� � v�xZ�L��
UΙJ'�w:�-�*���4-��a뉺�݄��m+�;�~Ο�i���I��}� ��� 7�� {[��ͧ`����ԏ�4u��޶h���<��Y�2tuqԫR����`���kw����&��EL,���LI�D$�¡ �Zd		A�P"DT�H0�#I �$����߆�"bD	C.i�3F��S3n\	xdIh[�[��	�h��4�`��k&nf�.�e�K�f�#�� ��@����3[4��	u�f��C3X]������4J��D*��3[ĔaN
g��U�4�83�aSUr0�U5��bk�#B��.T�R���B!�R"D�y��hь�J��M�Z�4f)�.0�$��5�k�5��#5��A����.�+7ҁ�V�,$�%��H$@  @��@���R�B���S��V�|E�h�D"�Ȩ| ����* S��(�~D��� 'ȏS{� {y�q�uj��S�� ��x�׋ ����)��׀�Ə����Mą$�=��s@�[����@=�����&8�c=K\����r�����n�3ήl��x�[�;N*N�ʧǍ�d��s�6�|_߷4�n�����_Hj��X�عM\<m�!����@=����w4u��ו7�L��DrM �Wx��ŇD)�}ذw���hwi`�
'�@�{���s@>�w��(P���P�A�n�76���-Z�*n�V�kx��J}�����^�zb�ߛ�N6�:m]P`�:��捬V�lw]����S1�e�s���/\�K�@��&��8��� ��� �Yx�� ޓ wsT�T��	������ ��yДL���X��X�[4�cE��7NPRM��u`��a�P�O>��}׀{�S�qkE��fa34nN�)�>����O{���kw�yn�X��Sqq5D�j����kw�~�
u�_�jo�`��nH�� D�&)�����nK���k@UUUmUm*�{\��	s]C��ri'�^�MƂ7v͢Z�N;N�2���*�jnz���d�6������ٻA����r�SxnP�9F��r��ă��f�6��u3BI`�����]K����H�0g>�ƃo\R9��/t]�E�KF:�t��=F��ƭN�Sw]�Pˎ��F�.
���V��2�Bd�̹�3D�f�>AOY�j_�5���Och��d���*5�}Ơ]l� ]y�x������[�-��6�j�m��׀y{^,��, ������M6�di�G$�=�빠{��������ΈJd���
mZ�4T��.�`��`�n����^׋ �Յ���cx��4�[4�l�<��$����`�*��TݐFӓ@=���:�h�w4�u����5"�F8�DR��y6�P���5v흻bv��.ꋳ�7&V����n�M�Ww�n�1`�b�oK��$�(^�~�xk��'ܠ���.���rO=���C�� H���Z��������=�^,ҷFqq5D�j����{]��w��Q3�?ۚ��nh�T�n	���DrM �%��LXt������v\�E�u5V��� ��x�Т~���~����x����	jT����-��$v6��m��v�&���q�S:�}�\i%Ġ��ɓ��s4�w4�k� �n�%	}!�>ŀt:GqT��WEU������Jd7�� �/����� ��U�L��#iɀm���a��
�G�m�b��٠�4Y��pI���h�)�|���`��x�����ط$Xr����;�����h�w�{ƼX�(����*����s]��Q��x�HTck;�C��gغ�\Wn�S����,��������h�E�Z���x�K�7N���1`�ኪ�T��IG$�u�@������� ����������D�&�i�̒I�w�b�7�ŀ�/ 7��z;R�իV�®�.�`~�P�_w� 7_^�{��ܜ^���
1��(F�Ax�EqA�*�EC�8D(����`���*�,�*ꦮ� {�� �
u�_�n�ذkx�H6�gr!��]�)�ۈ�x6y�ǰ[Tv����&���z�G$vn�͝9k��5��=�X��_����@�}x ����I�'RI�{Ż����H���`���kw�DL�i�6�A%P�Q4�kx��ڳ�D)�ͻ�<����Fqq3Jh�W3V�?%3��x��x����7[ŀ|�Y��ɪQ��I&�z�4g��h��h�n�
�� IA!$!��U;M=r�m�I%�`ݰݰ�U�T=���2lA�uyn�L�=k�w� �7gyj����k�\OCۋ����Rq'�5���c�s��s�B +�h����O��ã-/:�N�JPodu����r\�]����۽��]b�L9kY�m�s�E�΋+�`��,���һ������ˬ�y�9��s�ZJ6(�7cve��\�Tٲ\���	�hM��
Uo��ޮ��0v��e��0�G�F���G$�:����n�}m�����\��L��;���Xt���%�䕀jޘ��]�k�4Ӎ�&h޶hU����M>�� ��� }�*��U�h��W55w����k�� սذ�w4޶h{��?�N!8`������?7���w��Kn�>��}r�v��T�ѹ����:K���:�/g]�YQ,^�M�Q�:��*���wI� 7d�\��[&,en�&��f��j�����w�
�J%$�T�)�e�V ���o�UM��M�h$�#�h]k�=N����� ��h��a45�UWe]�)�|�}ذ���<�נz�2�DɊc�$HRf��V M��}%`��	���R0eѱ8�2vp^ۊ���C���mM���7�NƷ]������'�Fr�|�o�Ϯ�N�X���/P>�� -��fL"�"iɠyu�@�:�h�w4�ٿ�H?u?O擘��nJ�7�ذkx�ߒ �/DD(�Z��t%e�"Q�F%HДW*�H�ٴ[ Eca@��������nC��_��=��[�,C������LX6K�5���j�1`�H��.*iU+T\լ ����~I�~�^���,��,�IәS=�Sr����.F���^YKb�3���j�͝�&K����s[]�K�k�Y&$�F�H"9'�r��=���� �����,#Ɔ�m㫲�� ���Y�
ɯ� {{� ��u��M�\�KV��.�Quk �݋ =�^���V�ŀE*W��/��n1�3@>��@��^���]�BQ����[�u�6����W55w�k�+ ս1`�b�l��N�v����Yt�0�����lt`�&�N���܌Y��zLm��p�[D\�3�f0�e�]׀���,zLX��}%`�vV-�A' F��h�w7������/��x׋ �Z��n.*iU+T[�X��x������q?b�:����{�e�q�o#A$�C����t}� ��� >���7i��t�����9��w4u�����rO/�}��Si�T%T*@0,�iBBJ<v��+F"B$.h�%"�͓��FP�[+V R�i\feѫ��Y��J$$A-�H�d!)�)i�M���ְ�� �H|s���a�K,	(V0� ���b��klё��@�ZIH�	��i*J4��	}�ĸj���X@�jK��U\XB0�AUv(��%�~��������   ,���t��z��v��S�6�-<[ȅo.i0  -� 	 �       �  �� �����q��k��z ӷjU�%@�0��"ݒ��j�ʼu*�W��8��9�@�N����	镪����+#�]����֚�W\�!�<��խ�=��b���o%��d�'�<.��[r8���7m�B��E��kƜ;�{((�qm��x�H[;��n���F1�nO&�nx�͈ݩ8q:w)��6��@pvQ;���hP8	�q��n'[n��3;�����ln^��ٰw-�6��s��:�l�`��"X��y��-�T=<�n�k����MYյ��>��$����l��������&����v�� Hԭ��6ۢ��#��Ѣ�[tͱ�M�6��ł{dM
�ܪ�Q���� �g���mӹ�g�@-����eL��e%��v��W`xU}+VҠ5X<Tk��q���:�j���Tp��HR�o+C�[������[x=Ð:	Q�R�Q�v 1� Tn�eu�+ 1�W�1��`%�7[Sj6M����ms� �^N��*�pzؒ�-�1�����%$�v�7F����g�nxꇣ�}�ؓ�8�&����n��t:o�ŭ�>I[v�s�{E�\�q���v�H���9ݻ���X{<�`��x�ە�)��˛��Z��MȹT�umt<�9C*;���&{r���4\q�쎛Z-ظw[�t�pU�'&.�Q�ui¹��SZ9�$ו��kd-�sI����e:孫<��/+��ܘ�n��ݭgs���ڬJܣ<ݞ��k6O)��ny_��cmu��&��� ʛ�.���M�,�_n�뭘nV���eYw`;[��>0`մ�֢7�v�6G�w=<���;W�uMմ�X����eNɫ�(������@}���߯��v߁|g�m�$[Z�+�U���f�m ��婝�iV��vĞuc=vx�U��Q��M</����ݬ��|�;x��)�'��3ӫnu���s��Ҍ���;v�n�"'�8n��<slv���n:�s���w<���x�n�Kv���m�@�c��I�Ψ�FpWk�wn��<mY1��َ{`ex<&�ힶ*H"���_�{��|��{��~qm���&y��Vy�����-��%�I�3r�����\N2�k��C�Eӡ#Tq7k�>z�`����n�/�5ov,�~g�~2)�j1�3@=�f���V�dŀoI�?��I�[#�7iZ���sSWx�������)�}ش����$r��q	�nG�yl���1`엀k�+ �\�1�D����ۙ�{���z٠yu�@�{�����WY&i�R4��cs�	λ\�� %��wK��3��N��1�������)�?�ly19� {�~��Z�/k��}!���.��Jj�Ԉ�ԳY�krO/�}��0�#�c!RI ��� �A$@�B,VDVI!!D$"BU�U<<��X�x��7y�D�ιeҩ*nj�' �zg_ۚu���������2�S##q�$XG3@�s@=�^�IX�� �Qn��%UM�M]� ����mwu|�}� �s@��¸�jllR&�l��8���aW�-ŵ�����ܻKz�;)�a�<ɵ�&dȓyNM���g��h��h޶h��ʮb!�7#�<��tD��v, ��^�m��-Sqn2��1I�9�u�����r~ �$��(@bE,�S�i�gV�_b�6V�s3qqDҥjjf�`tDDDϷ��������舖��X�]k���+���E���䕀j�1`�b��/ �W���q��.�⣗�x�c���6dݽ%;�l�X
�7Nr�s@��Uv-<�,���wXæ,�LX6K�5�+ ��SWV�������S7k �or�� ������׋ i��b���CmFӓ4�٠y[^��31.�_ۚ��nh}��D̙L��&��m��kŀn���$�aDE�
��%�&�x����2���� �tŀwI� &�x�%`�-}�9�ې�5�μ�3��Y�D����d�hu���k��AY��Q��'[�H�6�Z�~�� &�x�%`��X%��RR1<y14�� �u������Xt��iR�:�t�n�drM���x�s@�s@=�@�렙I90x9	#�=�����X�k��	(���{�W+�V�j6��#��w[��{��<��I<�{���6�� B,`��B4e�ZZJ���-%4 U�aJ���{o�kW32V]WY:I�� $�O��g���Kb� Y���v�����@�˻8�2��Oa�C]i�ྲྀ�k/h�9�M��ǝ";��j��e�����!d�ġ��˗8@��6�K�k`�;vd�{+ې\Z7
'�;:��+�17i�8����غ8�n7J�b��sí�}v:T�6�u'N�T��c��-qO��z���ۏ����.m�C]Rյk��Og�(��@y��,�wPZ�5NL���������s@�s@3א\���"I�4��<�u�{ƼX�x��k���B���S'��1E�q$4܏@�/����� ��f��mz�����C#Ndq�V��1`���䕀n�K;8����ɉ��h��hV׀n��1`�.d��H�.Ƨ^�q�\�\l�v+VD�5.�m�3���؞��7��"�drM���{���;������=z�&,S$m�&�˻���x�"�A�r�
 S
��	KHJF80�hZ��%	X$%Yc	v�d� B�Z6���#	!E���"T��DN(�����ŀw;�=-��=l�r9�j6��D�h��hݮ��3��Հn��X��ȝL�d�S"�4��4.���+��w[��א\��d�"4��<��@��1`�b�wK�7h:XU]&�Ӗ{yz�v�x�\����g�g��x�^��t����+C����i�ȴ��?���,�LX��x�%`����b$jB8�s4�w4��4+k�7zV,�\��ݠc�JӧUk =�� �[u���H�S	
Pm!)"��� �@h/�|�f�Jŀv�ŀv���T���n�.���(J}]�X��ŀ{u�h���>�	��b��Z앋 �� wt�mH�{��q�p��Ɩ��X�n9�v����M:z��756EN���Xɬ�y�n��R`&��X����ny(P����XQ����(dK2!�3@;���$N�X�V,��X���i�V��Pi�&��}V��Z�4�w4�����rW1�#�!�$Z�k���ŀ���
"!E(IGmwN�U���"�A��s4�w4���/��@��{���ⱸ,x�#�Y�
��x��ԝ��w7��ۑ�i�O\,�c"0�<���� ��4�j�=z�4�w4x�b�&��"��I�_;V��n�@��s@-�4���ƤNLQ,N(�Z�]��{��^�4�j�=l�r9�j&��RC@��s@/u��h��4p��T�2,X�DI&h�@�v��]f�{���R�#O�iV�I�� 	#e�n�<t)�s(��gRY�nC�WV��v�M\��p8u��z箺S\c\`9z�`�a���{WO]�ŷe��C�-�*�u&-�&4()s��O'm�q�0],�7jN���EO�ts5ۮ�!��m^�wc���63���<��4g�ݏ�o���V�񶵺�8h��s��m����pk-Ƭf�9��{��͟�;e�aU���Wmی�χgz�։�T�d7	\Ek�� ��z�H�d�3&��rx����m�0	�1`�/ =��n|�����G$Z��4�w4�٠_;V����Q�/�5�y��/u���f�|�Z��4b��C�4�LCnf�_[4�j�-�Y�^빠w�&+n5�E25$�@�v�I2�wLX6K�#�1U�5Β�2H`�1ӈ�&��»gx��v�C�n8ў�3��pq��)�m���]� ��h�ՠu���Lr�����]�x�e(����w�?Ss�6�Q��D)�Y\T���,�)�r]]� ���78m��w4Y՗#&d�F��nM�hI�`�ŀd� �M�q+���8�@��f�z�� ��h��@2�����)�$���6����Kۭ�,.�)��=ye�r�Y�e��q�3����"q��w4�٠^v��u��\���CNf�?7x�np����g(P�G�&/�&�XdS#RI4�����t74b��	4��9���M	P53)mi&��+,�2��J�B�Әa(FiD�@� 1� �CB(Ȓ�#���4��2*,����6����h� Jc�B�l"�^h�����)MM��{�f�=Xl����c$$c ��K�a�@�# �760
i� �AFHBdF$k�F$D�F��J�֖]��[Km���B�Ke�PM�h@�ڠ�H& �"*0�/�lP< *}t ��l>)�)�W�����%��RQ_oذu��=��)UUeF�,N(�Z��w4�٠^v����G H�M�2'�4����� {M� �ZŀrI�<������TYwny�wlW;Jqu۟6�θ6g��ipc�n؜tOj�c�F��;_^ ����Zŀ=o����d̄PPi�&�yڴ�^�s@/�� ��.J�H�)c�Kxދ�LX7���#�;����5�<Jd���� ��4��g�/���y`��#*�
��tMLլ ~n�����~�� ��s@�B�k�dq��<z�J��K��Ѷq��\z�nϗv�Y��x�n5�E25#�@�v��\��=m���f���76��D'R-�ZŜ�)�{� v��v��|�;�̙�n)�<��z۹��f��R<oE� �*S9b��:V����	�/ �;�ŀl��Yr2fB((6܏@�v��]X�x�>n��p����ݔ+[�[$�U�m&l��n';J<1�����j.����c�V�݅9��%��P=��v��]X�;��S<�AƇ�tl�����-�!�˜7X0�j�e�[:��Y�vØ̐[(e�3�C���=`۩vy����Bm{g���rf���݋D�$9{Yն{p�N��S��dVJۿ۬�3��3���7cZ���+l�5�S�vF���w�uo�c�k]7�j�����{O �F��c����O(.�q�[<�U�E�x���c�G�������`$ŀG�V�R<����w_D�'��4[w4
�k�;��@�����eX�Rt��Mլ=���ՠ^빠z۹�{�D'PڋE28�@;�����^���sqco� �9�I4�1`$ŀG�V wIx]�q
�dL�(��`��uY��R�ԛn��I��n9�Nrl���礇��멁b�7|�x�������(��7ذeuL�9X�T��ssWk ��Ȅ�`Q�E�z����X�x�J�C������rM �h��i�1.�݋ ;{� =�2�ZWr���Uwwx<�|�ov, ~n���x�A)rG�D�%&h^��}�h{��/��hP���,y��(���r�s���g�hz.�$e1A�4,�9��@�$�D8`c��1$���uz��x�x��s�X�RK:J��R�m]M�]��]�D$�L��b�=ϱ`|�g(��'��b�UJ��K%MZ�����X�^,"�QJaD%)$�kֽ ��f�޳��"R
8����D��|��� �k��������:��I�!�b�2&���U�^�o�� ���׋ ����R��.PybRwV�4rƜt�LZ���"�G"u�J;��N�Ru�ŕi��g�� ~׋ ���С(�C�_V {�U/�̆�,nI&�{���빠U�^�w������cD���X�LX{%`oK�'tŀjw8�p�ǉ���s4
�k��Y�=׋a�O�^,S�%�UIb��dq��w���]���s@/����e�/��Ǆ�8�
�FX��-���L����:�+��]9�:�t���W�H���I�^빠}z�hzנ�@�Y��r)S�h^���J�ޗ�N� �*SlQX����t��`앀�/ ���빠rά��3 �nG��w�?kŀ|�����%=Z��ܥT��aB��h�w4�]� ��4��h�q�"Y̄t�5U+�U����R���9s�3n4�KEu�eYRzu�چ�u���W,����.�kkn����͢�r릴�t��۵���`'u�N�E�[v��� G�� (�N�L���S���N+�g&	u=Gk���LDog��ŵs�{`)5\��m�^�6�:��B#��J-����'�ϕv�9���v�;"W���w{�ݚ��$�C4ɝ���7���7����5=&��[*��X^���We�<����扒�<��4����Y�]� ���2��;�M�Uk &�� ��xޘ�N��]L|EEY��)�����4׮�_u�޷76�c��� I&�}�V�� M�x����j���v)S"s4��h�Y���ޘ�w��	�۪�e�MU���H֐5���X�ra�g�b�y�4�^�d��C"ĉ��ɚ}�h�f�}�s@��s@�YcJfA�(4ܓ@7[��Z��
�BP�:���=�w4�٠�%P��?� ,nI&�;�,d���J��/ �܆��cDsL�=m��*��@;���\��?�I�I��#�+ ;��t���b�5ht�|��캱Ӯl�lG9��F1k��C��s%���[�6mVc�\��IMx�%�I� �&//0$�`l雋y1�Ac�$�@����s@;���l�;��q��8�%"�<�ŀ�."!�	$$%
��Rc�DG ��]���m"�E�#��X ޻��� o^,�(�����`Yߙ�5��($ۓ@;���1`$ŀt��:@ut�R/�j�ՠ����v��1+��C���h^z���rm(ӑ�I�H`���$�-빠zI� $�x�%�����nϩ��ǑI��w4޳@/[4z�h�s�� �y"��Nf�[�hi�â""g��,�v,�>��őL�I$�/;V�o]�����*E_HZ�{�$����L���(<rdR-޻��w4޳@��Z��+�I#���k[q�v�ͳ���\)�z�;A��nB̺��q<�3$��)�I��w4޳@��Z�w4sU���Y$H5��t�uH�	:b�'I� �[(��g�Ƞ�nM�h���/[���4���*����rE�6�,�x�����Jy�t�m��!�D9�"�4��h���78m��5JQ	M�"�HA-`ӌ2P����m4��V��ٹ�,!,ԥ�D!F! �$ BP�b���`!@�$�$H�
B�G0 GD5!�P����H�"����F�)f��d���(���
�0%��a�R)D K棅$&&���P0�"Pc`�Y�ZB����!H�r�� R RV�q�L��IB6�X�1$`A"� �"�#��$(K
���JQ�c� ��,ɢXԕ���(@$�#���I&�HAXB0�I0�Ks$H�#F1 ���HbA� H$B0i�D##�t��u��'���? [Am   Z���vۤ�z'I�N��9	��-�n�ݻ����  � �       m�  �`    ��;j\�k�Ct����Ӭ���'^�� Yi��dڶ�`�P)j\ss*���l�(m
)KU��B.%Z�9�cl�=�7#�a������4u�N+c�W�蹋;�9�8w�Y�TǺ�Gm�л��,�.D��<j��͝��P�t�%yn#nr�gn�2ش�{r��`cc�LP�#��ϻn�]�ꚻI�ҶWn4�F�[q�G;�;�wm���+ �>���2灖�\�q#�<4�cn-�[Q۔4z�;{�KJ#�U�A��Ȝ$e����[�T�ع����ɷ"���j���g�e�ܕ�Z�W�۳�r��Îڭp��$&1�������<:-����vLνR��Nʴ���V�qڞ�S l�l�Tl
�UһcT���|�-��mä6劵���p qmU�<��+U� �u�F�����`ձ�GX��[l7B�oK�K��Ҽ�yhC�U�SUR��%w\�U]J��Ofx��B���mP�䭸 �x\[��3M�@��h���Wyg��nWf6�X����=�q:�o[?�s�͸m��{v�(�-%.��s̾N��4l�qǃҶlۭ�B1�#8-�ikX��؇v���s;�����'��/���t��ۃm?5q��|�tx y)l�� ��ƚ8s�F4+z�;�ua�k�ؑq����͵���N�ɺ����k{�e^v�w��׷mZ���;Pa�̦y�����wF'[���wVjM��Y�S���o7i�[�����t;��c^�]�ŝ͋)�RM�)s����z'X���s��"/c����6�/v�� \���-)W.�WT��S-Ug���;&�	WP�r�tD���e�%;���|�fPz��y/kexܘ��pf��N!�ĖVMk5s!�h����D 6��S�Q��x��_Q�A�߭�u�d�L�M]i��%ܶ����ӷH�s�X��`�-d�Y3��˷a�1�6lq�]v^78�o6�s�A��~������8g�6��ۍ��^;3g�q��q�YF�����qlqdՇ��;v�d���4��xN�=4��v˼ɒ�(�X�윗Ba�@�g��R�m�!�i;r�q�:�3Z6�a�[v��8x�����I�v����aV�ˣ5q>z��8M�s&f�3��EŖ�c��D�sd��
�y�#���Nh����c&<CD�0��'3@;�~���I� �&,��o��+s#R94�ՠ[n�z�� �٠{��,m�a92)�m���w4�f�yڴ�0�� ��bRf�z�� �٠^v��w4sU4Ta����� �٠~\�~�� ��X�֊�d��\��Z7���/m��gqv�b�
�l�p�v��3�C�z��u%��'E�j����~��o ��\�!G�wu��I~q`��c�H�m��/[���x������Ⱥw�[V*v�Zj���5�b�ۼӭ� �x�[�Tl����	9�m�@��^�$���1`O[|F���V�];�M˭z��h�w4�f�W���߫����[J\�,\���6.ۨ]�{y��W]���٪m��lt�;E�j(��-�s@�[���4.���aqI�	�GĤ��n�[m��n��Ŝ�%
d}S�Rt��,������X��x�[�)|�"#!#�BI�JA�,H �A����+�%�$���Jܓذl��5����ȃXH�nI�yu�@����n�[l�{4����nG�6�,���������N�X �n�v��e�ݠ����t+ۭ��:T<ő�˛����¥��]s��+����vV���&, �K�5���I&,�����0��'3@-�h]e`I� ޓ����h*�Qn�jG&��ֽ�w4u��m�@�렱G��(<�Gz��h�ٹ$������ă�-PҢ�?��2f(�נ[f� ��LjZ�7�ŀIx���	$ŀN���g`9��"c�;��ۈ��[�g��Ng\2jB&�7lN:�6��$���X$��k�+ �LX���,�eQL�XH�nI�yu�@���zLX$����7.���Z�UwXm��=��á(��N���6{�=�݂%ȿ�8�0Ȝ���� �K�5�+ �LX�\Fe�(V�F��� �٠y[^�m��u����9��#X�P2G� �$����yj�Uɰ]�A�1כn��c80rWm�F�;Uػ���/;���\�l��l�����]�˶��+ڹP0[�N��lvĀ��:��:���u�j�^����n���-�X���#{t��m�ݺ��3�Q"8�8���yR63�P^�������{�vG&�O$n���O��N�3��6�Ec��m��3�0�'5��K=y�=r�'�#�Fڃ��b�An�-������A�O=E5������o��/СG�wu���X��DPy$�H�m�������� ;�� ��� ~v���EY7e�nL�;���m����۹�z�SEA������4*�`���(R�w� ���:nm+��E���]��m�В����_ �v�[l�;���4PlRbO�?����GB&'��m��C��=.���l��*rE�xR���*������, v٠y[^����Ȳ8��"s7$�߾ٸ(����D�$�}��kp#ޕ�I&,Wq� �ZvLsV��� ����
&{��`�b�>��T��4<�H��<��@������ �٠wu�X���K$���m��u��m�@��pK�4��⃌�LO�)��iհzi$�5j�l����On|r;������ug!&7&h��h�����m��=Z����F�ڎL�m��%`I� ����.ݥt�w35Ww�z[u�6�,�U	HB AE� H�>I>�1`�/ 7S�%[��wi�i��m��u��m�@�W�<.R�WE�+���n�� �I(��������`�y��1�c�0���g)�4�K��g:���֮��U�P1˓V�ѵ� ����x�[���`��`)=:����$C��M�����h��h�f�{���Dm�c�8��'tŀwI� &�x�%`e�����i\ݗd����o���׀k�V�$��WLXJqӍ��.�2G�4�٠y[^�{���n���¸�jllN&	��&�2@�䧠4��h�hnz|Y-�ڗ��wU��s�����F�rM����w4�w4�٠�*��"�$B�ۑ���h�b�	�^�IX.�d��V��`����� ��hVנ^빠vw g�A24�s4�٠y[^�{���n��r�bx�N$$R94+k�/��h��h���<�""=7��ݕr�l]M�r�J�Z��veؖ�F����h��6�N�V�Y�="�D�n�[��sF�b�ѥ�:+��h�.�<��ZOc9��[d+v���5ͷ(��93�t�v��X��D��-���nl ]��s�Y�6�����k��nq����`S����#m�n���r��$Z�{z:���^�z�l�������t�v�b���1���{��{���]N<�s��2�!�]S�ђ�ԧk��bm�`L�t��i��νi#'�$q��?u���w[���f��mz��T9I�Rɚu�� ���Kn���g�J&G�=5<ĤQ�8ܙ����y[^�{���n��A�+3�4��h䕀N� � M����8��P�$B�ۑ����;��������Ͻ��c�b�Hn2$����vM���q��G���b�Ät&tR���<�r�Uw2���W@��^��X�v�w���s@��� fA"di$�hm���`�� �o��\�O�ā�G&��mz��h��h���\�X�9�7�%����J)���`��`m���^�}fF��)	���n�I%��J�$� n��Bq���	�K�l��2�s�����θ�H,��y�d���S:�k�m�߿e��J�$��&,Ɇ�(�F1<$i9$�<�נ^�s@�[�������#��H�#rG�^o�oʑ@b���J�"H��Q� �ȶB0`�"X�Y1M*{@Ɣ�p�ĕ��Jer�� H f.���d�$��B��,@O=�B!$0�
�|ˆ�B4���`KHJ�C7�x��n�n�{[�ֵ�VP�; F*ԃH!c@����9�Qe%މ�k5���!ʄ�H�4.�Z��Q����"�D !�A��R����ty���)$a�H��y20��	�Ł!�pdt�!�hdP�sIJIi�����Q�+s��,��̬��!!ZXA�aAAOPS�\�D���� |�_Pt���O,�>�h�נ{;���K2bR��oI� 'Ix���	�b�5w���)�$������Z����7�ŀr��C�Ε:�]7hn�z4��]c:����zt�[M����n,���#�)<N$$QI4.�����=��h�f�{�n,M�4Ȗ9#R=t���1`�/ ��V�ֈ�#hy��rf��s@/[4.�����=Z�օ�"G�0�w�zu���� �Q�$��"`	,HH?(i *�BN��X����)P��E�L������ z�,��, z��	G��p:�6T<�uí�'g���;J�L�<��`k�8&P]����\�M�[�������݋ ��� �}	B_Hl���56v�h�����X��X6K�5���N�~M��?3.���ڹ���XϺ�N�X�x�u��s9�Ӄ��RM˭�wLX���l��N�4ꋶ�D������h�w4�٠zu��"!D|骧wsU4�	�u7".���6�`�	��ݘ<��7Q ���]���Yx%�t;�:�r����7=��غ�:�m���B�z�s�[c<ӡKvݲ�7dH�x�T���Վ�:*�ClrYv����>&:9�{p׆.ү�9��nl�cK���N�nN�N枛=mGn��Q�ѷV�������Ew=r�ӹ{��r���JI΍��M�<D7����2p���!���r�^�WY����9��X��}�ny���f��Ej�v�_v, ~n�N�X��`t��D�q�H�rf�^�h]k�'I� �� �a�J)P�t��n��@�u�@�n��빠����j�s@b#rG�^�s@�u��	$�Ϥ��pژ}h��[�X�LX$��y���I&, _{>���e�5�ڥiW���]�:s�6�F3�BՌ�9՚,�����ɫ��㋠�����xӭ� ۶~��/�5�ۚ�T?э�D���M�ֽ�����b �DP�U	D�6��x��� �뛋d���c�5#�-�s@�u��m�˭z��T9CȤ$�4w]� �٠|���-�s@��WR#����I�m�@�wJ�$��� ��t uHO�{W����Sp�ٞ�v˳n�s�+FQ�e��ۡ�'�	21�1��#I�&���@��X��, �K��T⻱�h������-�s@���h����^�˸mLAb�UZ����� $n��B$D �����AF0!�F0��H# �!���Qs���7��`gZ�q���L�$�� �٠|�]`���%>o�X���U4����E#�@�wW�[�s@���h�f��� ��,��1Ą�Q(!aB.,㍮u6Bv���jǶ��uɟa+[���8y���c�4��-빠}�w4޳@�wW�_Y�C��<�� ܙ�}�ugB��C���K}Xm��Jd�T��!uU�����`wu�N��w4���� ��ǌ�m�m&�Ӻ� m�XۯP�$A�d!!�"� �� Xł(����������+Dͩ.�q�۹�}�w4�f���@;�n�v��e�]�fkUQ׎���P&��'+�a��.��n�u�&m��l�g�:��{�b�	$�ϺV$������1�dI&�h����^�m����s@�3��mI�!��R94�uz��hu��m�@�ֱJ�Uw3E̪������Q=��-���� �l�<���/�aP�M��9Mɚ�n�^�h]�����_r[dI��,R M� F�M�Gn�r�4Y�	Qm���ݷ`~0�Hq�S���;�N���n�[�*<��pg&۶�x��Ƃ]�3��i8�
rR��G�6z�&�%�N���T�a����[��/Y�awֹ�{o\&�m�Ƹ��[�d��Mǭs��z�l1���7a����δO
�u�1���ͮ���Q�[�n+�;�����|�?>v�;��unt<���w�n#��z�g���Oh�U�:L�|��A�4m>�uwuWk ;{� ���=��`kx�b��3�6���h]��t���%�w"��E
�nc#qǠ{��hu���[4.�X��2�ȱXUZ%T�Z��	(�>� y�^��u�{u��>ZܙSj��2$�s4�h]���n��![m�7���G��v:�=GW$�n����nl�790�oi�)�!�H��h���=�w4��� ����K��#L�c�D��=��a
�##Q��� 7�� ���/�aPأk$r8ԓ4��� ����uz����h��G�72A��U���I%3��x�}X�m��n��Aݗ�&�6��M˺�����<��`���\�KB�l���������s��6���ʌ��a�N:����p�9"�.����q�������_� �I� =�^ ot�WpڋBs�9�s@>�f�{��{�,�tFS�_X�]�n�`���nI<�ߵ����({���0Vn��[��^u%dq9�"	H��� ot�{�,�&, �Ixޗ�2F��"�ɠ{��hu���[4��h/�cx6��gGOK\�f7Yhnx�,���m1�]�b��8ΜNr<��ؒ��9jI��n�}�� �u�����h� ��nd��mɚ�[4��h�n��Aݕ����NI4��ht���%�w"��E
��-������ {��j!}m\��s0!��:*a�VH��H!Ib�22FH�fGY�kL���h%�!Du�J�D"��E|��^�֦SY
�J�D�uV�t���%��K�7�b�7���k�s�l�D�;7��4�{]��$�9*N�uq\���֧j;i'n�=s�V��%��K�7�b�=�b�/:$�qI�d�5$�wY������2n�ŀy�b����%
�7��'d�2%�E�@4��� ��� �u��L*4)�#�Ƥ��}������n����}��=�'*�niIV�U]�U�����3�DV����V{ۋ �
$�"#��B����1U��U��
��" *����QU�������$ *
��"�
�X
�B
�
�T��H��*`�AA
�D��A �ATb*T`�EP��
�A �@B
�A��AH*D��@B
�D�� **�� �@H
�Q`�DE��EA��V�
�E
�Q`�E�� �EF�`�EH
�P��`*@��DB
�@`* "*T��
�*��AR"�B
� `*A��A"�*@ *@ * `*Tb�DD��D��D��D ��"�X
�P
�
�@b*T�� 
�D`*��@�
�`*E��@@��AD��A *@��@A�
�@ * "���DT *U`*Tb*`*@`*`* b* �� * *A"*D`*",TR"�A��@ `*@
�B(����"�P *
�� ��DQ��D�"���EV ��
����
��� *�D@Uh���U�dDW�_�D@U�U��DW�" *�" *������)��������l�8(���0�'�P 	
� R����@(%KZ"P�T��*T�  )�T   �)U�T@��@� P  �@�$ �JT�����R(QH �  B�
UAp    a 
R�@��@��$��uNC^��� /gt����jFZ)��1�Pҙ>����O@<2�NN]�� ��x�rk�N@'��n :\Q��wC�Ȭ���A���"���(��   ���à$��7\�C\_]{������g{a���B� ��a�b����K� �E����Y{�@t�f����=�X6�s����� h�۽����Z���`<�P@ �� ( ��� �����.�˽=��@�e((`}D�)�`R�N����gG��o�R� =1Ҕ�=�)�q4� N{= zx��(��: �)�N6PR��t��i��� � �J��)�ҁAf��  g� )A@P 
] ��LMM)� Ҙ��Y��>���<}[���nX�X��� �L���|
�ϰ|�4.�N�e���`2� z`"zG�2���:� $�  �
�������|����}� ���a�t�,\@  'A�Jb;� A�ϼ�P�@��8�siɓ��t��4��uq���2}��   =F�l��   �	$�M 24 D��T�   "{JSi(� 4 ES�Д�U*� 2 AG�IQB�#f�%����_��G�]c�Ұ��q�X��JJ"��_��@]��"�� W�` 
����*�O����(�5)�F	� B������)��Sg5�k�O��ީ��F����F�9O=�Ge�
,
�E����Ʀ�b`ApM@b	C��U��m�e�|�w�{�9C�z�c��U�Ƚ~��4�3\���udzzn���(e�+��3/׹ÿWvOK����
��tw���s>I���,��M��U��[�gЮu�{;I�f�oKѺ���j�L�e�y�4�߆j�L���y���B��>���g�'
�w^�^a�}u��m:<kP�w6���2�蘣���a`�)Yu2�M�#c:�W��ǽn�����5ʛ=hr�z*ӽ�PV�)�y�=��v�T���r�ơ��"�fVM��gB�^j�'�j��&�t��o/����f��2[.�7�V,"��1o&�XiWޖZhhR��B%D�P������ӣ���'�M4��,6�η�}sju7�/�]���U�u�9�G;P5
�a�O\����C�+ո���z��8ɻg�s�.�``���@`�0J#�Z�Ԧ�y�>z���ө�Vxt�rՅO6l��S�a�,��ȡ���B]|
l���Ŭ
$��`B����#���ey����q~������<`�4���p捲��y9u��������k�ѷ�	.�q+�T�bQ���CB�M��E4��D�0�n��
,-Ǎo�"��}�Gy��rjo
�u��b��D�Q��Y��WO)�h�f�̀2\˨t�/��ES�;r�#2�9i��з%t��$53��z�_�LeY�R����yV�Y�G�(��;�
�9�Z��5����=~�2Qx^[��U��q�"Qc+������e͹��:�P����j���D�Čd��7�SI
�*B��1��դ�`ez�ə2�=��n��E�[f~F��0`X&4�V�����i�|���°��Afh�ԭ	�)YV`�4�H�HSI��:^���GA�b�Lv���F΄hv�[:CC�!cC��
.����x}��O����ݿ;��u���0N*c�0"�j�x��:�>�T�>�Ǹ���|��8WdC<x�|Rm0�~��C����������WV�e!�/']f�~����X��U�Lk�8!�44�k
�<�%!)41�D���;m.�B$w� � �GJhRRP"Xǰ�;��EY�g���Xl�k8dU�bf���i��U�F��O.S���#RPЄ�4�
��T�V��=(��*�Y�W�������B�g�n��h�&�*�i���/WzU�3(е�a��ý;�J��\Q��,u6d�5�Ƙ��ǯ��3���ҴMQf�z=�"m��71�Zuk��J��N��I����⭊UӼ5��x{-Q�F�&!�!���Ӛ9-�H�wG;�aǽRVGJJ��Q�e4�Y�T԰ �D���K?~�`«� 0a@� �ԍ�0��$��@�B�$X�15h���O_�Kѻ�r��ўh���ү�N�+���\��������8�ΣȨ�Vn8�[ZV=��::��ոh�(����d1��L�ll����I˕�ɚ/fe����k���y�^���cM�w��Ҋ43u�᤺��1�����	Orz�|'*� ���2s	��F�9݌v�$Hy��C�9	!>�(qF���C,1Ց9�lW0�u��w�wÄ�:�ŭ�Y7x�!FVSȻ]}u@�Ϋғ���������K�XZ��!�T���;A�]�[�ʰڍT�|��SF�ZV��B��,���H0p�Z,���	cn�V������	���}��O�@�#4���EM�hܿ������p�Ֆ�WFai�XSI��I12*�3�m7�|�ϔ֒6CF��$6�-:�Ȅ��b�T�g/#�4�8)�!}�T�j���|���hm�3Z��,A����mk�橰�d@���<�h�f�orF�J)� ��ºٳ�MlH�&�h�t�G�@�;�)�m5�����t� ���J<dV�k-X�8�ȓe;�z�cmA��Cl^Zhq��B������;)"�i�5�ύ�55�`iF1b=�B���I)RIR�
CW�7�#b���4Y�X�S��{��ђ���]$M�{"l��K���N��jd���+JЂW�����ǧy���
H���!��u<�6�B?
�z5�'��@�u�&�	�gaWB����."�����]��`0,�B��DN�	��+��!��U�1c�g����������{/���U��5٦�����)�����u����A,�L�=\&Ju�W�_�OC���c���>Xҕ��ݞss=�,��I����A��]�-:G�@�4k�����6G��A6r�/{���q��/�%�P ��Z�x�esm�Ma6ٚ���:�ƥ]�93Һ�Odh����|g�0���2Q�ͭ�S�rq�ǃͮ���Jf��9�6����O�^{�u�	�(<a�q��vU�[�f��42�E�ifl>���&�H8	 �U`0�H%bH`(���.�pzTc�M�C%��~��ny���d�kA���`��ǒkU�3r�ǁ��+&�
/=�껬-x�b`��J�,�a�3�a�o;�Ŝ|����_�c���'m}۽(��|p2+���_�p�����{+G��RM���b� +�GI�74_���:�H*Vw�>��l<&Hi��۟Nf������P�E��Wc�v�>=�~��S�H�7y�V���%]���ˮ��a�`X0�b�]^6�Vr���������CQ��C
.�Ɠ �"i'x���%̦F��&NzVy�y���2S�m�� �»�W�5�'v�}=<�X������	��V9��)8���F֕@��e��_�5e����YHe�_����{���p� �B!zk]vGGő||P���QI$WI��F�c�"!Sd�G�饜D9-���˷8けU�a���@�QV��c�~UH�z�y��q���x�5�hPd,m�	G�"1�RH-bЉA;xv�ߺ�ӉN�o)�]nw�G��T]�*c����u���P�=�2Y��ި`�R�4J3j�!ǏX�nX,�k�nR�I��V{�3����eg�d�u��@�����A�3g_��S�2���͊�x�A%m��γ�*�L�7������u�S)#y>�`� >I ���>)eW�x�:r�JldT�'�u����M����}^ή��C�.e!��>�ꞯyt�py}��yמUC���U����u�y���Ǆ�����2E���8cb�����0�ƫtN��Q�����N�s+�ha�V��^��8s����@�.����
h6���<	 U �S�0��"�ԣ 逵���!�X��ϩ��1B.Ͼ�s�1�0<ؠ!����a�����!!~�a H�Q)"R!G@J��B�CR'�<xHU���փ��4ݧ�$<�������T�m_�F��2!SN�|VWFÂƚ�ǟe�9����U���.�Y�s��Vx��
,4��f���D(-a�OB���ﺟ�Y�a��(m@d!Ef=����ː�*�e�}�x���WnQ<c��+IM�x���&��(�Ƨt����2����4�"�=�v���a8�Z�k�
/,˨c/����k��=Ŷt,y���rT}ƣ�bW�ֵRa�쾂��!�5���fa�@���QI�i�73j�����{���A��/r���k}�+!WW�Ӷ�s{Oi�Ϋ3����v�~>�ì4�%+�Ϻ��<4���������^i�ߣ�ʗ+f����>k�"�H��
����V[��b�!*����o����C�2"��.�:]Uz� m�Z�  8,��[�d����M��y�!�n6'�*=[ ��
�˥�� �f��5�P�!Cn5�4���m�	Жkp6ؑ�� �n�ie	 � [M��H�8�^^����  � $�m�4��84V�Y�`$m�[Cv��5I)��       ��     �    	           �           ��            -�  p        �� �    ��                              �        $���g3�@�#��Tb���0�@��*Ҷ���٭�^Z��ˢ:Ltڮ���Ut����YVU�^��kk�mz�$�v���mr�D�a��o��vط�/3d8[xI��$��m��k�m�H @:�8v��۠*���5 �m�h[L� H	�F�v�ہĔ�Uݺ�8-P[@,� � �:� ��Bs�tiP� Ԑl-�';$�ʺ˱�#jG�ֶ�8����v�)0�ڇ��9�EAݢ@�S��p����M� �eB�z�[��@yW�^�`F�s\/_��:6�����iPk[)l�L^� t�-��f�ڳ֝���k��ڕ����OW�l]�CX�͔k�X(+��Ūe`;�cYNB�@����ʛ Il��p[R�	(F�j�Z�U����	���/_�u��v��$dYbl+���n�z�92�-̎�Ye�ͮ�"AsjDc��j�56���l=�j��hV��۷}��}.ַi�T�Z���嫳`�ӡy�ȆW��MU��쪸���	t��<��ԨY씣;p��L�p$8��n�,'6���'�U*�UT�����;���w��t%��M͝�Ɯ^9]���z�%�Y�I��^�A5t�U&�V7U�WVVX��<p�k��V��Dc:oLu��å,�ˑ4m���\���*p5����m�K���3�mu�$*v��^�j��Gr��ə�oM� 9-r۳�3^�Ö��m�jݸ u��WR���Z  n�\�d)��l�h�6��n��B�@UUK�s=:�T j�����@Ue��@kiX"6�u\ ��vj���Z^`v�� l�8  p ��uv�2"F��v�I���  H[%�;�[@����$�:��Y˻:n� �۶� HM:v)��j�:��i��k(� r�.�[@��`� �@ � ����8�ɶv�3#�m���@�6�	 6ضJrI?��*�	��6�-P ��  v� ]6 m� ��[N �e�	mvN[%l H�>  ���#m�   �]m�I Ʋlm[�Ԁ��-�ɀ ړj݀�H[@m  �`p -ɤ�km�  [M�m  $  �   �I�6�  d��PÍ�   ��-�Uo��  E5�  pymBk� m�����    ��`�l &��mZc7Y��-��`-� �   -�;v�m��� 9�u��`-�� 6� 8�۶����Jݶ� �K�ņ �   � 6�[%� ���   p �  n�[pH    K��m׭����H�M��F�dݺ�kp��A�`ݶmmfn�&�m&�6�6٪��Z $lq��'6u�� lݮ$���;m��}������  �`Z�a䮞���&�i` 6ؐ�`��6�m���0 �[{  6݀-H�m�����C��Ӧ��mE���mYo7�k�t��k$p��[x$���V�.���ܓu�Q��3���\(�d��Ƅ4@�j��a8i�qN������J���VYv6�uU,�G.�SWl�]��4rR�+�R���<役��l����zq�=H�x죰<p`np����ge�[յT��9�m�8h�q�z2'(b]�d'$l-�%���[[cd_�����h�ʻ����=4�uɤ���m�M�o�k~����Z��&ڪ��r�;r��!V�b��;c��_��}���WUU7n��p���^��^EE��%�m�M*�WVՔc���q��J뭮�9�[į5�ܻ�3��d��]]mi�����\!p���ڒ0�� ��Rp5P]�aZ*�
�����wP�m��L����������n�$�l�$��N,�糸n-�q����6�咚J�����e�lr��	6ȧ	/Y����K�c�_5J�ݺ���jAi���Z�]0�M�̀H�h�rU[uUmR� �e�� -6 ��-��e�p-�Z�N��l-�m��m&���Z����s׶ͺ�^��@ ����@H� �C��6���[@ ���m��� ���� L�[.�c?D�[��0A��,�9�Hi�];am�r8�//-*�UUJ�G �ŵ�ӄ���H  ���L`Şv���)�cs#��i_��|� }UV�Jq�UF��ւ���mϻ햒�ê�Iv�H��G�k5�i�U/\v�P���ْC��nm�I��@[2����q��mհ�E'-�姶�q�1�m�l�J����7� n�(c���#4մiz��ۍ<�!�x'���^vk�vŴ;#/�I'6�M��8Ŵ��Ѻ�@�m�l��k��   n�˗� 6�]���D�c�-�A��h�k�h���/�Mm�l��@[Bln� C����Ȫ[d+�ѳ[:kMSO5sw;��)V��겳0h���K:��m^�����ONؒt��m�Hv�k5jۖ�@��\m�ݰ�$�\�VpXcI��n�{B��1�JK$�dZ��c);-.����R�+%TۑZ��j܌�I:3Q��6�܁�RZ�֞�R�Vҫa�R�[��o�ұ�����M���
ƥ��.&��-ڪ��I���@Nں�UQ�*��*Cn����D��� ,kv�i��pq�i�J�YYî������  $ +j8�j��\⋕����;���[kK.$ m%lhhٶ��]�]�Uڲn��I������NKX�;S����\G��{f�-]��WiW���Jm��N��B�AN��튃����]��l8ګ�Y�c�BTkn!�/2�5ml�݆�񑠮ej��p���͜���u���$�6nؑ�3��*0UM�h��@]X�T�@VV%�,��+�U�¹�yn���;$J�Ol R�<�Us���cs*�\��Z��Z��(�!�ZE�@m�  -�� ��� �H �,�-+v[B@p  �s���Y�0(-��%�ڭ� �6��  ��   �(m��.�֭���[@ �Hkl� ���-��	m�ڢJ m����U]*�J�V� 	��� 8m�-��h    3����@UUR��Rj�`   p[g@ò@ ��m�iv�HI �  �F�|����  ����m��  H	;l݀ ���kkm�  , H     �h���ie��'�k�����s���mm-�8 8l@6��݋h-���o i�@ hl���v�8$�d�����l�Nf�j��%%�iM`%UU���8��vv�W�]� -�ٶ��f@����m���h� ��:�f ���  l۶��kn��  ��.鴀$ Em�:�� M� HpڶH�kh۶n�k��#��6�b@6�`  �    *�J:P�U(ګ����KS���Cm�3.�-mu�b�tۘ ��bմI��Q�m$�1�j�r��Rݲ-F�����.�U����������f��]g/m��k$�Ͷ-�S/
����8�+uUT�#�x�����;,iۃ���}Pv)�[���ju�����r�%����� ���΍���q��#��A"t��pYd�칅Փj��V�yq��v|p+�La�^���AK���t�9i��ٚ�)k�t�R��f�� 4\.�7(H ��s�ju�;mm�f�d�^��ۋl�   8	l�޸���﯏^��5�U�@R�6�@ n�u������� 4�� R��\��v�MV�]G)�ݰ��,�)i2q� ���]d��yiy9�:���]5햜��*����5c
�ԫJ�Jj��nn��N�k�$!����i,�7R�˵㬮��e͹�Ԯ��������jOsl�v6�W��JTG6�I:R���O���E��7��PT�"���(<P8�� �!���l � �@O������	�P�����N �T��(q�+�A]!E6�M��p!"��#!BH"���#	$a`��� @�@�Y	 �#,���D��!�B0�E#��"HH@�H� @$�F���$"�"I�$D!$B0	FX���`�D��B� A�$`�	`�HA`X	�	�0H�HH! @) �HF�E�$  �FE4�DA��+�E����	
F,#��b'�U<*�T��tT�|�a##$�1 �H��B��$bā "��F!���HB	 D*���`'��"|QZ(�@8�@Ҡ�#� �
�|"Q��  ���(i
 qF�'����� (�u�
�$V @�B U"�"}R��18�A�PMQЁ�
����v� 6.��=�>Q"��iD�A��a`hP~��P(�P�}Ca�~�+�G��<�y4 �Q�� `��PG�:*5E
)���`D:*�Ut�yA�1jA_�SK�ҭ�6*�@O��������}A**z�{�]�Yw��l�ً�v+�38z��s�r�m�K�����H�(�&ƪ�8m� p �� � ��I      6� ��BFA��c��MKn[b�ϗ-��Tv9�wjH @$�	�Xh�_4��kc�W��-�.m��qb�]r��m�]�g �į/g��Tr��)�]v;r����ۛ��0��v���>L��9u&m�nv��5�R'Q�ˊ�;γ�(<�q��f����u�j�n0���Mv�0b<(�y�X�skT�3vXT3A뵓���s�9�V��ru��$鳁r�],UB�F2�X۱��M���[u/0V;;I��!�p:��H][����m�Z���L@��-��V{f�¨
�n�$��wVm�:�W�����<dn����hr�P�Q���r�jkbx�`� �iܼp$n���u��9.��H�����G����0`*���<\��Aۭ��/pf�<'Z	ɜ�K�Վ���q�e��=�΀���4ȸ;�u>q�nq�;t���4[W'm�.��Y�H�)D��Dgav�O<��n2�fÅN�s��*�R2�:��s���i�n}���ݨ*����n8)��	d�v����=e�Өa!�Dk]v�	6A�ݵO�\(��0W��+�;�wv0pg{�@��8��n ��m�4Y�l�2�a}i�,��CktlO]�y�W&���:dE���
<+�s����f��0�.wg���v]�jUU����VW���6�*��z�*��]`��]��=3��ʴ��-S'9ڤ���Ĭ�F�U��2�4�ZK�;Fkݶ�V۩��</=�gNɩ�rg�n-���&\�Aqڕw���%��Uu%�>#���ۋ�8U�֮ѨۊC/k�l��h�^;-qs�g�t�9�=�)^�kY�<o*�.�]R�K��I�ԍ%��K/Aq��<3��V��8�޵��Y�u-��wZ�A(�* �<�DO� hp^!�PGJ(h(�kd�����Kw�K���R� �A\�{.���l�P�Z'4�ύ��)�d�#��;&���B�i��;�`���W��oE�2с�����::��w3ѹ3�5�Bp��;\�W�Q�p��j��'V�k^^È����ɹ�����6�+���x:�,�
4�#@�:��5]�mO0ی�<
��SCN��	�JuB�j]ݣe0�����8�S�)�� �c�	����M�^ʻ���i�9��w4�|@=���S@콒���S��9��ܲ�{�4l���빠weʛ��2BD##����M�)�}z�h��>�\��`�pR(�4l���빠[�S@�t���0�5�!�O"��>�w4r�hwJh�M��A6�hX�����6���V��Lh.V{Q̚,gn���g�kI�I���9��e4��4l���u��>Y�U%\hjb�L�N�`s�x]DB!%�J"*L�vXw��nYM�v!X��S19�73;ܵg����guk�������\�SI�M�O��4�]�ܲ�{�4l��Ƚ����S�9��ܲ�{�4l���빠w�ĵE29�Q����s��+��{e�bn8�P�n��ݖh����ܦ�tpP��@�t��m��>�w4r�he.U�0m�9r�S@����-�)�w�S@��u�<Cb�i9l�9��Vbǅ�DD)J"{���m��˖���JO�q�a�	)�[zX�zX��9��V�=���4513&%��@��S@��hw]�ܲ���('��:��J�
��\�.���c���ꛞ��eq��hܱ(�G1
Ed�l�p�-����s@�,���t���n�m��m�G!�}�w4r�hwJh�M��;����i��h唰9��M�;���>��Vg�K��L&IA�@��U�^�������@�D� �����'$�e.U�0m�9#�-���>���>��hm���lIn���kv�s�G;0ۛ8wB��z�6�l�,�A ?��"3�E!����m%4�ڴ�S@.\�1)?�q�3@���z�h�����s@�g��¹��̘�4���/YM׮�m%4]ؒ��3&8h�����s@���z�h�-�4ډ��'�r�]��(�����zX�xX�Iu���;�p�@!�UN�=�vc6�͹�GF�Z���ps��v��:;��w[����ܖi�3���l8����qe���VN���f���\1�N��.�\k���흍<�U���ӵ��q���C�&�8n�#�-�`xj5�c���#��}��R�2�<m�Es�w�������kk���yu�kW����i�
Ĉ�2�����/�j�I3�NV�9�N���#�i�u�&h7/H�������Bz0�8��񗛕!�܍�M�m�~쟍�e4�S@�빠r�X�%�e��%ʦX��(S&�4�nh�Jhe.U�$7j)���=z�h�Jh�)�}�a�6���Ȥ4^��뒚�e4�S@.\W*hpĤ�i����Z�e4�S@�u���~����g����<I5�0Fn�ۢ�wh�zƝ�P5�EtKץ�w=]�ك2b��hu��/YM��s@�aV�˻N�#S1�dQ�@�e7�͉(�+	Dj+�` ��y��m�������})�v\�P6�M6���4w]���Z�e4�S@��,dN3��0#��^��@����z����s@��p�/�"JF�
6E�}�R�ԣsw��w3mX�fM���-TRC���@s׏n���{ng\a<P�Lc�7��Y����sϱ]���0V�m��������z­�fA�h�Ш��V��Z���ɹ�ٰ=OƁz�� �q\+�JO�q�`gq�6;�6 P�J#�
�kvՁ�͵`rW�8��Ԫh�5.�s`s���z����s@�aV�˻�RF�cdȣ��z����s@��U�}�S@�z���ئE�"Gd9��u���p�Wc/jQ���nKp�`�,�����dmD�o����=�w4��Z�e5.Hnnڰ6Mծj�ctEM4��/;�hu��/[��{��h�.U#�S"$�`��=�e4��h�w4]U�e.Pų r8�r(�;�j����Ved�X8Y�IG37����;�è<i���'�9����k���w4�(3ii�����ܭk�!z�p��U������rN8�zq�,=�|Ѻ��]��W�����l�X�<,�e���-X�������L�QG�}�S@�n��빠Z�@�>�l�H�c�28�^�s@�u��-�U�}�S@칙rT�K���T��5a�Os7����;6~ǅ��%;��VI���QLm��9���Uzz�h���=z�h�G�kcc�119*�
�
u�v�1�9h�[v!+�z�k�g����xwjwNs����z�ӡ�n�5�4�J]:��>���zו���ٸ��c2v�c�;cڧ̺v�{���q6�a��v4�ܳ��v���I���WnS��˚r%��Q�pn-հ�薛;<v���~��C�]s�V���B�GvW
���6�\�[�u��P�Fz��{��ߝ��>�#����L9�˞�=p����|�u�um��C���k��J`��m�S�RE0IE�{��h���=z�h���>�\�����Ƥqh����L���V�ٰ;�fM�ϨGPlM���'�9��]��Zyڴ��he�pW�&19%5a�wv�f�������V�ܵ`|��F�rb�1��F��;�ՠ^�s@�빠[b�@>��+p�H�}����M�P�lSe�����I��Ӻ�F�tl�$�(���QH���h�w4lUhs�h�-�4�#f���g$�>��|E�@!A�UP�(QTf[����ɰ>�e��f,���"?�s9�����v��n��빠Ur�R<D�RH�(�Zyڴu���]���V��R�=`9jG����׮��b�@�>�@�ISY�8�F�W��ͳ�1���* 1����iDG^֋p��0pk#1��s4�]���V��}V�׮�v\]��?�1����b�@�>�@��s@���݄�L���6F�Ҕک��]K�;Y�~�_��_R��$�d��RڲI�
�,؝�����8"�RD`�	7�Ie4��F�X�0� )4VF�%.�+�q��J�m`	"�7������H[t�:ZK)��{)-x0n�堓{��%N'64�)ޤ֙�V:��Ea�y2����T[�4�1��O�ٽ�(�2X�$c��MSu�O��kRʴm���R��{���<�c�ާ�o��ah�ᡃ�R����	tki���TIutI�	5�6-���#cU!BYHV�%�)�(R�Z��;4kWF���$�͡���$�Bm��kl*J�.����n�ٷ�榘�.��Ih�?8�D� 'Q��T�+�O�G�R�m@ڣ���C=�߽��wX��=ϰ,�)��AD��;�)�}z�hz�V��}V��r�@����0MŠ}z�h�����Zyڴ�ι"������9nMuԜ�:B��N�<��;�w(!rg���J��6)�&�$&cN`G3@��Uh�6~���	.HwsmXN�ZۥC��j5��v��]�׮�߱�M�L�-5hQW@St�u-ӛ?_ۚ�]��b�@�;V����PlM���&
L�=z�h�Zy�גh��"��Q�P!!"B"F$"T:������$�x��W"$ic�����V�r�����Z{�@�6�i�2"Ad��ֹ;;y	�cn��L��vh0n�%�v�۫�c���6�1G�$ƲQ���h�ՠ}��Z���!��;6r�4��s-"AE"�;��@�빠{�Uh�j�;.[�i�Jbo�9׮��X��;�ՠwt��ȶ���d������U�w��@��M׮���e�<dm!H!��Zyڴ��f<����V;�rl�r$DO��hD��0�D!�"!�j� ���X�a.b�$��u�ӒI-��svKd����WF��!�U�y�7	���<��0R:��r��-u+[H8��nΝ�8܏Mev.��vmL��m��)���,λ+h�S*z�u&x<N�iy�7cTu�w_�;m�~+g�8��[��\&+&�y��M�c���8	��]�c7>S=bz+9{Vc�p�u�ا�Om����߾�{�;�����߂qj��Wl��^���r�n�Lm��s��m�6�I��Iz�/$�F��FH�~�ߖ���s@��Uh�j�>�0����&I"�=z�hu����Zs���x+��&H��#s4��V��v���Z�]��-.�d��@J5��v���Z�]��U�{�"f�:l���K�����ܫ��w7��w�-��Z�u���q�C��@�u�@n�z<�v��E����d�i�`^բD���obo�����s@��*��h����r���d��T�:j����&���&��D*$ �A�D�%)B%-��)�)B�B[ �`@�YP e!%-���(K)(r]�+�6}Y�`}���R��2ubْ?�B�j5�k��hϪ�=m��>�h�\����L��8���h��h[
��j�>^è6,Bs
H�[w4��Zs�h�)�Z[��R4,n`�81�/	�Y�@g�Ar���ܪ�͑�n9ѫ�1�x)��$#k���>�h�ՠwt���n�喗	�x����.�s`w��7�"!L��zX��VסV��>O,�%3	�@�t�}��a���$�뾻Lm��ՠv\�P6�F�x�
Hh~���߷x���`w��6	D)���`d��?D��d�������Ы@�v��������ꄵE!!�z��\l=�Bܚ��B���n��s����u��iLy&H��"JdI�ȴ�j�;Ϫ�=m��>�
�e.PMjH�#"��;Ϫ�=m��>�
�u�����6����h�w4�B��e4������$i�$Nf���U�{�����M��������;~��-�0�4�0Q�-�e4�Jh�w4�B��>�݆vX���h���̓�*v�j�j���cvP�����q'KY-$���*8h��=m��>�
��)�v\�P�yCx�
Hh��o���H�k��3^�~���!%�ɒn�٩)64�i��Ձ�u�́���ͅ9�zX��VӋ�n���e�3R�\��<,�ׅ��fZ��J"'���́�����5�$S#qHhz�h��h�Zu��3?����\�FIo�Y�^�|m��m��Y�p�}��œv� �tz�Y�t��۔��{[�=��wmuԴk:��z�UĖ��;`�[F,h�b��5���p��;f��=Ҽ�;rQ��ҡ't%�!n\���n��t��b�kb ��ݞ��-^���7n���69Aw�B�Ÿyq��9w�^e;lx������m�O;چ2����e)�M75H��|�%wE���&�C�
�趃cX���^v�����]Ď�Ø�y�65�G1ʚeML�&�K	mt��Ձ߲*��)�u빠��x/�&Fc�ә�w�Uh�S@��s@��s@�˗h��`�j-��h��?D%=��Vw\���tP�'�H)4�w4[w4�����h�-���!�LB�4[w4�����hz�hy�B_�D��[��]mY����C�z�����w;�mɎH���ƹy�/0���r7lW|z�V���hz�hm��>W.}e�+��\�.��m��_�8/�cP(�Z��H(D�)�"@��`�X
#EJ��TD�%F�H��"�lcP)a
�S	D�T(�,�wj���ڰ;�9ɰ=��A5�$���!�u빠{�ö~*��\�d�O�~��vI�{���!H"5$�[~ϾI.��ԒVݧ�$�Yu�I{9T�x��L�Ǒ�3�K�Ÿ�$��i��%�]F���߳�IWr�q�I#��D}�ˉ�(�ڴ�t�����0����N$�N��\�W��`R�������? ]e�jI.�g�$�u�qjI/�pcc�D�a 7&}�Iu�Q��?��i[}��I�߮a2I&���n�'����꨸쪧dr�<�I�{�7d����$� �2fH�O�I.��5$���c��y#G�N`)3�K�Ÿ�$��Z��$�˨Ԓ]�~ϾI/+�6Eɍ�L�5u,�$�o�}{�I������I��~�Ԓ�n-I%׋��#Q0nc���;�����f��x�v�,�7;�ku�z!���	��R8�bNO�I.��5$���>�$��[�RI/���H^��M�1Ha��F��]�g�$�u�qjI%��}�Iu�Q�$����*�!c���O�I.��ԒK��}�Iu�Q�$�{���K.\h���nO�&�ũ$���vI=����I��׻$� .-&���B UB{���ym����N�y�E�r}�Iu�Q�$�wY��%�b�Z�I}m�|�Iz���أOl�2e�ƹ[�Ӏ�lc��G�vA��m�t����Ϟ-r���u�(� �����>I.��ԒK�l���.�RI|�v:�'�0�m�m9>�$��[�RI/���K���I$��ϾI/+�$�LPJdI��ũ$�����%�]F��]�g�$�u�qjI/e-17� #�B5%]��'���<�I�{�7d����$�/���H^��M�!Ha��F�������I�%�߲i6I$�߿^�{��#�$��G�����t���0�x��nh�/�N��8D	!���	�����`ˠw
/5R-_E M�bK��w,�3I�]3qB����HE��&��:0`@M�3f�an�ka5��݄���7B���$kl��������D@�d�1����V�r;n�Ax�YE��VQj���F�B�Gi,>wv���ު� �J�#�0٧T�V]���ֵ��6?�4�kC�@M�|YMo���h�QU��+M��B�(e(��t��B�Ĉ|�Nw}:�j��J@@!��6H�!M��f�	`:6����H�Ј����5��>�&��(��+@rB(�PQ+CP��ʢ��>F&Wa��3��@�{���J�M��kca��
��<��n���;������Yl� 	 -���`�    ,; �p	$      UT�,X3u'X�̣�R\b�ɍ���{rK�q�vf���^
�ZUБ��/����4i�[1wc��Ioc�\�����ck�M��(�)�7��0�����{�u&s<�ۍ����3�vԲ���Ѵ�<�u���M��$���ogH�m;��a�9}���s�g��(=D�)z�����<�k�ˬUbhqf^�ݒ�-����+:�n9�x����8�6��]��'*S��^I��bV��괁�ʂ&u�.��-F��	�S���[k�i���:��F�+�9w:*��J�T�u���{(zg]+`��f��:t�[Ʒ�j����-�vMֹV�W��վO���{>��ix�v�`��֬�plf�͹�y��9�ӌd����l��%ö��}]g�<e�g/9�hr6S%u�r����P7O;����c�6�r�6���v���%�*�ݙ"��p<��rm�x�Og8d�fU��
��X%ەS];��R\��)2�L�q�n��2�;�ed�6�����z���秬tsˌ	4s�<����5�z�6p�4�%������x݃�i�yF簡���X�+>t�[v�l�ӡ�u�u���0<��{Fu�������v{Y�D��P�3i��h݌���gYN}grU��YP�!;�[�� ;S!ceL������PI����e�ayx�Xػ���":�c]u�9�bu�i�Z4$���H�VK����m��ae�[kr2v 7^��ΖkI�Ip��)��l���8sPjg�4��ۡZWx�J�
�F�j3���HT�iv�}Ϧ���t�c'��n��wj9yN��+�v���ɹs�H&�l�e�ͻ`���GZE4�;�h�g��iB��h,��9�j��,'%ֶ��kk	�l=5�9��n#Zƴn)�u��]n�}U|�tU#��DM!��Q�(p z T�HH-������S�wU�Tp;����ې9�z�������n=mv��`��>�5f���<���D�<2Y�$�'d��(�CFj��%h��n���g��wS~�E���-p	lld��au��Y��l�����vw(�K�:l�x����5� �i:h�x|{8���5L����u�\T�tp��1C�4mv�vۖ݃Ar������Gm�7%�IY��]����{�绽���i�#�F���q%��T��h��;7�n9�$��\=�t(�9�F�ɧ����ߟ����>��_[g�$�Yu�K�����$�\��c� ���M��RB_[g�$�Ww�����}�Iw]Z�I%�NlN�ywC�w�$����d�Ow��v�U_}�&#RI.�ߧ�$�e��ܘ���1
Bd��U{߿q�$�}�&G�I'w�^��E}��i2I'�~��҉E]6����ٻ$���2<�I�+���������	�I;��{��?�~�K�v^e2��Ǟ�mr��s�h�v�	'�,��z��L,O&��������]V�����G�$�w���K���RI{���|�]�V�RI{)i���RB;��ݒO}_a2���1���GJ�Lo����ӽ��{9yg-�Nﾽ���UT����G,��Kn]�$�{߿i�$���2<��EUO{��ݒO�W�&I$�=$���eZ��U��O�U����<�I�~���{��	�O�*��߽�|�B���?GA9?��"5$��~�vI=�}��$��}��{��y$�w�����e�{t۬X�d����n��k�����^4�Ӻ�cF�t����ܸ~(:��r���$��~�d�N��vI=���?�%��������ə�^^e�T�J���˲d�N��w�UT���yI$��~�>�$����$�g�Oa����,ݒO}�<�$�w}����$-@�������;�s��p��ۙ��N��~k�����'Nhr\����~P(������$����$�o}���N_���g��������������X������7;�I���4����ǽ$�~�Ǒ�N�}�ߟ�����|'Z����ہ�(1!��]Y1�����*������U�7!L��'0Ԓ_z߳�K�t�jI_�>��
~ �~�������o�,�?��˗N�n�U��I��G��_��#���{?t�m���|'-���ӽ�S����z����<��P5�WF� ����n�'{����@�������I�c��I&���EJ�U�]�˗vn�?!"���b������9m����ӽ�ߟ}��9m��$�$T( qЎ�(��%}����L����.��H�U4Yu*ǒI7��M�$�����c�$��ߴݒN�׃�$�|}�wwM�U��i�u8���/��	�Em�Vݘ퓜e�˞7Fr-Ȯ\\�ȑ����w������|o�'w��vI;�^���rO}����U{ɦ���ت��乙����9�%�Bm�o���fg��qs�3?w,�/RQT���~��O��#�9�8�}�Iu�7RI���n�'{�yI$���n�$�O|�i
GC2��4\�����P�s���$3޹�`}�rՆ�����x�-�j��3-�KL�j��3&Ձ�^���|������ٖ��b̺����������d������K������uu�;VV��sZ�	�m�q��u��}���z��6�K�N��5�s;l�fM����;utl<�ݬ���5t�]���"m���Z��R;rn��-|`�k���z����泍��kL*�\���#�sv7X�Uԏs�e�[XJ�u�$Zw(َ{�z�)�b���7]k=p��5�'\��pn�Ŵ�"�j�W;Aps�W+�M�g�<1[6�ހ8���۱��u:��\Q�1�t��T������ǅ�ϻ��	G��%a��~�Vz�5�i̦�r6ڰ9�x_��EQ��Z�3��ڰ>�]���B���m��ӆ������2mY��~�HQ����=��,��х"�r�USTKj��Q
������?;�Q�A*���V����l`�NUP�Z�>�<,w%4u����s@��jkI�s֮�, ���'m R鎎���wF89��f0��8���BⱮ5ʩ�ӗMKsL���Z�>�ɵ�����7�Ł��w�UH�j���s4���Z��J2�T�Qי6����ǅ��P���B�a�~�~_�I�n�Z`��V���mXw~Q
<��!7��ߦ��~�j�9�,MKr�c��K��j����9�̛��Z����J���~��=^TM~t�M��L�9�̛��I�o�����6���﫹2�i�a4(���r�ˮ�Z��D�w:�6��.C\[]C�N����t�}��s-Xfdڰ>�<=о��׽6���ҩ��U5D���2m_�P�%��B��{��X���l�2Ձ�VfL�d���������hs�h�*	�� ~C\��߸rI������,*jn�7T�S�e��Q�P�'����`o�߭Xfdڰ��S�������f��i��2��9�>��V�	~Y�z~_���`s��6t̰��n�ێ[�x��<J\&{��[��ڜ�s<�r�l�29�ƹ�?����|
R�j�6;���s@��Z��Z[w4�\�Է)�7N�9����fM�Q航;��M���Z�>�ɵ~K�EQܭJ��T�M��[��^���e��̛Z��h�:���x�ɑ��섧3w����ͫ�ɰ���BR��$�"T�E�BBB��BJ�@> /�;s��^I2�٬��x၍��)3@��nh�ՠ}�ՠw[��^w�Y$�B4�Q�"�H8]D�#'D�.�s�޵�vPx�e:�����5�i�L@�ʪK\�[�`s��6{�kRQ���j���*jmT˦ꚪ%��9�̛�D)�3vՁ��V�Wj�������$��LdȔ���~��=�ss@�v��v� �UE92-���1�V�)�f�+�[�`s��6
�n�X�j�Է)�6��y3@�v��v�����גrI@t�FB�dH@�XF��$��d%�߷����9Ci��uUJ� �@W[n��c*G:6�V�s*��<�z��ӂX3�k�=��-�8�]�쮺.@]#��p�+�ՅN��F��o]unܵg*���]%�g��p�u�䶷MƢ���o^�t擃<^�X�nzx������q��[K]Ǎ۷7VlzMƛ�ٲ�
v%.����v�U��Ͱ.f�E�u�<^w7Wj�=��m�j�a���xѡk� �k�
,�X����]Sdۀ�L�Hz�Z��?��w/�m˅��Wt)G�m�����w[��{��h�ՠv\�V*���MRi�S��̵�(^����7}a`g�ޛ��ɽ��L��v�h
T�m�iI�[�C@�v��v��̵`g՘�t�Q2ئ�S(�Iz!%Y�����׽6{�j��(K����,�T�ک�M�5T:e��;V��n��론z�M����Y��gG]�+���:�c��rP�;��A�y�65�G_��>x�Qܥκ�d�u�����ܰ�>�xX����ʨ�H$2d��}z�j�D>�Э�-�]3ZBhEe
�&�heQ*��N@UPS��B���)�Fhf�P�Tꨴ���JG7�����mX�e�؄��w�j[���mҧSL,�,��ʳ�B���ݵ`}��>���&�*\�i9�t�(Q9]ͫ3vՁ��XXy$�N�ޖ-X͡U5UJj�S-��3���$����p�zX�����	U�D��"J<$d3��˵i4s�B�
��Gm�a�۶�Pۮ^x���<�sRf��n��z�h���(\��ݵ`}��M:i���UN����ǅꄔɓ��`nnڰ>����(��4����p�9u�@�n�����&����T9T�&a2�7���	�މ�y�i���JB�/�����M���Nďz���M����D���v��lbB�)�K��A@#�X��a��L{ �����w�2Zq�	����*���Xp�����2�Fٽ1�u����d%>'Ё��M	}�� ����0���vq�|e���!N���}6��8�����k8��Њ�����#�b�����4�Ri��^pO�;M��f�VP*���e0MK.�iϠLhN����<b����|#bi�e�׈��-]��}�]R$@9߆���HS� ��'Ez b�U>�	C�'���E*���F��E�#��_���~4/b���)����:��D)���;��w��J�߿= ���R(�ɐnf������9u�@�n�z����M7�Ӑ	�P�v2Q���լ��Wc���$.'p1�������\P�*��p�zX��U��̵�Q
>��{�r��Q5J|�I�ӦX��U��̵`}��f</RJ&LZ��-SmS�5N���Vٙa`fYM�uzgYZ�c�F�4���
'���X���;?w*Ð����
f_���+i�M�mʪuL,�xX	Nw5���V3�a����{�߿�����O��	� �7-��ֻ�8���596�z���ks�v�������� �Q��ǒ8x���&�z����C@�e4/b�$���D��@��Z�Q	L�nm����K ���`���H�H��&A��׮nhׅ��%2gs]���j�>�KsN�mF�L�-����4m���������`w)lU4Mz��Nf�2�;�f�m��׮nh�����1�
L
"!���U�
��wㆪ�骀�m�=v��'��Vݺ�����q���e^�{G[�9�{��U�n��0jgu�6�` ���6"i�Xz�?Dq��s���o1��k��"d�V�n
ڍ������6�7=�#N�-���p<��O�ݞ�B㶞bӆ�ۖ�kDĘ�aƄ�:x6��lݝ��|�6ts�<ېy�'�x ����e��!EՍ���!uN\wCrg�m�c%E��c��]B�[��#lۋ�����
!J��r&Z�ڧL	t��~��֬�\��/YM �u���̫��USU2ڰ9��j��2nk��3����̵ȅ�
*��y[M�i�D�b�uI����`�����V3��X`�R�UN��MR�L�؏���;��Z�9��j������~S�&hD�T6H�[n��̵`l$�ۺqpݟ� �u�u����9#$2�,�ݗ�ͮ����:��4�a�ݞ��{.�Ѻ�H�85L�s>߿~74�S@;�q�#����zՀf��5-�b�l��SCVw)G�	CH�(P��
��ǚ���V30�{	%䒪;��*��Sꪤ�Kt� ��;;�j�$����t�`nk����,���ԶӚB�m�qlD$��!~(������߿\�~�L�}�`q|���TR� ���2ڰ9��%��(�B��(����~:���`gs-X:���`:
�ڹR8�c�Z��Mdˮ�q��wZ�w8��L,OE�)�d�O�9n'�^��߻����Z؅HQ$B!	$�������QV�sM�R���߻����Z�9��%��ǅ�Q�!!B�BIU8��UU�R�̎e��o�j��f\�LB�B�Rgq�`������g&D:eK��*��ԔG��%IABB�P������������vv�� �.LP� ܃j4�4�Y�&
!�@�$ "�*�����zՁ�̹,�b2���sRꇷU�쮆��F��H<���`��8�v��dS$`L͉`�L�Ԏ��4'���9$��Y��~ �$BDDB���=�~,[��)I.Fڤ����w4�������]�T��Q� Du���zUR�b	*�s-���\�w}�h���;�͘�����c�kvrL_�M~���9$�����'���9$JbEU�D�����{�rI����TU�GM�j�:e�g��`lDBK�$�DB���/��{�%��ǅ�߰��f�'K��݆\���9�\��n��3J	��.�2�=���_`��7`gs-X�˒����TD/!@��D$�����-�>� �.�Lnf���Q�^����4��o�f(�(Q���&�|~_�R���:&��Ӓ�����`����e���rX��b��Ect�N��2�b^I*���=�zՁ�̹,�xX]ŖR�Z�m:�)�݁��j��
!}����n���;�q���gJ	�n����}����5Q�
tv�9�4;W0�c��?��׏�sv��Y��^g��mG��h�t��Ul&hq��mcJϕ���<�z��7����;=����Jg�;������5��Ң�1� �mgoN��u��2�᧰��X �;[/;��F9h*i�(q�l�2� \�ǈ��M�9ݗ�wn����[�4gu鷵�3Ԍj9ӱ�n�!��a:��nMn���Cl���<�rc�FO&���W=��9xmؒ��2���v�31�`���
!~"!/�=�zՁ��+��r�i�U9�%��� ���`ffZ�9��%�B��L�jҨ�D����&���v��h[u�S@��+q��%19d�2�vȅ�
{��������ǅ��Q3��v�'I�� �.�L�j��f\��DB��Ӏ��`e�s@��+jF�F8E��p`�cܫ[h�+˞^B��ooF�]�]��<t�}$h�G9�D�Q�@��h{��-�s�B�ۛa`}+"p$F���e��~}����!�� 5�����ٌ�ws@��C@�e4ιth����t�4۰;���gr��(K�"!Uo��X������
�4�Ỉ9�ץ4�S@;�f��������+1n�N��[sT���c��w�����ץ4�Q'����" i9����#.��az��=�n�9˸�oG������}�?v4�\�����z۹�}zS@��f*����,��[n��3-^��>�?���@;�f�\�������L�j��u�`w��6|��!Ik)�hB�
BѠ��c--�hBT���X�b%	 �i$!H��P���V�����QC�{}��I��f�{��&G�dȊ������Z��4[w4�Jh,�����H�2]:nl�w��$�wwx�ۏM�ڴyڌJG��Q6َ
�)9.j��j�v��ưw/�<>�t�nN����0�����ץ4]r�DB䁝�v�Zж�U1�SQ�3@������Z��4[w7���J�3�[r9�ۚ�M�Nnրw������ҚS.Q�`!�m�Nj�Xy(��"�s|���k{�����$�ĸH����mco��⪨	hr�Ne���2Ձ�(�D(�Ȅ�g�}���~�V߻����߶��t�<�aPV��NȜl��s��quJ�Zi�,�vy'6�\���d:���}zS@�ֽ �u�����LX������9����ʽ�	/""U����zՁ����䮩;$�Ku.��u`�q�fe�5(J&~�zX9�VWqe�$�Jm�Х��?(P����`}���;=̫B�3���Z���J��&��u4Ձ�ǅ�興����fk�>��V �U8Du��WD�t!g��.��WZ F`A"A�}����!u�a�| @ֆ	+�1I%�5��Ca�Bb@�bDM�Pѽh��P��!":�D�@�����浦ki�uu��CaP�R�)����$Jiq�2��\Q��CQ��`@�aĈā-L i�d!���wor����+����l����E[dřr��5B7;J.6%�
�Z,UtX� m@�`	     q� [N�       ��Rl&H�9ʜ�u�q���mS4������P�!��U��F�rf�s��:����cg�p�5ƛ{6^Z۵7&mەꆮ�)�CF���A� �<J>�;Eam���q������.�U�]��؋Zv�2�� ۙi�q�\��N3�k�GQ�=,ݹ8zvn{O�3���1�6�6�Ӱ��SFHٷ����	�0��y��2���S��]o\�2v�`IGҩ7+T]�؜��e���V\�;^�.��텃ll�zJ$��6��B٤I$�&ԓ���e��� �pJ�..rJU�l��eU٭�tUWY�Ce��`"G�n8]���nڱǩ����d���f�t�uݮ����X�I�q^˜���� �=���.��'[�eyU��1�f���ufD�vɤ�.)�J�� �#nvq'9�;v9ɲh瞱�z��9Ogu��
����=Y[n1��p�\�W�^H;���ʵ�d�vÄ��U�Ƽ��g���R�ø��Vj�n���M�<l���܌����Kv�I�t�([���c��|v�:i�<�s�[s�/M1g�0ce�aS�ܓ�)�������5�fY�vv��ΐ�:v$�	ji���:-��;ۗ��[�K��<��,y���;���5�vL������UY.�7c����c;f��n�����r;�`�kj66�v��Sƽ��X��ղ��	61�1��))]���]��,�Z��l+W*ƧbT��UF�{����kj�@���x�}��5.̛-m��g��ڶ�R�Ye�n��� ��t�W;{C��t4
/k��9;v`9�݋�X����s���q;�#��q����cN�t��W/�q�n�S�UU6�8�V[��Uv�I��&�ݙ宲tw:�DV�^�l���!�[հ���P 0Ё�>�
*�Eҏ�z�W�����B���?����kō��U����m�$����(f�kd��\�uk��9G�\i��'����T����.'8�@y�'eLn�8�d���ԫٵO�:ᳪݎL8�=�;p�\�r%vY#Z���Hn˴Y+����C����<�qn�c��u�ë5��{�mS�@���Z�4kJy�hsB
�鎣ѝ�s8���:��f�#�
f$NH���؝'ZϮ�/Rgxެ9��3�S�nx�#�)""S�Iq�x�Y�ݎ��3-z��H}���3E�J��TG$���@;���n������w�/(IB�3�"J$�Ne���6�o�j��c����eX{�v�����%�vI
�ܫ1��B_� +��<X����;��3����1V!�DA�q89���wY�^�s@��M�}���$hȈ���]��*���kk��f��:^r�e�u�s�������5�F�F�a#rG����/[��}l��WZ�ιthDC�I2{��$��{����K^� KJF"�+#  ����"@�:Tꁂ M�w7٠r�����@�vXYYۘ�i���'��f��;�����ۚ�[�)""S�Iq���j�wY�^���n��˔y�$��n�)���>�q���[�zp�v�@��Z^%Ƙ�I�sja�d.��nz�k������d�W��3�$�n.�9۲�!L�A�M�4�S@����/;�)�)b_��o�ؖ%�b_��Y?Qu�$*�r��5�4F���~���,K��g2q;ı,K����;ı,L�s'�,KĹ�j1��j��*��\!I
HRB�����Kı/�{7��Kq�ԃ`B"T����|1B��Q A�CF��@ &Ћ*u>���5�~�'�,K�����#Z#Dh�GџI���XK�����,K?!Q5����v%�bX���?N'bX�%��ٝ8��bX�&{9��ؖ%�bx�٢ۻ5��{��{��,K��g2q;ı,O�����Kı3�̜Nı,K���|Nı,K�o-˻�w4��;Q�u;P:��ڧ�^X�ַnN��ݝ�9ۮ^|�����m�nR�����7����ΜNı,K=����Kı/�{7��Kı33�8�������[����s.%�5N����ı33�8��bX�%��f���bX�&fs'�,K���ΜN�y$��(�!Q
HY�<��U�nMz��v%�bX�ٟ���Kı33�8��bX�'�ft�v%�bX��̜Nı,K��f�K/w,�ѻ�o{�v%�b"ؙ�̜Nı,K�:q;ı,L��N'bX��@6�+w{��|Nı,K�_?�O�]Gv9
���x�h��4|�gN'bX�%������Kı/�{7��Kı33�8��bX�'�nx�M}AR�t�i�UKU2M<d�u�1�ݭP���9�p����-�K���{��s�gM��)�sL�j�|B�����z�\.ı,K���|Nı,K39��ؖ%�b|�gN'bX�%��G�Y���4Җ�[e��
HRB��3]��UKı3�̜Nı,K�:q;ı,L�s'�,K���7�I �6�hR�w�)!I
H[�{8��bX�'�����Kı3�̜Nı,K���|Nı,Kǌ�%���j�[,��8��bX*'�ft�v%�bX���N'bX�%�~�پ'bX�%���d�v%�bX�՚p�܎eæ��5p�B������d�v%�bX���o�ؖ%�bg��8��bX�'�����Kı ���	6A(@� B�"�-)`А�I}rK���n�N.8j� ���v��e��n,�i�u=Ne����v����j7�l�q�/N�r/F3v�!VڕB�6{-�;{g��)�*�]�\r.ѹqm���*Ʃa7��"�lrnnr̓(��ý��%�:�X+lҞ�#�-��.[wh�ۻg�v�Eڣdl[.��p��nr�:諏ocV=v�ltF�v����v�v�j�&����I7����X �Pc �D QRB/{���R�%�;U	�湹nqc�[qd�y<�D�8�z��y+s�vn}��;5�SQ�N�8�bX�%������Kı3�̜Nı,K�ft�*$�Q,I!{}~.RB����"J�S�H��o[�v%�bX���N'`�X�%��3:q;ı,L�s'�,K�����v%�bX����\ѽ�{&����{�Nı,K�ft�v%�bX���N'bX�b؞��i�$��5�q �ޘ�T�I*iQ4U8V	"(dL�s'�,K�����v%�bX���N'bX��������1�#Dh�F~����Z��K���,K�����v%�bX�9��N'bX�%��3:q;ı,Mͽ.RB����@mW*fS�%��ؙшz���ڎCn8�I�ɱ�*[6�8\���*eI �7N�MӸ\!I
HRB�����Kı>fgN'bX�%���d�v%�bX����Nı,Kǌ�-p��]ke����,K����8���D�}x��P�����b~���g�,KĹ��|Nı,K=����Kı>��N˽�eæ��5p�B���������
ı,K�{7��K�X 5Q?g�~�Nı,K��ߺq;�I
H]�5i�n���*��e��
D�,K�{7��Kı3�̜Nı,K�ft�v%�bX���^'bX��=����NW#�(�.���X�&{9��ؖ%�b��"0�#����'Ȗ%�b~���x��bX�%����v%�bX��{?�55���4�un�:ܙ��ڮ�����_e۰�nÍ�c�3�N\�Ό�=\Wd����wؖ%�b{�����,K���e�v%�bX���o�ؖ%�bg��8�!I
HRB��Uj�	e5N��SWbX�%���e�v��0�Mı/�߿���Kı?����8��bX�'�����Kı>Q�g�C�V�����#Z#Dh���o�ؖ%�bfg2q;�j�2F1d"!#"�$X!!UG�C�D!q;>~�Ӊؖ%�b~���x��bX�Bś�&���M�L����
HR~H�D���N'bX�%�����8��bX�&f�/�,K��D�f~��,K��܅��[)��l����v%�bX�33��,K��
,�~��߯�Kı.f~��,K���d�v%�bX����Qm�e�W+gkۮ���j6�,d���6�#���R���s�sD�ů�����bX�&f�/�,Kľ��|Nı,K39��ؖ%�b|��K�����$,�5i�n����'4�ؖ%�b_{پ'a��@�*���b~����v%�bX������v%�bX���^'bX�%����!TCj�w%%��#Z#Dh�����'bX�%��3�8��b䊤���j'���׉ؖ%�b\���'bR����d�&�t��T�j�[.V%�b|��N'bX�%���e�v%�bX���o�ؖ%�����A�,L�s��ؖ%!I
wLZ��0�ST��e��
HV%���e�v%�bX��(&�3���"X�%��?s��v%�bX�39��ֈ�#D���U.�
�%�՝�2��,�x���ݜvPU��;��d����7 u�Ơh�������oq�����v%�bX��ΜNı,K�g2p?��&�X�'���׉ؖ%�bb�x�ԒSt�8�۸\!I
HRB�����?,C������b{���Ӊؖ%�bk������bX�%����v%�bX�<g!k��SWZ�f���ؖ%�b|��N'bX�%���f���bX�%����v%�bX��ΜN��$)!wi�[r9��SN�.bX�"���f���bX�%����v%�bX��ΜNı,K�g0�\!I
HRBNKuT7Rة�\Nı,K����;ı,?�U �����'Ȗ%�b}�����,K��ff���bX�'���k7���(��kp�G5P���1ɳPp�����O]�ԭ��kM��s��;[����\Il��'J�ƈz�*gA��K�}��7Sҙ2��ۮ�,�4��NJ[e�t�qq��ֲ���b���7<�L�K�[��<f��n�\�{;���t�Ui��'�y�&*L䝃A�%�v�s�۷D���K�������ϴ�Dɜ^�rY�u��&D�<�4n,ϧ�\���� Z{vvږ�TWˮ���jW/n֊o{)�toWz����bX�&fgN'bX�%��3�8��bX�&k35��Kı/���'bX�%��OY��N���U5$�W�)!I
H]ݽ-;ªEQ5���߿k�ؖ%�b\�߷��Kı33:q;Ĳ��:j�C�MK)�uNi��p�$)�bf�3\Nı,K����;ı,L�ΜNı,K�g2q;Ĥ)!}K$Y3:2�ӊ����p�$)��}�f���bX�&fgN'bX�%��3�8��bX�&k35��K!I
HX�t�Q3#T�t�Km�.��ı33:q;ı,O�����Kı3Y��'bX�%�~�پ'bX���������3�y�c��r���/���t�;Uc�ס�m��L[nu� ݅w����}���v���r��kDh������#�,K��ff���bX�%����;ı,L�ΜNı,Kd�ڦ��t�M:l�\!I
HRB��ڸ;
�DA���D�K����;ı,L�ΜNı,K�g2q;$)!I4Zr[�T��b�6��v%�bX��7��Kı33:q;ı,O��d�v%�bX����Z#Dh����eQ5ݔ[�]]U�#�,K?(DCQ?~�����Kı=���q;ı,L�fk�ؖ%�b_����,Kľ���)�{$5��.�q;ı,O{9��ؖ%�bf�3\Nı,K����;ı,L�ΜNı,K�=�3Z�ޮ���I׋;`�UU�9�UB-�nݳ��h\n�5��$�{�����}m��t���{�"X�%����q;ı,K�37��Kı33:q;ı,O{3���4F���Ϥ�J��\j�U]�#ZX�%�sٛ�v%�bX���8��bX�&{3��,K��ff���$��$)!j�ӕ@L�-�Iĺn�v%�bX���8��bX�&{3��,h�������I	�=P�*�UҏH	�aX�C�',t�4�B�.N�$�)!����B�B�)�d���.�c-]�v�wq7FmQ�R1�P�HԅY;@�6i�&JV2��2�Jc.U���,�825ED��*�r��,a�c%��HAY$%abD��D"�`�1�PC�'�[�CࡹD�
|C㧊nI]l���l��~�CA�`M��C�M�i�!�2� ��#��a��#��bh���xPJT$)q
4����tv����-e֊M�L��I@�������C�wn������x��lт���  ��O��B��H������x P]�
u��_"' �<)�P0�K5�>�ؖ%�b\���;ı,O3����RkZ�wu��ؖ%�bg�:q;ı,K���'bX�%�sٛ�v%�`bfft�v%�bX�3��7 7[�n�������$)��w�,KĹ���;ı,L�ΜNı,K=�Ӊؖ%�bg�a�j���k]E�!��vU!r3��np��c����dx�n����:�IS�۱q;H��,KĹ���;ı,L�ΜNı,K=�ӈ�bX�%�s?~�F�F��=^�~TK�e%�&���;ı,L�ΜN���MD�?g��8��bX�%�����;ı,K����,Kľ���)�F��Yu��ؖ%�bg�:q;ı,K���'bX�ؖ%�fo�ؖ%�bfft�v%�bX��f�7�n�o[7�joz���Kı.ff���bX�%�fo�ؖ%�bfft�v%�`|QЦ�D*&�=��q;���$/�d�&v�����Sn�p�"X�%�fo�ؖ%�`�fft�v%�bX��ΜNı,K�fo���7���{������
{<�]<�se[�.D�zq��7g��1����F�Vےө%�.����w��ؖ%�bfft�v%�bX��ΜNı,K�fo�ؖ%�b\��|Nı,Kǌ9-�&��5�or��g�,K�Ϲ�8��!bX�%����,KĹ���;ı,L�ΜNı,Kǰ�MSr!�ɪrۦ�RB���w3|Nı,K�7��K�0�MD����Nı,K�~�Ӊؖ%�HY�n���R��*��w�)!I�PR(��k�g��;ı,O߿s��v%�bX��3��,KĹ���.��$)!v�9�UL�4�%�R�|Nı,K39��ؖ%�a�?���É�%�bX���߷��Kı.{پ'bX�%���D�Ъ�;���籿��^����g5PpU@S��=���#���)�v�Z�Nvn<�v6�]pݸ�n��OXWZ�cv���m�rlv���vEQ
���c�#.�M�xuN,r�un�
�3�r&kv����s�6M�6븐��������+�7d�Ź̈́�c��NL�D���ۛ<��n�(yե���kl�q�1ƃ^�'e�=���Z]\nB�.YDuWe���s^��Y꜎X(<�'7HvW{qn�s�us�i��X-��#n}�w�������sX�{�Nı,KٙӉؖ%�b\���;ı,K��o�ؖ%�bf��p�B����9��hu.IN�uU7�l�v%�bX�33|Nı,K罛�v%�bX��̜Nı,K>�t�v"�bX�4z����oWa��Z����Kı.{پ'bX�%������Kı3�gN'bX�%�s37��Kı0�d�	f˽�z6��{�v%�bX��̜Nı,K>�t�v%�bX�33|Nı,,K��o�ؖ%�bx�%�Cvn�Zٻ�os�ؖ%�bg�ΜNı,K�7��Kı.{پ'bX�%���d�v%�bX�~�-�n���;6��;s:+/�u�4��wF�/�gl�\��ݝBѻWB��w����2X�%�fo�ؖ%�b\��|Nı,K=����"A�MD�,O���+�����$-��-�*n[r�.��'bX�%�s���;��H��;���'����'bX�%��߿t�v%�bX�����,K����5
i�i��-:�۸\!I
HRB��d�v%�bX��3��,U,K5���v%�bX�=���,K����}?\%�ʻq˷�ֈ�#F}����Kı3^���,KĹ�f���bX�&{9��ؖ%�bNa�Z:���UCt���
HRB��fk�ؖ%�a�D��ٟ���ı,O߿s��v%�bX��3���{��7����{���#:�X�-b�y�L':ۣ]��t�w�����Z�0]�.��Դ�����p�$)!I
w3]��Kı33�8��bX�&}����>D�K�����\Nı,K�r�D�:n��[n�p�$)!Isog�D�,K>�t�v%�bX��fk�ؖ%�b\��|Nı,K��Kp���.��wz���,K�Ϲ�8��bX�&kٚ�v%�C���%ڎ�D�/����;ı,O���\.��$)!bR܈m�4܏z���K���{3\Nı,K罛�v%�bX���N'bX�%����\.��$)!f�V����ܚ%����Kı3^�k�ؖ%�bg��8��bX�&}����Kı3Y��'bX�%��?~����o{����sf;;��u����۠|�<���]�+�ӶF�us����w��N���v�+����,K�������v%�bX��3��,K���e�v%�bX��{5�p�$)!I+'*�R��i��$�˃�,K�Ϲ�8��bX�&f�/�,K��}�k�ؖ%�bfg2q\"I
HRB��Z:���UCt�'bX�%������Kı3_}��v%�bX��̜Nı,K>�:b5�4F���}�~���K�*�bv%�g�(@�O��~��,K����?N'bX�%��}�8��bX_߁�����et(Q������ �h��ʵ$FD!�X�P�Q#4E�j2T⠧�_�'?{�ɸ\!I
HRBո_�D��ۤ�޸��bX�&fgx��bX�(��gN'bX�%������Kı3_}���#Dh�����˒�U��-�ڈ�}<�䔳��Klܐ�swn�˙ӂ�n�y��8�;��*��.���4F�������bX�&{y��ؖ%�bf��5�� ϑ5ı?g���v%�bX�=��M:`��3M��5p�B������/� �,K5�ٮ'bX�%�����,K�ϾΜNĂ�$���*h����U4�X����ڵ�=���r�R'蟽��q;ı,Oٿ߯�,K���{]ws[6hջ7.��q;İR��fw�ؖ%�bg�gN'bX�%���e�v%�bX����q;ı,O�߭�
j�f��[u�'bX�%��}�8��bX�&{y��ؖ%�bf��5��Kı3ٝ�v%�bX�R� k�������k*�,Oh�c��U����v44[@Y�8�7ke[f����q��,݃]�5�Wm��.��#m%���m7)s�kd�ZAd����KZ�mU���flpA���Zq�]e�mv��i�Wm	�vX5�N�uV���u�fM��"���8���ݛ�E�N�8�&��DC!�s�w�s�jݚ�ækt۪=��;+=��3��ֵ��vfj��B�{�4�;��㘭���H��e��n�.ػ6��{�o�����u7}���bX�'�o2�;ı,L��f���bX�&{9��ؖ%�bg�gN'Z#Dh�G�_O�]��aw%]�F�X�%������,K��g2q;ı,L�����Kı=�̼N�I
HRB������i���@۫��ı=�̜Nı,K>��8��c� ������^'bX�%��Y�������$,X�Y3�9��i�k{�Nı,� @�O����Nı,K?o����Kı3_s5��Kı=�̜Nı,K��'2�{�	��[����{�Nı,Kټ���Kİ5�3\Nı,Kٜ���Kı3��N'bX�%����޵w�yV�@S	��sr�4��X�w�\�v�N�FŹ��o��.����?{�7�ı,L��f���bX�'�9��ؖ%�bg�s'�,K���3\Nč�4{�O�%m��e%��U�#Z,K��g2q;������H��bfg>N'bX�%�s37��Kı3_s5��Kı>f�m�aR��*lS-��)!I
H[�z\.	bX�%����,K��}���,K���d�v%�bX���n�L�tӪ��˅���P��;���v%�bX��{5��Kı33�8��bX�&}�d�v%�bX�4aa�ʩi7SM������$-�ݫ�Ȗ%�bfg2q;ı,L�s'�,KĹ���v%�bX���L� t<F�5�1Q�@nx�卂vԛkgY��=�.�Cɩ�6���,�;ı,L��N'bX�%���d�v%�bX�33|�>D�K�^����p�$)!I�W���@�r��f��os�ؖ%�bg��8��bX�%����,K��{3\Nı,JB����p�$)!ImΔ�B)�g[՛��8��bX�%����,K��{3\Nı���B��A�RU1F��g_�Z�HB@�t ��J@�c�eE���
�(qT�"j'�~����Kı?g�d�v%�bX���r\��nUi������$-�ݫNı,K39��ؖ%�bg��8��bX�%����,K��as�����f�޷�'bX�%������Kİ�0O�����Kı/�߿o�ؖ%�bf���'bX�%���o�zjS&����Rt6!�MSщL7Ug�Ŷ6�5��N$l�=^�v��;\'P��w���ı,O�����,KĹ���v%�bX��fk�ؖ%�bfg2q;ı,K�ٻ��i�l޵���s�ؖ%�b\���;��Q5�����\Nı,K����8��bX�&{9���%�bX�4aa��"i����n�p�$)!Ik7j�p�ı,L��N'bX�%���d�v%�bX�33|Nı,K3ә��u.��t��Iu�q;ı,L��N'bX�%���d�v%�bX�33|Nı,�Q3y��'bX�%�����C�%�UYwUv��#Dh��d�v%�bX�33|Nı,K5���v%�bX��̜Nı,K��w����Ӳ�)��es�3�:��D�F���s��(:�=�hz[]���Wn�`mY��g�,KĹ���v%�bX�����,K���d�v%�bX���8��bX�'��	��wZ��ٽ�M�o|Nı,K5��q; ,K���d�v%�bX��ΜNı,K�fo�ؖ%�bg�[fwz��u)�vn[��ؖ%�bfg2q;ı,L�gN'bX�Xj&�_߿~��,K�����\Nı,K��Y0��ٸk{����v%�`6&g���,KĹ���v%�bX�3پ'bX�%������Kı/ϳ����m5��zַ�l�v%�bX�33|Nı,K�{7��Kı33�8��bX�&g���,K���>T�O��%�,�r�S��6��uXF,H��s�M�8uXE��j�J�Ʋ���)��x(R�!V�!k!+E�)IB�='��@�V������:�[;e�@�E(�"D �F2!"E����'h�"D���$w����ٻ�5i5�� }���.���BYxB�
1H�b@`�$���d	�N2�aIgT��4m)u����� ɵ��m�U]�J�������
�]tS���9��z�v��'�M 8@$� �    	 !�H       IgbX܀�բ�Tp8�Q���7 �n�q�km�����i�e�US�od�n�:�ŀ)�9���A�Z�ns]�b�8� ��.��5���n2���k/���;׻n\��71��t:�=E�1��]����5�i姇k����F,�S���cN�d��(]��U��T�ױ�Ȼэ�= =U�p��v�ŹklT��l��� m�9�I,���c�	ZVveUف	q��G5TN�0e2^p6[,�(l [�S��I����k05W*0�hci�Uu��j�ہ� ���35eUٮƁj�Q�\�Р.@ h�*���"oT���Y��ޭ��Ѧ�+n�2줚�0Nlt�.���񐃶�+���SiC��U��45vٸ�nR�F٫{+�\ai��6��n{[VN��	6P��5�\C��<��Y��+x��U�r�eؚ�"�"9k,lg@ s�5нSkm�Y:��ӑ�sִ�*�Rd�k���E������+`�Üɡ���=�.p�wۍ�M�
���n]�|�Jm��v���Z�#�t��5�n�)
�8�Ձͳ�i��.v���!�x��	϶8i�}��^��G[]]x��x�b�ͷ��j�w�c=g.�x�7qcS��Ϸ9�^�la�N+s@�!��=��eUkj ��U�`�wj�77f��
��/��m+�0g��@%'�mU'd��V��[:�^�� �D�,����-,�m0����n�4ʬ���4m�=p�\����7nU�YW�ö�jh
��K�nyv�܂<��P�|�Hc�w��n�۷m�Mmٹ���qۚ$�:�d�AmY%���.���Ö���-j����du�bu�W�t�ԽҲIg�˪ɳ�N��<m�a����ݵ� Sh�A؁�W��n����k���C���A����2��n���z���/u�:6�p�B8K[����Ǚ�n݇F�c]���d�3��[���́țU��2o�s�d[f�|�n���[s�+����`*��.��s��d�g��A���]�-�n�U����c�������Z�7]��U�-��5�r�ci^gm��u���G�wo���B���eSr6���]�P��ip �����q���wY��9���M/�l�0�8W`D[�6�:v�]\�����j޵���,KĿ}���,K���d�v%�bX��Μ�Kı.ff���bX�&g�0��Ժ7��{�&��q;ı,L��N'bX�%������Kı.ff���bX�&k=��v'�U5��a����v]��[7�k{�Nı,K���Ӊؖ%�b\���;�,K5��q;ı,L��N'bX�%���r����-�6Jn��\!I
HRB���p�%�bX���k�ؖ%�bfg2q;ı,L�gN'bX�%��0�]���-KnUi������$-�ͫ�Ȗ%�bfg2q;ı,L�gN'bX�%�s37��Kı=�&��e�mb��d,і�x�MNzug�:z�v�E[.E�=v�|�U}�����7������v%�bX��̜Nı,K3�Ӊؖ%�b\���?>D�K��{}W�)!I
H]�hHyMM�
�����v%�bX��ΜN	"ŋD�!"EB��0�Q�AZ�B�#�*�DH)�Q9Ĺ��|Nı,K5��q;ı,L��N'bؖ%�;����J���˪�����4F����'bX�%�����'bX�%������Kı3�ΜNı,K�-Ri�*ni�7T۸\!I
HR&k�f���bX�&fs'�,K��{:q;ı,K���'bX�%��p�M�D�lcmn�RB�������Kİ����,KĹ���v%�bX�����v%�b]�?���
<��tv9�Ω�sƻ=m��G+U�׬r�aGc[z��nʸ��P��-�ֶoZ��8��bX�&{�Ӊؖ%�b\�f���bX�&k�f���bX�&{9��ؖ%�b|>�.j�{�r�ro{�����ؖ%�b\�f���ؖ%�����'bX�%���d�v%�bX��gN'bX�%��0�]���˲�{�����ؖ%�bf��k�ؖ%�bg��8��cC�H��+��R�`h�7���:q;ı,K�?~��,K���M+��t���MS������DB�����N'bX�%��3�N'bX�%�sٛ�v%�`~Q�����ߵ��
HRB�i{�'�SE5B��2�p�ı,L����,KĹ���;ı,L���q;ı,L�s'������oꔈnyi:�m����r��<��-q�Ǉ.�s�ϋ�;h�ٵ� qXQ��� �~�^�����{���X�%e
���lM�۰2~̫�S&�,��V��vgG��Q4��@۫;�;ܵf�(�77^��w��@�r���8�nB6�4�rՀgs���eXZ��V�*P�""$gs�,���Sl-���5���^�����{������7Mֺ����V�Ķ^Nt�s"Pq�=���gY�g���:󱪹���&�W�zu��/u��>���=�ň�`�����&��=��/u��>���*��@�:�.2A��1)�]��YM�Z�{�4�.Yq��Q5���>���/>����,6!BS���>��P�ENi�Hd�$4Ϫ�=��/���>�ߧ$����%�)D��@�) ��RQ��#�ТF26ԁ	IX�X�b4H�$�b��1"0`�����W���V�J�v�bu�:�^�NP[M�&�n�\����m�}�?^���,��d��l�F���z�pΟ\j���h:VL�1fr�O;������<�z�z�&��v�W�v��P-3�n㫷dRsn��o4�,�6�/Yшs�ܞ7cq]����*j�;c:5/( i�.;n�=�����y�Sv0����8�K�E�F�d��w�{�g��Og����G�+p �nL�Վ
��:.e�x7'���Ѯ����	��P�`��@��_[��}�)�^}V���캚�1(br�!�_[��}�)�^}V��t���P�S&.����t��9:j������h�Jh��hr�͑��)�H��$4Ϫ�=��/���>���=�ň�`�����G"�=��/���>���/>�@�u�M�mg�@���;w&�Ou�m�v�L�Q>��ڻ^��Cn��n.՝�n
�m��w4�e4Ϫ�=�����R:S�j����u�� ��;#�j��D��pC|��NZ���DKٜ�|���S@�빠|�љQ�)���>���}ׅ����6Ձ�u�`[Irn8�$�)��t��}�s@��S@�}V���캚�1(crE��/��h���/�U�w���o��x��tAMj�vm��ѩ11�k˪s��:�3��x�Pl'\N�vs3F��7�I������h�)�_u��:�˛#d�LRE�)#�/�U�w���}�s@�^��"����)˖6���}ܵd�R��B�
��J$Y��YV	BX�AX����{\�{���J��6P��L�Xl%
w��f�������h�)���0�J27��y^�@�}V�޲��]����'4�6A(�pB�F{7A�3&�5Ț.ź� h{#���F��ӝ�2E! B'z�����/���J$;;�V�SS�,m�fE�w���$^� W��9{�����Y�b��9"mHh���
��@�YM9�&���j��s�VNfU�߱�a�.�QJ��S���`f�X����5-�U2ۭ�k�;�S@�����z����Y��nzn:��x⬝#��s����؁ۀN����]ts���Zϣ��#?{��h۹�y^�@���,���qD�r���m�����
��@��^�}���q�!��#q9�����ՠr��@�n���FQ,�IFH8��/;V��ֽ������i/�C�(I0�E�r��@�n�z���j��;��ٻ[�x��UJ� �nf[L�tR��H�&�j�y�a�i���Iz�j�LH�9�n݈1�-��yz�F)�I�l���:N�B�f��q�qٞ�m:�]���<dc\�������\E�`���=��4�:B���uK{%��u�f��E'on����@l�;��d�z���$sVP����ty��eݹ�'Vu���H��׶md������|}�6��$J�n��G��smy%��$<�w;��TӵۉG��R��,N*��Q4ۚn�X���׬�/;V��ֽ�X��Ġ���C#s4׬�/;V��ֽ�]��\��D��b�,b�M�ڴ^����h�Y�{��E6��qE�Z/Z��w4׬�/��@�Ρ�W��1�dn=�]� ��4�j�9zנ^��8��Ld-�D{t����p��J2�_7;p��Ck��&I�8$6�dn73@=z��ڴ^����h,�e�6�ԉ��M��fM�	|�"Pw�n��̵`gqߔBQ2n���#t�L"�h�ߦ�{��z�4�j�:�f
�i��ۖ�7`g{���l�/��@�ֽ�X�7	 ���C"s4�٠_;V�˭zm�?��~������@D���ڪ�3�4cO8�Sɽ�uЛB6-Ͳ]��b���1�94�j�9u�@��s@=m���*3dF5�(���@;��}ܵ`}9�V}]ɽ��d�Vh)'b���Sc*��7����3*ƚP�S@�7<:����jcbl�Rk[�;u�{�,Ѿt��بĈHD�c���ʚ�D�ID�)�.�0vD#�ERFGZj���
2)>å�hhSWO)��"蔕�}(B��$�-�!�9HC�k�c/�5!�	t��45HP	G�V������ �o{�	MheP �A�p���7d$6�)`�*�`�HT/8˳k� H������:����O' ��Co�Eڀ�� yhxPz"�@>� 
�	%@I�W�o��׍���n��F�dn73@���Z�l�/��h,�e�I"�AI�|�� �h�w4+k�?fb���i��Y�\�n�������]��m��F�B<�^�X�9wk+���踾 ���_u��<��@�}V��r�Ads�rE$rh�w4+k�/�U���ޱ\nA��d�D�hVנ_>�@;���]��ZTI����4��@�}V�w[4��j������eXt�N
���N\�i���1��D-�o ���X�)�^����jA9��?�<F(:��9�h{������3�  i��۩�]�mp��\�M&�Cq����s@��Jh�נ��Ph�%27��zs2��%2nc����ڰ3��V%f�K!$������S@�ֽ������i/��E��a��˭z���<��@�Қe�M9�����Ǡ_YM�ܯ@���`v{�VQJKm���jQrM��x�n��ql���k#�0�M��B�a|qe���^2��G[��X��s���M��b`Uʫ�c�λ=K���q0��e�5���v�n���Nm앺U��n5��tLԮM�C��W;Q��N�v�;c(kn��'.��n��"���:]�� �����ଥ�w'�f8��Gd$�{I�ؘ�m�t�*e�fd O�����nX�4SSbz��֝h��7M�a�w8�{���m��-��(�7�H)1��29����Jh�נ_YM�ZTI����5ȴ�)�r�^�}e4+r��.V�z�2,qE$4]k�/����aV�{�4�u.!�M&�dq��S@���@�Қ.�����#ILQ�!�z�R�/t���ֽ��h��$C0GU���U��v�}p�XZ�[n�DXݻ\��.����pu��tEP}�;ׅ���2�����w^���=��#�M���T���e]BP@��vf�%4��-�Jh�:�%�ds$NG�}e4u��?f%����*�ߞ��X�p��ƚ��M���6����ǥ���2��\����28��N%�^�M��z���=l�h�涱D�I�^L�������m\�"�c��{gm�Z3�vx�u��A$��#fI ȱ�RC@��]��c���1��Hnc����Fȩ��M2�:�3�x^�J"&N�71�`v~̫؈Q2�d���r:m���kڛ;ׅ��C��%� LHE?O}�������oa�ξ���K���6�l5(�̽,��Ձ�c��TBS��ٛwG�S��5T�7��z���=l�h�S@�����?����g`l�9|[BVt̆}l����>�n�a�5����v���`��i�u�7���>�y3`gz��P�>AW~����~nE��hr����^�M��z���:��A8�#�Z��9zנ_YM�ek@�8�[3d�5����/Z����=�V�7�3����v�@嗃
�a�ɐqǠ}l���wt���ֽ��A6�h7��x6�p�l��Z�zq�!�clxE�\�v.���QBB""IDI$���wt���ֽ�e4�Z��("AőD�h�)�r��@��M�ek@�I�"A#���4^��[)�{����)�v\�jKc��i���>�S@��S�;�SCRJ"r��VWu��'M̍̔�%6h]jzwJh�k�>�S@�s��_�:+���M�j����
{[g�-�I#�E�mE�`<�޶��}����Aݯg�:�e
�b�g���g��vj�
�N�"�����vݞv��Ѥ�K��k�Ʈ{nKkw�(fu��]�KJ��T��s��7���7vGq��h��UZ�0�m�md���{���)�*]��Y6�՞v� ]�dkPc�lnv6�����w{��7#�]յMШYfRd[;ucb�]�;n��dy�;����m��3nk�:0P�m�g�@>���e4V����+fl���$JHh�٠}l��˭��Қ����Fb&7�@��M�Z=��4�l�qQ�a1��%$�.�^��Қ�l�>�S@�g����E�#�;�S@=m���h��z����&j.,�=��c���KcVݪ��@��	�XRy5�g�m���cv��b7 ��h[)�r���)�v\�ԓ�H�jI�}l���ϒL� PF�3���������m���*�ND��' �!�r���)����e4�r�P��G"ȅG�wt��z�4���9u����+f�k$D�I ��h[)�r���)�u�A6Rm��INyMܛQ���۬�ݎz2)YH9�@cW\W,�n�ջs�;N�\���}l��ˮW�wt�g���qQ�.Lk"J4��C@��� ��8�u�@��M垶0PD�d"�8���^�f;-.%�B���I�D'
K��]�o2�d�i/��#���z�4���;�fM��B�����ūt���Z�	�F����h�h�)�����!*�(�Q̍&a'�"�͙ծ�u�բ�qq�ce7��ݽ��M���"Hh�h�)�y[^�����^�bp&<�DDȴ��<��@��M�­��޷�0d��)!�y[^����~���J��?=�?��Sa�#1���9��;�fM����`(��I@�(�]�ݫ �"��S��S-��`wXU�wt���mz��hy�S�U0�i�ӊ���˒&Gv��z��]����ɪɰ�t��'Z"�C@��M������;�Jhi/�Ra������@=m���h�%4��;.Zh��8�ԓ@��M�%4��[f�����G"QC�D��:�S@�酀}���T$������Z��Y%0y2EA�@��M ��h[)�w�;��oǒ��ڀڢp��
����"�$����H�D#cH�!H��,&���V�� ��	� 1c
(R�T����@�B2�"�+
������eV_�%���B! A�
nٲ#f�v�� `B���� ��"B0"F �H!8T��FE����*�T�tK
E�A���H��d�GSM�m��4l)	�XB5�)!	4GdD��-" �5����ꪮ�_�Y2�cVͻ(k�u���ov�k���$u�[�� p�pm�     [N �HI        ��XC��#�������OV����q�ݸ�f��S�ـv�\W��n�93�v뫴��S�q���{tGɴ��\���eS��ݼZ��ŻF�,£�7�ԙ�v�+�vF7�'�N8�ݬnx�p��,`���m�z<�/�Y�xP'��=V����/(SD�(���m�+�=�3��h���at�)m����}���70x55ݹ�;l�c#�UXr�+�c!N� 5�s��X!`Ȧ����m&�nB� �)޶튔5���nunQ���T�D6&�WV�cY�v�������L��l��U�A�g��\sɶ]�(=/l�*�U�Z��
//3�g}��ٔ����m���6㥎�K��H>�v����;u�[$q�4� /�u�&$�mk����)�������*tƻv�vH���i6��u��n���I�5�Cg�r��d��`��Y�[w69�E�hJ�v�F�S�iض�4���7O�ˣƦ�QI��v۷hi�D;�@>c;:���Nq�c��v���Ў{���lzݣ�%S��b��n���"�-���6���Ԓ� �,��Lv����c���k�y�����R��r�a��n�E��M�؝�vp�Ǚ��`�Zu]��q=`�٭����9Պ;7=%��iv�-Y滣zq�����DL�:�T9㊥UZ�]:V���b(W���l����q#�ih9�96�r��r��m�Rrc����T���oS�*mUT���Y1.G�R����F�`�[9�kj�t��j0kN-��.��f���R��Ɔ㌭USd7�&ɫnf&/&O\�%�}\:�!�z�;'�'Q�;q�7mN��^��6K��X�v7m�`�m�pT�CnnM���T^���M�^��9+_My9:G&G(�j�v��t��ww��ww�A �GB�}@v��S �1���U����]_oZ��r$N�i��^��Kl퍅���7����Y��J�ݍ��o]�c3�;MRF仩"K:!m%*�����Lp(��\�Xޅ�t{=�Z1���9��7]�ȩ��:ܸ�zu�'�`Vz���Kd��u�vy��Ku�aW�O��p��a�wm�ͤܖ���H�V��ۭӶ�;<n3�=q'�����vQ�EU=wiBX�bB\l��sm�(��X�q:����Ҝ��g8%Ln2v�f����s�����ڂ��m�������e4���;�S@�x�cX<��Ln'&����ZJh�)��� �����JI$4���;�S@=m���h,���,�H�B(�$4��[f����ZJhi.!I�$����}����G۷� ���`w�xX���o� �+�:���4��S�J�L��%��c�4�n%����p�X��S�9��;�<,��I%
9 wwf��ߢ?8܉5NAC@�IM����>��`s1�{
&Mūm�(s	�$Q4]���٠}l��֒��K��^F���'"�[f����ZJhϪ�>^:���Ȉ1��@��M�%4��h��@���8�n�4�Q�rk]F��.4$���az�𙱤;F��DLq����%4��h��@��M垶0ő)�HӃ����� ��h[)�u���ġ%2f��I4�L���4��;��{����Sl9"m�DC  ȑB�X�`�J:`��c	@����"D�UV��뤦�|�Ze�u!�S�#RM�e4���;�U������jD��' �!�u�����1�� ��ڰ9��w2[�|���h�t�YI��v8Ox)�>��rn�v��l�I�S ŎEI�ɒ(�s�[w4���:�S@�)qVk�`�ɒ$�Z�����hlUhϪ�>��4DD�I��>�S@�b�@�}V��n�{��TLq��������Z�{�9'��z,+�`y�ftS@�gs��%#Y	q����h��h[)�u�U�z�d�<���y�ݭ��j]�V�r�mmѳ�!�ܻ&�^M\a��u�mh��h[)�u�U�wt���h]X��1@Qnf����[ZwJh��h�X�cR$�171���c�����͈Q	L�wmXn�Ɓ{.]��	�$Qj-��4[w4���:ت�>�\U�&<x�ɒ%$4[w4���:ت�;�S@3��3���5
/� �[�����Iz�r�u���7kdk����RT�G�1�a���A`qS��+]6���1)e�M��plČ�8�]��7��t�ԛ�������[#��gR����I��6���t�pݘ��C�۶��I�;���R�u����aE�KZkك��Zc�Mp�y�^K��Q�乵�mzm�̦����m��݈��N���l��}��^��cMd����p1��85V1CӐx)�lۓvv�g,�������rl���!rC��j�;��F�t6��T�M���c���
&Kl�h�����e4�z�Rő)��$�Qh�)�z۹�}l����V�֒���2bp#p�=m��9��;��&�aD)����źr��SSA.FU5`s1�`l(Q�s��-��z۹�vu�0S���ɋ�ٍk�I;dnU�v���w s��k]-�]��!Hӈj���!�u�U�w>�@�����h�˱djL&L��M���I����b��QT��"�c�`}�xX�s�`qa�r�mR�.U4�m�ُ��5%3��~Z�~4�é�0���Hh[)�u�U�wt���e4�Tc�)	�pjG$4�*��ٖ��|~�?��h�mH�Hq%,u;�<N�sFN�s��<����Y�r+	�v��]PLq���)��$�Qh��h�S@������V�֒���8��qh�S@������V��}V��h]X��10Qr�e4��}y> 	�"�m��~��|��M��W#r4�4��9����Қ���>�)�z�.�I�M7.AԹ�>�^�����Ӏ}���;��&�����R��ԍ��֯<:՛���Sj�0Alm��Ak�ݞ3�Zݎ�t��i�T�K�M9���;���9�S@�b�@�t����u1��"n%!�}�S@�b�@�t���e4Ԩ�pR��ԎHhlUh��=l���YM垭"�/�"N5���M��h[)��R��dɍ���ʶ�*�e�p�=l�����[ZwJh����0S�at��-��g��G��N����y���)�.�v�#��P�d�+�ñC@��M�����4[)�{=�
�n(��nb�C@�b�@��M��h[)�z�.ő�0�28�F��;�S@�����h�he;scǏY!����>�S@@��M�0�cF5�D�JC@��M�­��4[)�vO��Ǟ��z&�ɂ1�"b����;ﾪ"���Y�K�&��ZL��'�`2�';�9���*�L��g{N�ݎ8
�p��I@X6�9��q���d7��md��bg��.9dָ�9+���etō��\�sq��8W������+o'mTn���>xnnƹp#��W�c�0Z��Kn�Ŏ��rs����j���a�t]�
R��ڤ4Z�Iy�w�����aJM��	�3�l��A�z�'cAr3��<#ة���;gҚֹ�7a�����$���C��;�S@�����h,�k�I�s	��Җُ����dߡ$�N�T��Ĝ��~�?��h�h�)�vZU�6��L2C@��M�­��4[)�{=��9"Y�����aV��Қ���>��h/�ľQA̎d#��K������: �6M�=�X��<�9�[��m�$Y�&L�1DȾ���t�@��d��r�>�.
�Y!��ُ�
�9�����`w���>��4cXDA�Ĥ4���u�Zs�[)�ΦX�L�⥶��JS��;6ef́������垭�I�s�@�}V��e4���[Z��~��&j/9J��c���t���W�@�x7l���[)[]+m�\a�0�f�(�[)�}m��:ت�;�U�vZU�6��L2C@�۹�u�U�w>�@�����Ƣ�# ۘ�U����\�coޯ}1�� ���R�F!�!����i%�K����5�����'$c5c���#F�G˧H�� w�HF2%��)�t o�;8�UHC�)h� wM $P�.�A�t@��ZR�C��5�Y8 `p�DH$&�E�2��5R�4i(��(H�B~R��H1H���DmhBD$T��F �$Jh�D"Ü+����RȐ�*F�ݛ$��MJq��p�[]$.�;;�U�0[�נ^0d���n���'��(��lY��(���k)	u��J�(D "�,B���a+/ǩ�|�!XR��|�~3�%"��D�	� D|"�Tt��~#�G�; _��O�s�~o���=��r��da2dj �E�w>�@�YM�n��b�@�)ث6FY!n-�e4[w4[Zs�hm�M��㑨��<l3�̽��gۅ��@�ܮX��ۙ((��չ75�2n
C@��s@��U�w;V��u1��K$�jI���V���Z��h��h,��\0��'0q���j�=�S@��s@��U�{�����9�'��q�`}������O" PD(%)H(@`,h�B�E����J�Ƙ�&���=m��=lUh�ՠ{����3�����[ʴ�ũ��y�*5΃D���R{6��s����M�(�p>��k�&7Y�7~��;6{Y�`}�xl(��HwwmX��?h�da2A�j-�ڴv<,�2Ձ�c���S'�LS�[��J(En-��ۚ�������ڴ�é���18���z۹�zت�;��@�[��gS.Lm�K$�jI���V���Z����̵`8�=��*�TR)�uB�{��8�UOkm�����t��q6���]S�Ӛi�/:�v�[��t)��ڝuĔp�63fo�^B0|�l�t/Nm@�	���1�x6����XͶ�ѣ�n�x�v�z�%���n�-4����qY��Ofᰔv�7�"Vۗ����^���J<w[J�;m�#�K�j��q�N��ۓl=�Ic��B�;9z�W�ˊf(�xi�U���N�{tV��v�uk!����0,u떹��ӗ��3��z�ߖ��s@�[��zت�;���"'��4�Z����n��b�@�;V��iV����#Nf��s@��U�{�U�{���=�苍EFA�0#��zت�=Ϫ�=��hu��R����h� Ȃ5��}V��s@����=lUhiw�-�D���#�7�.ͺ�)�H��N��w-7�nN��u�w]���8�9c�3M� ��ڰ9��Vs��DG$;��6ݠ�H�P6**��5rN���rR,QX��"�B	D �2E,��F�lUhy�Z�����eɍ��d��H㙠u�U�{�S@�n��[��|���E�E�s�@�t��z���s@���u��B��!�j8h���>�w4i)�{�S@�x����Pl�!�$qr��ER�خ�]�����$�`�i����ɵ�f7�'�nf��[��[IM��4��h�RPj(�?���f�m%4��/[��}m��;�����R4�Ƥe2��z�3������		�" �@�@0�$�)�P�$!Ȑa�� U6*��=�p䇭%4����@xE����{2Ձ�̵`f`�؄�3/K��g�1�	cdNf���s@���wJh���/���j8�o$j2cS���!�GX�pò��ӓ�M�դ��pg���L�ۘ�I�Ԏ9����;�S@�n���s@�g��.,�$��%������B�S&���ݵ`f`𽈙2pŵ.\���4�.�`no���n�m%4�Jh��Ս1�L?�s4�]��Jh��=�HĈV1�XD*��$#F8��χ \��A����s���Jh�Jh���������#y��rsm�\��t�:ɨ�ն�.���k��ᑷVd�1c�'�h�!"��M���>������>�vT����H�r�)�}�w4i)�{�)�}�F&�b$1��Hhz���Jh�Jh���vZeɍ�S)��m�j�b"'wK���q�`gl������>Y�j�(�A�a8h�Jh�������/\��33����v��of�n���TTu���Lmϧ�A�1ƕj���zݳ�q�{$ļm�۰�8���Z��h��Vv�^�Ʒd5�^���W���������^����z^=��]�9�J�Mؼls��-زT�v��M����ϯ:8����D��x�r9٦F[t/#�ksF�>���}gE�Nغ���^�D��"��2�M��(J-BJm�.��c���z���h��K4�qs��5gGn�pؕ]g��d�Kў�#�]�v������)�}�w4�%4{�4�B�Ƙ�&���hz����M��M���;=IA����s����M��M���>���v\���H�m�%ʦXyB��r��75�}�w4�%4���5�0x"E��z�hz����M��M6��~��N��/S�q�6�$c�X��~�������iDj�ֺM�b�6͐^xձ��H|������M��M���˖�Ә�I�Ԓ9�뒚�#����w������x����1���I(�A�a8h�Jh�������/\��<��T�6L�����IN�ޖ�ݵ`gq<,���@�n�i�bm&O��4�n����zp��wϖ`ܱ�xl�n
�O\��hą80���l��.D�X9�5��ul�-�<ݡ������4{�4�S@���h�r���P�$�A�@��S@�e4�n�m%4���5�1��DH��О���rIߞ�O/�H�G��E�6��M��4��Pi�x�cdR޷s@�,���t��m��˖�cN`�?��G3@�,���t��m��>����୩b�RS���WZ��V��<��L���ۓ��틚5�IG����dp�=��-��޷s@�,���݈V(���Na��m��>����e4{�4e�ucLsi2G!�}�w4r�h�Jh�M��J5��i�"s4r�h�Jh�My���H�E�j������q����Ą�� �! �HqG����4\�D�`(L����{�)�[e4�n�nYM�s[X�C�fp��uk¯m:[��k !�s��
�p���z�u����x9lQ5��~���hz��ܲ��Қ�ò�ҥCb��r�`s��W�"!L��^�{�K3�P�C���*�(n*[n��7V�,�����ǅ�ϳ/4�{�P�451c&%��@��S@�ǅ�ϳ-Xj�S����;9�I�.YRҚhuL�31�`^������V�&������~ U�� ��� U� Uh���@_� U� ��� E�@����A�"�A��@E��@�"�D��A�"��"���DP�"���AA�"�P *T�"��U��D",Q�"�A`*`��E"��A ��  *Q�"��`��(� `* �"�(�`��F(� ",`���"�@�"�A�"�E�"� �"�(�", ��(�",P ��F(� 
��"�",@�"ň*",R(��"Ĉ* ��`��b
�H",B �E ��b
�@�"� �@�"� �F(� �*��� �����  
��~ Ut �� @_� U���� 
�� �*��U����U�ي
�2�˵��0�
�����9�>��|�P
�A@i��RP�RD� @)�!�� x��P   T��(*��(�PP �  @ �( J�P�TA%E*B(H�ER   	IQX    0"�(
@�6 �;�K&���nz�����OR�� >�z�\]�y4�s4��aӀ �Wq����� 8d�vr������=��.>8�z )����C\ZUc�qjG  <
���  T�`�������k�;�{n-Kg�Gqk1=ک��wud��r;kg;� n^̜L;�u�y��` ��k�j���W��|PzUgo!��S��N���k�{�| ��f}u_o'^�����<v^���@@P   ��@�}]������y�w��o��U=swm����G�R���{��콇������[� 9��n-��q�|  ���^�w�m^��lﯶۗ}���:��r���{O}� >y�\w���;�x�f��}��> ��  ��  ր=�W�Oyo���x�� b
  �"��a�h=� � )Jv`R��{�P  J
N��(h�t@�� K1����M�  � ;h" ��@  ���P  	Q� S����4��0 vt}���� ާ���YWw������r�� �m.N�mŧ� 6\ڗmǻ�_< �Vo|�*�e�ˋz^n�4��x Գ�z�^;���+���N i�	7��D@  5O�L�IJ�  �=U*���CL�=��&$�a0 ����j��@  "B�*J��� 3Q�}���7�?������Tn�P�q�0�BJ"��_��]*�"���U�������U�"���QBJ"">���R�?���?ʾ,��O��w
�ȥ�d����6���B����O�e>���8a��*�fs9����.�F�>h})����3�$���5�l3d+��?T�~�4F!�¼O�m�d?!)�к@�1A���,�4@�3F��p������$%1��p�����3N�e5���H�������O�Bie'N��Z|�˾�����gY)Lћ�g)��}��IqMo����Ml�~>e�Le��G�oe�z�_�aI�W������[Y�Azw�)�vh��gƍo�e#T�1��!t��� ��rr��G����T�*}7�_d�f�����#�zvD�o�� B��݆�4P.j�F)���0Ha��C���E:���������r����h�v�d,���`����4���D���ϊ}��vu���}Mx�77��j��>U򴄫�s5��gܦ�#C�!IBf�)�h8F�	��
� n�����+���]}�l����B�3����[��q�m(1�0��-3�����		yM:{O��3^�d�c[�!^4����]�T��>$��
���wmvr��{�][^���J�Ii��;e�=3o�NZ�$*�������k8��]r�e5n�|��_/��:^���Y����R�۫ei��6}���O�����k~iR@��g�_B���8����-��l�va�4�C���N�frɘ~��S&�=�<�~f�F�?�6F1���|�������CHU�:���^�+1�k�>6��$ Ukz�m.#-�m�^���}�j�ǆ�����F���:6q�#s[8�;juR��!E"Q��
�J�6p.�� @��������o|ɼ�����d8��w�ܙ5��}Hԍ%��<Gg��lh����}Uk�<����3ㆾ�J��|q]�|�ĄI� ~J|�ө���C����;��韏�6a~v�^����~^̽JB&@��8i����$@�F�����'�l��F4 0\$4o�h��u�i+\)Ń]g8O��a��$�4�4lH1�ՁU�4�*@)d!��8~�IL�B!MlcrR����*�����Z�lt��Q�~�Ks��~����p���7'ژ�H��Mh�9���O��M�����Q�x�r�,���翵���'�!K'�j;u�K�yb�mjB1[�~[ά�.�\|����ܟ�zuڤ��i�c^�=�w�����h!!�H�N�ӆ�/-��~������S	�!�sy�+�<��!RV�2ג�}��^fV������Sg6��BV��ƥ7�2VdA� ��&�%r�&����7 �� ��J����\3A�l�1+M;�@�!���89��&Ӄ�
��0�͐�it;0as�Ø"U��D2cȵą\x�Xt��cï��{7ٷ��Q����^�W��RBU�"qѠ٣�o��F�������}SA��i���Ɲ���
}�p6S�B��@�ld����8pza���kxk���m&���\������%04D�0;� D Upb��,@�Jm��H	�i�F���
n'S�9f�j[��g������K���W��Uk+t٧�>>H\���E�7�S_a��N�t~O�"S�GƵ4�lћ6]}���W�ԯ<�gR�[�r��Z�yywWy�=�!U��x�^�]��ڻʙ���f�/��3�����me5���e9���~��j]�R�^?R�W���٦�gؒ^fQ��Vq~��%��^ͥ~@�u�BU��3��.���)eu�����^y!x����h����F��~g�cX]�M����U#�>�@`QD�@"D�%C�"�~�TW���RH	 �R!�7�����wy�|$!U�n���x�~T�Ի�i
��k\����w�8��L4lٜ7/39��j�b�����ڽk�RB�Xז&�!L5����W_�n8��?$�@��4f�%��l��!H�	sG8l�{�j����e�"�������f'Y��U��e�/_���ȥE�|�OD�B��\�!����7����j1�S0#��t��!@�����B�.�Xa�3��Hk�����H��6�Wy�!R�T�^=�yjϐ
�v����|!yv��Y��� ?G�f\�Bn��g�����f���g��0��ԩ+�!���������y�Ǜ�#��T���LI!k�S�#!cD�	p��R�:MV����RD$�̄�hm�Cdha5)�p�ӻsd.j�����V��d�-+�&q4�c��f���SG~��n�D%!���l,B!�I
᧌�j��?�M�	�I�u��>�Ydj@���L��	���4d���a�C��!R%�"��g�S0�n�,�aB�P�a}�:i��4[�:2��D0c
9����kA�nd?}�SD��ړ�d�!2p��k
h6K��Xo9a�ҘCGM���O�6f�}.CVK���f~�֓C��B]�!��6K��T撻��j���7!��bYЖor9�����na~+3F�t��QZf�I[]N�|/��ݿ/��c^Hni�G�s{�wF����)���O�o�!�WE~7��>�a;�7�I�HP��M&�0f7�8��_�L$A�> �bDX�U�X��ģ
�p���z?o�kzr�]~ͿF�?	�b�PX�3K���
}��Y���p�G�7�h����N�����W@���D�5�3����ۯ�
/�Q���S�L��0,$FA�,&�,�#)s�8��
2�3�.��/o>o���RLT��{�{�Z��>��5���R��E���-RNO�^O��W�&��g���{����-��R\�)�ц�k��wFg��t�?h�#�z^qz�k�6����w��ԭc�o[�}���!*��;��^�Y�γ)�^�9�ZX��B����x9�����D@(Cl�+����߉O�,,���/�]X��e�I
�ˮh��J�������x��nҴ}J�[v׻o���������9�F��J]jѷ�t)�[to���e�����j�P�0h(`0j����Dh�
4t����E
*����������Ţ�6ŉ"�+���cF�����V�k�5e&/$��~
-�*�J��՘�¯�9rK��	�|�`���CGz������E!��îh�8s��f�d0��n�}�s[�۽D^~>aL4s��SF�H�04�$jh"P1��"�����[�����: �H����%Κǔ�A!N8p��~qx�b@�+�H!������4��������nsA��)�9��8}����BL0՛�
|LtƘMg뛜����$�Z�{֩��|����Ef$*�+X?ufW+	�e<�m7�Y|�ڪX��b1�VS��Wn���}ٍg.�����{�
�c�.�x���\���R���tO��5����F��4l���x�G�]Y���8K~�J�X׳��G�v�oX�c���w�k-y'�R����hϲMt�A�C�"B�,R�D
�&�Q#s#$#&��/9x�4	�����U20�L�		!F$H�Y�� f��M����a]&����!L5�g�������cß�p��4��r8��)Ņ�ہ��Y��f�^l�ڵ�����*T� "PƱh�(q��8�?�46l��O�������CN�=X~d�Z��Xc�=#R\4?��L?H�T��6a�����F��[�k��nJS��_�1��?,
Z�,J�D����	:����`� 1���A�ls0�p4w�u��,��?s�\4s5̰�~8�������k�����o�k�9�/;�r��ˏ�����I�$���A�\4ˎ�������5��6��B��g��Vo./WsB>*���[MrE_����-��������MP�)��8�u��;O4�W��4˦��㟈ˉ������������Xk�ύ��Մ��ٹw�n��������Ӌ��
c�f��8�tq!��۳\#��p6e�d�q�M�Ѧ���$�U�à����
�.�<6�
�
|�%
&	��Lt���绺wt��=�����| H �����J����#�m�����Uj��j�96 �� k9%nIiu���Qz�z�e9�wD�G��8C����`ְu�@���R�e]�jU��Z��iVڥS
���T ��l6�Im�N�`;m���([vض�h	6� q��EF�b�e�Z�6�?�}mm�����[�鳀rY+6��Vۑn�����}o��6� ���}�O��am�m� 	H6��cm����b�#^�ʹ��J        $    -�m�                         �               ��     6��           [@   ��                    >�        �         � ��        �                               �m�D�v�5��J��n��j
�V��b��z�`Gm,�2�����n]	���p�P�܌-����m�4a����⧃'H���N�m���v�pכ���a��[%�\M���t�`+��Ֆ )V��\   8[�ڦ�� ��j���Qm� p   p���� �E-�gj�l v�9$�nb��+�V�U�a얥@gv]��U:�������� ���+�K\�c��V��{>�[����V�[b�l�@YyFG�m�n"7��j���x�e�2p5�g@6�tk�3I$��d�"�o4��,M`�{.~;0�&�ʜ��XQ71(��kd��F��ĵPqUO.L�tvJ���pUm�''1ٓ�S�eBV��`U��K��HI -��mdY��=k]!�Q��X��#PY�99#�ܚ)��uV��-��햬n@�t�ջmA���0lԫ�){<љ�]3`⧶�m��*�d�T���x����6�t�u�USˌ1��K�Mn�PQӲ�jq��	�=<O;7IU�,��ܑ�j9�<"M,u�XJ�q��nn����-���R��[pj1���(�%�6�W���@����(+��,�ښD��N�� =m$gdř0[@I:WpUj��V�Vb�'��D��T�v��u��5*��I,F�3�ڨ
]�wD�]
��F�ڔ��s�m�@6m�&�p׃gQ�8y��#��m��[I��U�����yn�myٶ�H8z^Ļ��m�Kh�P5���ɸ���yᣕ�ۣ���˻����WYӳ=E�s��QBN�S�����ָGc���],�7"��'I]���ͫҜxyeh+v�@P<���Y%��ۢ8��Q�S�� �zU��V�ȑ�Ӗ�Kl������l����E����� �A���i��M�k��di"�[�\Λ����$pkXr�}d�(Ȗ�h�ĉp�ѩ��V��U��RU٬�a�v� [M��    sm�����n��`$    �t��v�nM�r�m�    �[D� �ݶ9�����$�   qt�� � �`	� �Ph ��N[�wIm�[@�� 0 ;v����    �n%��6PZ�
�m�=��޷  ۫�6�7m�sm�[%$��6�@���  ��������H6�      ζN[���  m�� -� �� 9 �H�l�m&�$���2 �]�   @-��`� m& �r6�H� 	���tR���e�k�H   ��H�[M���6���-�m� ��sj��� -�^���m� 8 On���-��[  �i2�d6ݴ�������gU��	        ��l �a X`�      �ٖۀH  �ZmSi4���mI��i
�Ғ����x�v-�m�6������*�T:��J�K!�J��~��phi0 -�ſI�| $���i   �`�my��     /[�6���8�G[n�Rm��l-�  -�Qm�zh�^� @��	Ě%٦�4�:�MΙ$�n�-�I��$������h�^!#��� p-� m�`�-�K(�&� �m�Im�:v�H�6�;Pk�������9^إ��+�v-���m�Ō�B�6zy�Z�7d� O-.�W�j�3�ю�����m=U˰Fl�6X���@Y���_7�9'>6� ��	�7Q2l��ܦ0a�5U��P-f�T@&�%���j¶��8�⪨���ͳ/=T��qUcv)��f��!�cg�<9^�� .�b뫭�y�ڌ�ۡ:�yj��"n���u\݇\�svR�ǧ�|��� Y�G8�$�#x1�v컇`A�=�Q���V���jQ8���X�9m��zŷ$M+�����{d6#8�2\A4IpJT�5�@Y�v��C`Yw#9�Mu���5U�b�C���P�	{^��$.����L��*	��e6��[nz��]+`s�s $ � ]���/Z�k�I�E� U�p9�%�ㅪ뢥��\�ƞ�y�VU������;*Ö�H����nBD�U�"���N��K��Xx�mq��d:R[���+mJ��U*�0PR�Z�!��&A��iV�
��n�bj�H8�8�nղ�!�Ъ��m�\�Z꫃iY��	�t�6   	����Z�6P*ڱ�X%}��B����*�t�m��p  ��ܲ�JU*�UUj�Z ֖� [�ͫ` �  �	�6ǀ��z���]�� 8�t��ѭ�&۰[f�p��^�6�$p6� �t�u�.���@I"FM�`m�k@%ez�i��HMU�P9j�	�R�:*�`-���P(P�ĥ6݀	!v�6Ӧ�kiА ��[@m���m6[v���n�b��u�嶺4-��[Ij��Ž\  UJ�ҭUHK0­DO��#z�떮LB�u�n�lm��  h �hڷg m&n�n"�	Z����v l�]�t�����QV��[�\ ��l�K=�*1Cr���@,T�U�Dv�箂wGUU��u�]� $l��5*ͫjO����
,�2�6e�`۪�j�_g5e%p��`��I����=
�my�p�=�����v	  -����6� an�j���:i[n � @�;����`u���3��77Y4C m� ��9Z*�	:X���M�f6Ͱ�`	�����':ޣ��i��n�PHUU@@a�!��A*�T��Zf��:�K��m�p�{N^�M���^�}�T�p��Itہ^��F�� l�������kjKa7qףci�j���a�%�^�nz�U`1�+]��IfV�u7Y�t[m�Ͷ7!�M��"��Y-�d�Yn9R�\��Rnwbx����$L6�Ӥ^@�
�T6⮟5�T�D����� EC�6L�S�hzl����*���,ns-'��G��xݍRc�l+̩e��Z����Ӧ� kCWt#3m��   ���:M$���Ilp   mn���;�q�]R�;P][�4����r����5lu�Ͷq�>�}�m�|���U*������lb��i yD9�r+�/J��]���.��6���F��Z�HoPI���(�}��С[`ÒIm5�fMȭڛu���%`.�]��^��l��Wf�����ÒH  �6��C�д��m��kJ�qv��6m�m���}�m� �	6�w]ܐ�z�-��l�$ -�۶�m�a6]���kn mm :6�m 8����4Sj�  H      ��[[m�` 6엣[@    ��(8-�m�����η��   m �ۀ8�-��m� ��u\  E�ms[�d��m�V���m[G�	 p  l�ꭶ  ���   ������@   H��mmZ�TN�m d     m���h����; 	��[d9�vӆ 	81:�[%-�I��`� �`����	5�l�����pGU��������[ )����oc��a][�c?'�[v�����4͵vn��$V���t��ѵWfqI����wg��U�Aviº�`-ܚ�fZ��-� r�3�k��^���]���
��VʵF!z�d���HF 4d�x^�UU���٣r�U�:�R��#��:�nn���v�t���z�MFӳ�H������7G�Nն�n����7mڣ�c��u�ֵ�[s5� ���(�� ?��@U� GH������"!��+ �~@~��]�v��q:"�DO�tD0Q(�4��tCd��F,B A�,!�HH��H,B
E�1!#�"��$�� �"d����d���2 E�� D�D�HHH����B!$ @�",���+$"�0`��	H��"�	2H��!V!$X �"@��d�Ha		s� �Ea�Cj$D� �,� BE��EE^� �W���b����Ԅ ��D"� H@�!B�#�!��H���A�� DaB2�"�D� E�ZAa!�S��@�Ej��� "�T> Ҙ�P`�hz��$c?�@�*�j �A���E�NFB1�EB��:? �@b*PS�Dڂ| '�D��E��z�� �x�ڱ�� �����6."� �Az�����@����z: �� �)� J� >��tx�N":�D�@S����A��1Q���	�/� B�`�C���pA k�"`)�:E��~T��A��:�� ��T�F��@օ��_��v	�r"��� �b�뙙��YMf����˓���Hؑ����3����X)��X�n�d�]��7(�Yny%�f�` [I     �6� � �[Cm� �l @Z��      ���-(VsvٵZ�݆ۗ�T��܊Z��P��ܲ5T��٘�![���ϳ���|��s�9�ɤX�FKo�9����r�6��ة��:9���=u���tZ�W-rs��t�G�7On���v��۶6�s{v��ڐ=u��Ѩ`mi�s�;�K�m���'t��*�+�}��t�5��i�|���BPxF��27�C)ā���F�>݈�(�n�!��󖪪C\˪�H�K�+m2H���tu<��R,l7��qb,�V�2�<�� ]����v��2KR�K:'���mL�Gq.�t Vyz�d�H���UU���*�����+t$K[&5�#�zVu��l��m��V�ȹ,^[�Mp�6�NQWeP�7�Cu�t�ޝ����pn8�n��˅��qE�
�rNca7���ն�]�Ƹ�'	�ܼ�-�rŹ-�f��(:��X]����U�n4��q�ezނ�s<o�ڸ.	����2M�[��ʚ'Q()�.٤
e;g�V�ݫv��z�c���0X8<mڤ�xs2��R�[#Zے;u��ģ��J���xe3�`��e�jq[�x��`sr�3Q�KM$K4�KV9#�b]��]sۍE�0LX��66�f@Y�K�I� R0駖'u�N�p�N�����8�\�\�Xe�����Kkt�K���/:�r���=y�nq�0!h��xHK@l��]*M�*(yy��q�sӮ�c��l��Z�7��m�iV�W���j�[H[! ���V����Kd�d ����
{Gb�Z:'P�M[ks�s�kh5��.y�^��!����k��&9�Ͷ��e�355���kS]�T �E6
u(~AOȩ4>���C�ӻ�������ߤk�{���h�G�ת�����y 
����C>xG#zg��V��	��Z�.�N����{+��Aρg��&��pd�@k
*�� Bn*ˤv<�����5�k�n�O�Є���'gݽѤ6^��[�t��t�1Ŷ���2CՀ�{K˘�G��쭼I9
�#�w)�=d��Mgc���9�jfh��k/�)6��f�R�ngo;�`��"/�=�<�`L��	����v<�aCq�Ǯ�)a5H���`�{.J`oa�t�1<��1��ɚ��h{�h�V��λ���bRI�D�DXU�&���A��4��#L=�`�(�'��1�$��)�yF��i�v���6L�u��y�������t�0ޘ���Z�UķcdǑ�Y"o VK�A8�v^���x����w��F����M�pI3@��� �z��j�<��s@��Rx���,i�I�������|�I%��*\t��R4��F���r7�ib�QdrM�j�<i�XzJ!L�������htjA�%�@�廚��hwY�Z�Z��STɉ�I�%�L�$����\���R4��}-]a{㎮�k�s�pY-�e�3Pc��7\���fLѼ��-c�qc���;�cK���F�H�vG�Ȣ�x�Q�I$�-v�˖�h۹��f��z�F(G&0q5W8o �x�ꈈM$��o/ �ڴ/)�y ��N ��&h}��%;��X ����� �M��Ԟ5أ����f�k�h\�s@����Kh7�qD#��	�U�Iz7U�%���뵳��<�����p|`��x#xF�F��#�x�?�Z�-��-�s@;���en��d�#���̦����4�;�cK���MS&'�9&4�93@��� ��%�wkvp�=ŀ�����U�2cs4��4]�@��]�'G�P� D���f����S]]!�QF9$�@��h\빠[n�w�f��eȱC ��m�Sm�oiw�ZWcNwmpҜ��s����X���٫V5"�dn�:�h۹��Y�[e4/)�y"�L�@y$�I`�1�$�0=F�4�11F8)3@;޳@��h��L	$i��聬�FK*���^f0$����I`�1����cc����C@��]����7wx� ���ݳ "m��mM)Ēn6֓_ 6��[@6�`�`����lS��<��v����m6�x��@�m����J��oAhwO5��Ҿ���vez-�\��2�zz�V���a~gYrV�a����=��gї���ӫ��ι]3Wb��7I�%(��c�[R�q6�{u�̾�|�-x5��Gl	O��m]�^7M��qc6V���Y2담3Z$�Z ��9���,�)���U�n3U<s[���tq�Nث(�I��<��+�[01'��&'#�cIc�8�빠�Y�[e4.t��g[b�Ɏ7$��Uk ;�]璄�S&�ޘ��M�w4=�`�(�%c�I4	&A����4�;zc���R)&@q6�yzS@��� �z��)�yyL��#rcN`(ㆁ$�0ޘ��d��`{N�t&��9����0�n�.mFhiy�y��a���]ەz�<�0���N�خ����	&A����`{zWU�ʺ.j��]��ٍ%	w�		EJA���'�j �M��<�w4��4ꔰ#y�RHh^��/[���Y�^����u��Li&�^�s@;޳@�e4/Jh[lM������Xߺ� �Q�sN��� �n����E1�?
$�"@_�v���f;m�<\n=96��GX�[��۷)�ӹ*�D�hJ(�$�h�����M�������;��$��ۆ���fl%2k�ŀ�o }v���j�$�I������w4��4�?~K����=�ύ��I��&
bi�e�`�1�6d� ��Ѧ�����iddI�94��<�(��Ѧ����*R���Eڻ�H��.;�l�<1@��L&��x�TٷN����$�DiE#Ȝ�C@��M�]��ux���|h�WᩑI$ƪ��`N��z�Sl�0=&A�e���H�HɌi��-����h�M�]��m�8(�hJ(�U7f��sLwoL�� �}D H�P�5l�>��]�e]ڻ���m�@��h��h�M�e4��Zc@��<"��%� ou�0�JE����I���\��G��A�<�7 ����4��dfA�$�h��L!�)�'�4l��z�h�M��������ib�n'���-���w4l���H�Pj5$��5$��߿~����0{��ݳaB��^�z�~�jdCrH񤛆�z���)�^���S@����O��������6�3U)-���V� *�t�LCĥ�n]�n�aZ�u���%�]�e�_nݜk�s�uδ�0<�:{n4�i[i!Cn�X88�lg[a��c��T�uݍ���dܝ�{�x�<�O`�n�'D���h��1\�k��--�Pi6HM�Mɑ�v0u�n�8�ݞ8q��g�w͸x�s�8�Aك�Kr�b=d���<\��@#Л��{������i�c{+j�vs��v�v�q
��.�;.6�X��g���"��D��&1�3�<���^��Vנ^�s@��v���2�Mـ>�fyBJd����5������;��$y�ۆ�U�����-���)�[T�<�H���AVU�`l����7v��]� ���KtM�x�Ɠ�I�� ��rST���i�wr�J垎Ɣh�u�=�����v��j�Lk�M�k���f�ΝP��_k'F�e��oϷj�*������ՠwR*�G5�Z�352�5��'o{��"�ň�D�DBU#��,�M� �M��գS"�G�!8���h�V�yڴ
��@2�E$Q8�FɌm��-v��h[^�z���m�8F�hJ(ǎ8��ՠUz�������=E��X	x3!��cBݰֹ�/=&�ȁ�'llz����Jx�~A$���2G�M8�
�W�[n�k�]�@���x��cmL��-�s@��Z�ՠUz�lDL���RYrR��S5dݬv���;��n�����ì�h1�+
J6�V�
$a0*YX�5�C�����ZRwz�i���ef��Y8���!YC{"�� �la0�j�	�$�J+)�7wm�n���}3��)^���Ų�.�����]���p�0���%��.����FB��B��hA�)k��c&�FZ�����	42��,�n��Q�R0�\GI
@dd�$3L&9��Md	Ȓc�����Y�f�����B����֙BW{ C$�K�f�H\�P��1֠\�GI`f�Kk���]\��*R"��j�q"��Ehn)� L�RҼ���X*B?!�@�`��� ҆+��
~A]�R�P�#���'�"�5��>��9��s@���r7�I�%n7�k�h^�@�����h�	E���&	��r-���۹�Z���)�r��)��Ǎ�H�X���"]ڍ���l��2!�����/L�n
�ta�oB��۹�Z���)�fx�����_���#I�H�1�����pݳ r�� m�Y�"d�wr�QEBQ�<qŠ}���@��z��h��@����ܘ��
&�4/���ŀ7]s�JWa
@��	(@! �vP�ww�4=�2����
Ǡ[n��[)�[e4]���Y��~k��j�C=n�{9��gΘ|���������fdc#��z!�"%1��� ����v���BQ���ŀu��ʬ�7Q��qh�M���۹�Z��ޡ(�#ds�jIT�l	$i�%��� ��WQK&D'"X��@�����h�M���u��#I�H�1���u�8�J7w4�:���ŀWP��,b'ʒ��_�g��]��t�h�Bdu�����ۀ�i��1"�]��9�M��t�6ٺ�n���aw4:�w8��n�g�Ӫ^�;ct�W�t��Ks�c�H���1uq��΂N�/��v1��r�<g��^�\�ÐΡ�C�p�a^\�6A%�(���t!��g��vU��z��nݎ�:ً���M�"6�n���P�N�BŲN��bwg����s�{�ھ&A{���rt��uH/2If�-����g���6�;;��%��8�x4�q���|h^�@�n�k�u�8�pm�nW��/[��w���/YM�T�%��0�@�n�޾�@�e4��KtC� <Q�'�4��Z�)�x�W�^�s@���r&&�JTՓW8�`J_V���w޾�@�޿�xтǏ�fcX���/�����WdX�������؝dt�2^E 7RHh+�����;��h���ݍvVL�RH���@�n����1HJJ�(D�J��!(��a�$�)�$�+F�J)�N�5�'�ޘ%��jQ
d�۪������.F6�h��h����^�z�����c�D�"8�ԑh}��/���z��=���z������m���m�@�^�@�n�޾�@�e4����<ɉ,q7�a�R��6F��pa��Ð:u�N;�K�H�t�ȹ2�m����z�w4��Z�)�x�W�Z[�H���i8���w���IDɯoL�׵�>�� ��re��J8��8'�z�h+�音�!$��P����� �i��;��Ww5svw5Wwf��^��w߫�p6!(�{�`����W$�����z�w4��Z�)�x�W��>߿Ǔ�sih��rn�:筱��2c��/\ю�nWk���wSt�P���w���})�:d�L`N�����d���Dq��"�/YM ����w4��[�bG�-���m<�(�p�~�M���z�����<�e�6��y�@�n�m���a�}k���%���R��D6�'�4��Z�)�[f�z����Ě���Z��}�l��=;g��^oa��=���Q����8��gd� �Dq%pN/ ��>4�l�/[��w>�@�(�B8�"���0���B�5������>�fj���U-m�I�����M]��q`����B�׷� }������)�$�	�M��.���ՠm����:�x��{S*��ꤙ��n9�yڴ�l�/[��r�����>�>������%V[�m��A���LI*����;cB9u�$��3��	�[ͣ�8�9@qkk��_�������t3�k&2s�1N����<���&���\h���E;y���zG+�sd���na�D�f��=q�wjg�\��w��˗�d�����=��mZN���d�v���W6��a�ч=��[N�u����Z�A�r�-ˇ�����^�rv�%�+2J�v�:^��Y��������A�F�8���J�<\m���P�]�����女z���uz�j�<�e�6��rM���.���ՠ[f�in�y"Ʀ�f�`��� �M�P�)��ݼo�nh{i�l"Dq%q'�y�8�������%�{Xz�����9qȴ�l�>�����[��/;V�޼�?,HƄ5�d�i�ȍٛGP=�Om�v�݊��Uk���f��c~�9/�,�Q��K����nh���/;V�\�>����u]�j�f���sUV�$���s�� �U4%UUU�BV%T�UT ���� ���, @��` T'��^p��zp�{׀>��6"&G�{S*���&�쪺��]n� q�xyB�EW��ŀl���Hw��.����n�j�b��wo ׻� ����5BS���{��>�<NF����w4I:ok�l���6� ��yU%Hx�nm��S��&�7V���9�y�����y�p*%g���vs|�y���(�]��彬�[� �n�G$5���>��l"�$Bm8��@��{����fca�{׀{}�Xg�u���ޅ�*�f�f�WsU7wX��� ��,1.�J�F~�<�U�=���w1vXL�Q��IWx��������9�u��L�����}�9�dI5�&���uz�(���_ w������;���ui���6��zM��	����s���Ƨ!ޭ��ݶS��~�>|��$JpZ��?[o�~���٠^�s@�}V���Gq�n= ��7䏯�nh���*�^�����L�&7$lh�K�5���;��5)���X��� �njO�ɍ��4>����|����';��r��!"2 �!AL�2}~���/_��a$�Q������5D��o�k�ŀw���WI���dyi5s��wm�X|�S��.l�>ke�mAZv5[����|�PP]��� }�o }o߫�uG$6^�`���l�Q��K$�/[��~�����/v����TD�'���]���P�"m��/;��*�^��^�z����ia&D��jH�>�ߗ�������[Ł��og �A��E��*���n������ �׻��i��z�`��#�DK����� ��L�J�E�H�?4a0�`�p�5�t���g�S�t��.��0މp�0��_�B���0�EIx��qm2f�����jk35ěn�kX�����鈐� h�ßk4��K�\��ԥÆ���,����6���J�	�$5��H�kD(2�8���#M�		u� p!%"�3��8h�y�\���J�!?s��ɛhM��x��:�w!���V�.�d�U�L�h0��f o��dʛ`��l٣nݦ��䟌����5�5��Ĭ�����\"I6����35��u��Z1E�+)�dIu�\���sNn&:k�"�$c@�9�X�
b����LHk4$]h�h���3Z!���Zŋ��Wv��}���M����x�ɔu: ���HE�/�N0�]�.	7#ŵtyLԵ�In(d�z*�i     ���`  ( ���` �  @ �`m      $��0�����ز��ug���p�$�#PNL��Z9�l�[]o;F�:Q9�p�Wu�.����B��vm���J#��A����vؐº�v�m\0@d��#��۳0Eŗ�g�T)����=����������nl=�%N^���NsGNz�M�ɥ�-�':�5�V�FSF{G�`��g��q��3�y�p��=h���x�\2�i�y5�e��pd&�s����v8%ݛ��Zx�j�[ۊH�و�&ݵm#ŸW�j����ѥ�[T�������c�6�n���Lr�NZݗ��^���u��5�-�ﾉ�}Kt0����������UX����*���@��� .%���m��
���cq,@��m.�W`wn�[��K���g��ݓp���&�h:t��̚tӛ/R��M��Ԝ��5v-��u���&�Ć/:b�笝�[�ݶ��8���<5�uv�4W>^��tX��]��6��m�Gb�Ok��*ݽ��gb
��m��̊kv�g:P,�5o�>2?�i$G
]f͜��xl#�m�"X6�&��������i�ǂ��Gk���)�j*���vR�ۑ�v+'Z���$e�u;Y`�6۞\�N����*;cY%M��|��1����E[�]���S����j0�oi9t�f:(�p�����ѝ�n�E���絬@��I�O�ܕOB4��f	8.��gc۹�I6S�x��F���h1�짭��)�z-�H^�R�=h�]\�*	5�<�F��$�$�����:I�H��9�'J�X�t�ș�j�P��` �[���ͭq�m�η�A����$�g[��΍�u�u�����2	�8@[�	�q�7[��Mh�]d�2fю��3>:�O
��\  �iT6�������|([y�_�:��[�44�06��%�#m& ]v�D�ת�-Z��ĻC�6��\xl�^6���pbl;>�!�
s[p)��t=A=v.M��6����e� �kj�k#+-�:xN�7�IM�Ϝ�����j-�p�	T�I�ϗ+�n���އs��:�v�8��v���6;<F��Y'�k��s�N�9��X:
8*��u�\�Z�]jHk4_��D�ɽk.d�&�X�����=�Pv�mŀ��{<��uɸ0�!z����H�t�i��߰���L��L	]%�=S��$$M'�	�y1��Rf�޾�@��Z��z�w4}��6JH�pN-�h+���__���/;��;�J,�&9��M�"�/Y�^�s@�_U�^v���ԍ�
9i`�1�:F��Ҙ�J`�1��?>Yx �Ŧ�n�	��BƠ�t�GH��;/F��M��s����Z\�5f���m�&m��뒘�L`N��w]b�L��#�ԑh��_�ٸ~Ł�hR	"!��!h8���M�x����]s��Q2} �j�n�T�Q%N- ����/[��w���/;V��((̏�64F��/[��w���/;V��^�~��}��dI�y1��Rf�޾�@��Z��4��h{رc�����D�18��3=n59a�s���ʊ�hX��ߓo�^2%$B�pn/ ���Z��4���Q�z��}8��M\���ND�r- ����䏯�nh��h��@�iu#q$����
I�^�sI>��v�~?#�X����(?�,f{�����~���z�d�D��5Uk��J���po�� q��V�X���2m�X�$M�'��"�;���zt�'��0;o�06�:a�^�6S2�G+�r�r�7�(6�8]�H��h;\ЉOx�[�T	0
��`8�� }o߫�v!(䆽�0���1@R8�l�I�^���~����=�^ޘ���
�(���=�6Dɉ�p�>�����SO�?d$��>���5��s�̲�
�j�.�U�W8
BKСBU��<`}�^w��rD���'Av�`/�\��>�h�	��9rHh���<��B�o���7k}8�78���,\ln�&ڣ�S�Ǹzg�l��竎��A���.�۵۬�����
��H�Wx�`�u� �MΨIr@�wf�e��9�`LSrs���2l����v��l�ID���(�Ip��jH����[f�z�hϪ�<A��19�q��8�=	yB�U�{ׁ���02ff{��rf{����������Ϳo%�L���J��I%��߲ݿ/}I/��k5$���<�$��w�}����n1�bmD[��%�m���hZ*�i�{���.��<s�ͥj;Y��1���tk��!N���$�f��ɺsö�{(`
x�^is Ʀ8ON�C��"t۞=���;�3��0j���g�`�i���z`x%��:6���yr�};[;sѝ�b�f�K�g	˞;q���h�2
��J[;���5��t����v������7to'c.գK>�E�%a������1�]7&l�Ϟ�dWt��o�|�������������L̺o(ə��6��%�����_��ۡ�$�￳�(r�pn/<I*��o���6�^����K��I%�:�<I.��8a����M�#5$��|���o13�P������O933���W����~I LB�������y����&fe�{<��˦�VL����v��Y�O�2L����RIwN��J�u��Iym�x�V��Ԓ^q�Z^��:�Q:Mֈ�GC�8�ʝ#�΋O\[�Wgs�����ϟ,%P�=ZjH��$�}�ԒK�l�Ē����<m%l�/<I!�Cq��q���Ͷ�y��\�@S��ov���ݶ�v�眙�t�Q�I$�y$��g������Ɠd�O<I/����Ԓ]Ӫ����!DB�%w����������&f_Gk&j���OiĜI%��O<I*��jS3<m�93>��
����ə����q\��Ԁ����J�u��K����?~���%��n�����$�o���F>{%v7�86�)��v��u�1aV�I�6�=c��$�;kfFݸz�B�;� }~~~^x�V��Ԓ]ݴ�3���֒����RI[��j$���6�NO<I+n�o�fg��w3��㜙��{�FL���|��̯l��&n3n@Ԓ]ݴ�Ē��w�v�<P؃�{�߽�s���{6� }}��}XJ��l�5������Q�W��}FL������3/�02f}�7m���HYo�i���m��l���w�L��F���32��9ə�]��I%�U��@E��⌘���n�+[[�����zPM�Z�.:{��.��]�����v7�Q��$��RK���jI.��y�IW�Y�$����%ifjMᑵRU]MXd�����s�Q	(򈻹�o��������&f_^`f�J��~nuq\�\Ӑ�p�Ē�ߵ��Iym�x�W��jI.��y�IwP�mņ'��6��ԗ��1�����%��t5$�{�O<J��d	 �*��(°#
�FFJJVB2��|��� �_k��7m���[�{X��)�ck$�Ē�wCRIw���Ē���RI//Y�%zd�x!4.�m���^z�e�3svy�GSg��9|�hg\�?a���s&(�4�1&�I^���%_]f��^^�����%��t5$�[��MI��(Ӑ�Ē����f:�g�{|��κ�S�33߻��7��Q�������3,�A�� ����__BJ������{i�%W]ǩ$��8��k�������w��_߿�_�� %����˞�U�3��%PB������I/���sRo��4Ɯ�RI{���$���$���g�$��7I$�~Y�P4�V�Ya!D�`EQ� B UJ0�	iI">�m��{��}��)��9z�6�����8t�6��*bVi�P�S���s��ӎ�띮�vz���BxwY��q:����Ó�'���� *82(��j�T��'�C��À�wݮ�ϛr�w�:�u�^nչŰ���9ݻq��w7�;���v�g��5��w�|��|���s��F�3شv��vݱmMls�{a-�u�'�\ck�Մ9,�;LԂl��c]��n<f���<r��3�e�Ǳ:�>u�5�����'����"���8MHj�k@����$�����ǩ$���<�$�Y�jI/}�W�$�u	�ȱby?)jI��m����s��P��VDM�w����ɻm�����&f\��؅US-��[u6L�x�6��O<I/��pԒ^�:�<I*��=I$����$gYF�LDNCrB��� C��Q7�{��������홻m����s���*��#��o��wm����5+RB6�I�F���J���RI/=�y�I^wqjI/}�W�$��f�X�!���36Ŷ�c�iַ���ɸŶ��[�9pxF��wﻻ����.�KXPn~��}��Ē���Ԓ^�:�<I*��=I%�ō��4�M�I<�$�;����|=V4�$IP%3!pqA��asf*� ��`A1�H!qE�TG.2 d�,����0�
`�Q�Sʿ@�@$ۙ�\�3.wث&ffy�w�~��w�۷z���|����en7m��׿�9m��wfn�򫙗�����m�n-I%���d�G#D����_ߔ/�BW��|�&ffz���&f_i✙���?7ݷ��%o�5�,O'�ےcݶ�����m�� $X��������g���J���RIw�:��1�d�M���]��'�z�I�$���7�m\��jKa����,p\\�i���Ϸ�� ��}��[oo�ٞ�b	/�j�~����������u�kp5q� ����s���H�CZ����ٛ��~�����j���Ԓ]�|�jHF��1�ԑy�UR�5n����&{Ջ'�$R���J�@ �RP��%���x��9���3��)H���@�sY��.́.h��f,��4kZ��I4@��Z-�j�w���8�a���� C"]�5sA֍c.z�)<$��iDH@d �����a��D�(���Z0e�XZ�3��j�̈́�4��˚#���4/�D��i$�*\�&Q�i˘��B�1�,"kH�<����"�߻�u�����*_��fu�05���& �g۟����,>>>pI��S����Lִes�mKL�����������B%0ٴ ����0��їY�%�h�\ Ca �.�������"��� �t�� ��
�?�_��E�8�A"
�������~�wm������� ���{r�Ե��q���{3?}�k���w=��[o����|��(?�Y�������7������)�#b�W׉%z]F�����y�I^�Q�$���<�$�K+lh�A��ı���;�T��|�S��i���h!l̙��50���d��H?�&�&� �'q��_��@�}ݛ�N~�u�Q_�Ā�B+������ ��?�!X+�蚲�ʫ�oF��L`M��v�S��_�>���Ow�O��kT��M��f�� ����	�`n�J`M����wYu-�Fh̤�k[��,�\�{� �o� u��i&�B�!\�УQϻ�krO���ff�7V��j�ݬ﫮p�^P�JIy�_ u�׀?��`��G�Wv�$�nn����{`�=�U�@g���d�tG=���R秧{��=�����>��}XJ�5��J�������i�zt�ލ0;o�0�V�K���j��X��y���IIU{�X�����K�ꋥW%�YUw�w���Ѧod�%����^{�X}[��;i����eJ&���0;{ ��Ѧ��L?|���?y0=�}��@�Q�Ln	�@����<����X{�f�"$�����eT���w����љ��3V��L����c��	i0k�:�L�Kz+M�zWt<�ڶ	&�xn�nlp�-��m��e�s�{u��O'p�qvYٓ�:���]�MӔ��ͻK�T���N��u�#z�}��n���+�nH�۝lg;<�*�V.�PW��]�I�{n�.^-�[���*vG{�n�l�>��-��6����3�^6?;�����>|��:7��������n��a��hc;s͛7a�'�v_j�V+�T{��v�-���+������׽8������G$>���kJ�Ѩ$(ɍ!'�}�=#n��7�q`t��y(���������B��Q7wk ��b��x�+�h޻���bL�
91����%:��`mn� �o����{��,s"$nA6���y]�@؈[��. ��X�^,�u�QR�6{E��8v8�ڬv�ksb��'OX�^qppigh^�=���#���/�O���,��ŀ>���P�$>�ݜX�zے���K����}��ٽ�?�ǂ�p��� ���w훒w�k�`?�Ś�/%����,W1sStMڪ�n���b�9�np�P�&w���������U��7��j��[	%�K��P�}��?o�ذ���}�XsK��7�DLi8�����B^Q����{�W@��~ŀs���K�����j��Nb2�e-�p'=H�v9x�ӈ:�v=;$C��Z����b�`w� ��,���a/
"		G��{�����r]�6�n��� ��,��� }o�z�f���!Dw���{��˷�����9�5-aE����� m�XLDFD$�W��ŀq�� ��ud�,-\�MU�]��$�	F$DB
Ps�����'}�훐����v�˝2�4bS �	�f��?}�vnI�A�@�0H ,R �I%�{�/��׽8m����*U~;��ҋ���8�ypLA�G.=Q��FÌ�hX��G����W-��6�,��� m�Z�IzB�$�
B�HI%���X~eU��3H�rf��;V�m������;��f��"�H�DH�Tn�����S$��d������`ݐ`I#Lu�L[2�gՅ+�MIsZѹ<"*�D`�AE=�x�=�{��s���!!$D%�F"� ���A �33���s@�bL�"$���i�h�� Ԓ�BI.�{����� ��S@��$��hD���14�}r��\���^�:���qփ���jyc�kX�Ѥrbnf��>�@�����O��~�P���>����X}K}ue�Z-]]M�]�SI`{� ��F���O� �T?� Ijw�h�Yr���H�Y���?���$i���#X�vZ�Ys55rMڪ�j�J#�������;�����X;�f���V+��Щ]��]�����5D%�BQ	o���wv�`m��-$�i}?V~�6N��4tRN��ڶN�T�m�UL˙�9������n���N��ݣ`x�x�̰�`{�4;�n�]��{NܥlQ@���79��ݡ^ ���]��)W'�b�^��^]��#3�Zږjݻ�ݺ����[:Ig���<�#��C�BD	��nzܶ�qh���컞9ώݝK�^�m�ܳ�ӳcmrQQ��d�O;3�x�1<�3��8ݎM�[�S��g�u�@�˶�1���y����nwI���1:�2Q���~w�9��0��zK�"!(_Pwk}8����HOɋ�ܓ4;�4��`�u���,�А�!*���\�+��JcQ�!�}�����yϪ�:۹�y�)���@�$rbnf����?D�%o���{��ذw���
����>�On���6�����j���X�%�""";����b�<��4:��Ś��<L�&H��Fv �����[`���jׇW�<�ȼ������a1��rJ�p��L��ϻl�D(��QPo�ذ��1M�MrMڪ���w���L����@"�!B�҅�(��3��`��`����x.�?F<�ǒ4䙠y�Jh}x���BI/�(��{��`��ذ���c�q"G�\��<��0��X�D�ך`=���.&�U��ŉ����F���0:u����^&&�I�x<j&��$Hn��Xx5��Sy�ۗ\�$��s����w��/��.8D71��!�����)�u뛚����^�(�$rbNfϻl�Q
!L�^�X�w��׋ ����Ґq&��4�ss@��ٸjХH�2,�Ie`F0��$#eD�P��)�"D���-KHRP�V@�0�Kh��%YXRUi�*�T%RDD��e��-Z�8��Q�Q
��7�w��]�JC�)���L�<��4�w4=�M�\��<���Lq
Ln	ـu���6"!y	$�����x���b�9�m�]u��T��J�\��q�9@�������p����	����=����؀�p�Ǒ��F��4=�M��6nI��k��� @U #����nh|����LH��lD���ŀs��0��,�vٚ�D/D(@�F(.d���e֦����5ff�i0:~���#Lod:&���ʥJ쩫���Q7f�	B�BI~P(P�	
Q~�ߺ������X�)CQҦ��ٹ$��t֮���waVV�}�f�%
<�B����DDF�������~o޹k|�m�x�r����H7�V�Y;g�j'\�6�Kq�㱱�ۭu�9�����806tM0=ݐ`v���ѦE�d̔���\�Һ�k �{l�IG�Q
Q��ŀwwذ�Zŀs�h�6aV^QY��
��4��ti���/�.�����ύ�x.���y�G7wk�Q�{ŀw^�X;�f�%�?+�}�h���n	����4_ZŀzK��N ��� �z�` �0�� Ad�X\ ��RR\�N0�S����#�L��	�ڙ��76i^C�����F"�)X����d�a%�������F"ap��@�9��$*B͡JS!D"�FF���0C��LB0ep2-4��p�6FOt���޷��S�I���$�;h���ճ�9�p�h��RЇk:5�ͻhe��!��j�6�Ih ඒ     �m�  � �h   ��  � 6� H     ���q���C[i֣��[HR�rU:P-���W=�
�E6�^vK�^0c���rr��/\=n)�v�m�Pq"�K	��Nu��]2]�ix0�(.۫�ś��s]�]W��d6��8�,=;���Yh���봷�����[ѫ�Dg�+׍�Ʊ�֍�m����6r�����x�M�m����g��Ֆ�Zs�c�,�:�r���g��J�A�\��3r�Un�i�c]�EGX�Yd��Չ@7�G��J���j���kg@�-�v���W@��eg�c���y%�{r��F�pTlg��M�8�g,<�vi�٪�ڀW�*�ݕځJ���v�N�3��c�U3΀����
�6���`��5p
�R���\v9C'V
YY[�γ�m���h�G���YqSTEpq���[��Þ$���ć"�-�=��ۖ�m�T�C�cv��S[�C�'m�;U��m�nt�6C�W]��,��6��r<����3��v�7e���l&xN-Y*Yv�lj��CiŖ�snj�ۦ��K�1�Jv᫪7<@�#���^��d��lpUt�E��3uU\K���A��(gG*�Q�0�ǈ	9���[�sқ�.�J����\j�����d^��N�\a؊�˳���ˡ������e+g��C�Q��֧U���6��@�9� �n��^�Z�-K]�t;�W[��=�W��\vm��^쳍v�wnI<n���=�j��.Ͷ�vɌ���5S˲��R����*�N����I��D�ӖK�9+�"nkM�	$�-�v��5��T,�&�tT�bC�	���u�k�0n�^5�.+a�ҙ����t4�p=�ms�������Df��~>V���U�!�C�'���;�UD�����>VS�	���QAä q��� Y�C��\���^�/�����=��*���g;%���g�1��tf�#��7����=g���������v�7!��88<c`�C/��K�69��m�s���$W[�\�6��Ev��M��<V��c��c�#ؘM�pl��d��F�����mm!DHm�W!��S����	m>Cra1�=XM����3#a,�u&Қ;s��'g��5!?&,sCrd��zS@�mŀs�x��J$;�V,�{�54aW�b̻+0`v���ѦΉ�;�fy(��(UA��+��E�wh��L����Ή����{o�Ǿ�&�27P,��6��w�����?o�� ����;�x�w�ֻtK��,���L�<��;�w4wF�:&�&K��
����������h24���c�re�ns��+��:�����tB�UZ1M�U*�&�UY5g�k��`�06H4��vA�����,�*h.�n�������Ɇ�BJD��Qj4��#XP$a�M@5)���ELW�"��o�M0:~���F��U��̢���R���`>�� �z�a��_ws4m�s@�:�d����q�L�=�`v���2�0=�$�$q�$lNf��۹�}��fg���x����{�LoTk.ՂUYUW�S�=��=���v���]q��n/݉�����XHI0L��y�S@��b�>�^-I(\�}�ŀ}:'�u7r$lM�$4m�����oۚ���<�)�uΔK���BO#d�{�L�e}_$%�-	R� I)BdH��>@��	�����"X��D/���^������g ��ŀ}�L7#x��������^��3@����>m��<�"'��ްܪVM����2�310=�%06H4������s@��ʏ�i��m�����uc:Ou�[��:N�F�n^�������FU�-QuyL�07�4��H��B�ηg ��ܫ��UD��E����{�LI`{��0;��$��%	U���+����*�ԓV������_J`wH4��ti�N�2�VXT�ڙ�UV�5DD)�����1`�^,���
!%<m�`O�뻩�DNH��mŠwZnhw]��n���\�����{SEHL�!H*�Z8����n9�Nk`O>9��n9�/�7lt�����wg������	䌙���ۚ�`{��0'H4��H!��.�ev�����?�ś�S#�=�^�@�۹�{���)�0��$���S�A���0=$i��u]��$��E)�����Q-��,��ŀ{m��;�U�v[u�����Ln�b`zH�d�0;��0;�`i~u	4��+���`�,D�	 �l>��v�kZչ!lƜ:װձ�H �m& ����bt�ʹ��{
��3z��tے�b	���=k�8�k;6P��Gi�ݸ�R���I̯��&��At�G�y�{d��bwv�4�f��Cf�ʒ���o;�:j�;������K�j{*�jb��a\3V�\t�ێY�ݰ�m�V�Ӟ_moX����nhw,Zjܷ`U��!H $ RFAbA@{��}|�u\�ob*k[a8��W� k��d7��a�=���;m�D�ON�i�*��T�V�����\��f/ВQ����� �߱�a5$Bx���w>�?D%
dotŀ}���6�`K]Ƥ��ڍŠwZnh[w4�ߒ�ِ��;��H4'�ǐ6��6����,����m��h�����D�&7�h[w4D%	��p�n,��X��J��'c#�K�۳��ۖ��nY�N�6l�.ݙ4�}��@��$�7e��6�Pw�O����A���0=$i���]�1���ar�57$��ٴ��U��RJ�/wq`k�X{�f���#S�sCo$��n�z��6"�2۽0z������YUD��x�����#L��0'E`z[��޸�$��M��;�S ԔBK^���n�,��XT���\��d��>{-��[��x-�I��O���C\j8���T�Ŗ���	�F��4��#L��0;�c*�������Wj�`m��$�<�D$��o�� ���>��`m��6eڣ^xe�`N��wd}�Z��#A�"�B���W
#b�K��f����,�&*˒��*����X��-�� ׺b�8�Ł��DN�w� �Z��͗eZ)MM՘lx�D(����p{���Jh���$����	"�&�,��%������<v��X��v=��ř2s3u\����d��ym��/[��wt��m.���i���q�dhnf���,�(��	U��X��ذ6�h��!H	I���wu��cņ��~��X��X���wSv�e�+UwYW�HF��4��#[�`��A)S�'��g�|^{�_r�6�J6�D��	3@�o�"5��p��6���?�8��ގƛM�j�O(q�p��Gm�t���ʼ��-�(t�l	18-����-�V��x�������rC��ŠwP�W�d��$nI3@�빿g�P���=�zq`��� 7� ��OY'���&���[j��<��h�w4�es$����"M8�`j���w� ����;޼Xm�,�m�ۄcm�9��9���������	k�|�����׋ >��sR_Gkg3��L�JK\�m�	i0�4cp�,qGC�j�C��y�7[����9i`Wy���au2�mzi{g�����Ӫ�%�X%
�{0Aʯ0��<=�!�V��7b�ڮL3����qb��ۛs�vQ�9�v.smу�I�I=�/My3�N���}��d[�+��f3n����=j{;�a�\�uƸ����=�{M�Ud�zM�>(;e.��%
�[q���^�5���z��i��t�	H�L��y�w4m[���s@�۹�x��\�&<��	�ԙ�u�8��""�J���`��� �z�4�ҍ�ҍ�$�Ȧhw]��F��0:IM0=��a�v*�Z��&�`jIOۻŀ|���:��4;���W�d��$rI3@�ti�����L�4��$ʫ�����Tv�w�=�-�v"��0v2vj��m�^ǌ��.?{��x��E�����^f/?~?4����d�0=:4��W2I�$9�$�$��빫����j$��B�%�� ��� �cŚ�Gu�cL����G�9�}�ۚ�F�!`wti�M��b̺*�*fiV�=���]��� �x�,����s@�q�\�&<��	������wF�$i��2t;��m��\��ؚlk�2�7<�.�v��*gV��u�����_?���}_YW����*��|���o��[#L�j���b3����$i��rS�����O��꣺�_f"թ�����`mn������pK~64#�n�1q�
�����0�lJ,	.�e��L�\��p05���n���B�J�s�) 6pџ��]hc"�`L�����Ȼ��m��H� � �7y�
a��`�P(J��e��T����bK�.o.$6@�.�԰$	 Z[$J� � � �?_�C���M�2a�Ѽ@� �VA�3��Ro�5������iBV]�j^	�H�W�?��ѳ����R��1�0�3Q'6��V�B�dB0H��X�%	���4F��7�).�5LI�K�@֍hYBm��(J�:�PZ��S�A\��� D`E���	��S@(G�z�D�� :	�����nh޻����E	x�D!���Ji��Ѧ��0��U����`E���28$��H�N)�w]��n��v���s@����bo�Et��ۨ&1��Y�X�s��s������y�"K����#o$cM�I��Nf��s@�� }�[	.H6� |�V����6H�O�hWj�/r��w]��m��<\gW1Ɏ�	�܋@��x����S=��,���Wm���4($܉��;��h�n��s���� �`�S���q����A6���\ݬ�7� ؄��ݞ�{� �z�`�n�DL�����7s� `x�z�-�֍��K����堶:ώ��<i%���L&Lm�7$�4+�h��0;�4�푦�U���0T���%M\��^,؈�{� }�Šy]�@�W28$��H��&h�`v��?Ē���?S�'����MYt���.��Z�ԔBKД*���L������ti��Ѧ���fdҪ*虥SV�K�Уt{��{훒}߻�rM�:�
@�R���~}�����iZ�\X���8Iml�� ��RzB�<v����"[A��=U���/<n7�WN����+'-ڎ.MP�2�������9ޡ04��Y�m���p�Ν����y�9���w�5�{f��;�ιp���s�wX�Fy�\A�:zZ��a��w=p�zmg�v<�q�����m��1KB�1��ۍ�˳ �R�y�3Z�.��\��v��A7���I5;h�4r��Ӭ�D@�����=�M���\r�6�������p;���f�[?�;�wߺ�`}x���N��u9��x�B�MȜ��빠{z�h��X}��<�D��z����me���L�?4��ܔ���4����@�u~�"&6��I���V��e��>���%=׼XgT�.l�,/QFVe0$�07z4��Ѧ��V���
�4�hCX��M�%�y�K��i�
8��=M�⁥x���ś��;�Lj4�$$HQI�����=�w4=�����%����X��Z�����������ѹ'��ݛ��� B,Q� ��4�>���4}�s@<�n�RG����f�MZ�>��0μXy(���w3@�_�4W�̏#��n�@�Ti��#L�4�ݙ��SE��\��\���>��X�DB�O�������r�`n�LԄ�J�f5���pM���ջ^�v9���;9:��]]���l����]�/Sw�������`|�n^/�D.Hw������1v�KUUE�]]��>��3�7vw��ۚ����qu"���i;0ܼX�7�p�"P�%*.Df���4-��l�"F�D��
��`z!)�w4�;����v�����;ޖcL�6�N5'!�y�w4�v���ŀ}�`��#�ݮ+�N�� h�l[�n;a�Wz"�<u��1��9�G�y���7�����/�<��`y��o�����Ji��2wF�\.��B8I &��4-�s@��)�y�w4}���g䏾�>R(���&����������L�`I*4���a����M���4���D%
{��XI�����;���ܝ_��&��1¢��V� ���(�0%SJ5�5P��|"��~��@��}���Cm�ܒL�=�������p�oL��,��TJrE��hQ�i|kԜ۠Hc��e�٘g��G��#1,n"G1	<�D�f�mWs@��l�>m��P�!����:�oUZ�1 ��!5&h�e7���H��s@����ڮ��ߒ/X�&4�M1dd�0=݋�URJ�0;�g�wݪq7wJ�U�3T����D���X���07fA��F�
u�xe�e�aYx^b`I*4�ݙ�07dkrLP6�"B2}>��R�F�m)���L����
S�H]J��S��&�g�i�����^zTo\u\��%�k�>���햕�r��|@/m����3c)���5�zu��3�7R	v�����;ch{�؈�EG�R:Skm�ۗ�nSg������L��_e;c�ZgG-us���ι5�6��\rv��ivyk��N�Ǌޅ�6��뮱�%�K�Ƒ2���2l�.:�lm�8��mt���/9n,K���:j�����wG7̳hÁMĤ����n���h�������ő�	��#L�`N�`ñ�:�1eb�������L�`N�g��|��ES~��{�iӒ��UM��K����N����;ݽ0�x��ws@�-�9��H$$HMI���M�;��\��ŀ6���9�׊����Lnk[c8퍀D��pu{9��{i�S�)�����.���Wg=H�͝��6�����vF�J�07fA�v����+S�V\�34nI��{�zz
hx�5G8f��,[�0�x���n����rAG&h�w4}������m��-Δn<��"I�����D���`��X�7� mͳ ���]*YfQV�3�`n��IQ���0�T�J>�EV��t]�Kn����.�.�c�h�V��=�'\]��\ܴP����F4Ӊ�$��{��^,�#���{���zK�����fff&��Lِ`l���۹���}��ds		Nw��ܓ�{ݛ�N� P�v���P�*E�H~'Z�!�		���H7a
�R,��BD$�%�B�(�ۿ{�}7� �,��"n'F�!�{m��=���ڮ��S@;�n�R(<o"�UV������z}��{o��o��Z�I��%HR.mJ$���qq���gv��̼�;i5�G�z8���p�ù��8��	���}��s@��4m���w4s��$�Ȓn%&h�ٛ	D���ŀn�ŀ6���B�7���#H&8	Ȥ4��4z�h�w4zS@��W�M�Ӊ��ݬ��Xn^,��0;ȈQ���~�4W+�9ҙ"X���[*4���΍0:ti�)t�U�v9rm�=��[7R�c\*v���f��>�mG�v�Z�i5�$�ıU�N�IӲ�`t��N��{�`䑷���=�w7�ؑ~�nh}Wۚ^����������!7�;X_^,��Ň�L�w��{� �L��E$D�	9������U���O�?�`t��E2�j�,YUWyU��; ��ѦN�0$�ݛ�	�ԀB������Sr�p�'�V?�a!'6L2L��#i@�BH|pᎉ��F0+
ѴajFmHؒ)���m�c4���	X2T�*J���leA�eYHR��c?T)�"!c�6$�A�$$�QJ���$�BA��D��T��� �� ~���tY.�BD%BXF1d#5�������	�(J��"@�Z�(ĂA�m�� �R!��"�JFX��,�߻֒W����) Т�8�t<竑���I���ꮃ���],`❍�y�J�ڔ^&y3L���l�� p,s     [A��  ( �m� �   � H     ��N�C�tѵYw4Й�׉L-�]%B�3�����jT�ev���獸�>��[\][uT�u�6�����S�.Ƅ㴅���Wl�C*Q�^5�GZ얀9�I��u�G.::��@]���Zf�z���v�ۨ� ��6�M5mՍ6�'z��$tے�f����[B<���g�FCi��<��[�����92�
�Ke��q�&� 8�7dr��Q����b�#��:�����Y_l�v�^Z�V��m�j}U�{hB�t Y�Vx��(ݠ�<�է���i�Anv�6�`pؠH+t��v�G.��[@D��0���������{e��gf�6��R�\Y5�gv�T�nED�u��F���m�qB,U�#�.���������fݨ#���.؞N�K���5�veH�n`��OE��p�m�b��ny���u[l�l�kq��s�z'���˶�����U*Ӌ�x��k�������N�G"�d�n/=��u�m�94�,��s�wF��ݥ�^������{I#�Jv���OLeUwi��Mt�0�����l�O�G�퉪V�g��Q�����=9.���ŕX1�2�Z�e�6�}vr
�fI���>���aP՘M
��[@:�L%�6�m�l:�٠c�q!�]�;���AIʓ�97Y<v)T�����n2.�]л��g����J�W�g��XO>:���컇Ql�v�g�4f����g��]�krK��zQ5R�#���mQ���(�&^�3Rl9�rLd�"K!:#tKM��$��6C 5U���f�4����M�1�ʑ���d�H��H�����eS���{s^� �/�&�¸��)���E� & �5�"�w{������agљSR�uz��c�X`$m��������g[m�v��c���� 7���v�΃�x�s���lr4�+�m�t���'�	ڧfN�u�Ievl�R,"��������nrat�F��I�n�bu�kg\�l2�W��C������J���Y�G;t�7n1bٓ���r�m����A��e��-��I�$z;�F��ۙ�nSZ˧-� 5򂆾�}q�?��i�]�=C���x�{zIC��������}8LN'k���k�b�+0�7di�ӣL	:�_�K��ύ��>��Gli�܎L�:���$�0:vA���O�$���_����6���$���s@�Қ~�K��nh����n�s�"�$ԙ�t�gF�:4���4���y$m��Ƥ4o]��]���ŀu�ـz!&��ܓ3T��.�ݫn�u�<P簷m͊[�[x���l{G:;oK5g���%�⧕!�n�m���w͆�/��g�G$;�q`t[�t\ݗeݓ7wWk o��ebBDBBB�&!�	 ��1�2�* �!FB B0�D-B,B! HBP�PU I	;	DD���)�ـs�X_^,�Q2}�}>���2$�I��/�|hލ0:ti�'Ti���X]Q��*�+0`l���F�uF�|�J�w�@���~�ƓƜm�$��\X�F���]�|��`zڲ^��m�ݳ���Ǘ�c�Zk�6��h�X�c�gZ����B�*�I�`t�gF�:4��](ɒ2(�MI�^�߿g�����_�ۚ����t��Hۍ�
U7f��ŀu��ê�$�DJV ���FX Ԉ�Y��nh����w�<i��M�Nf��
'��� �s����
=
����W���5���JH���Ws@��`l���*>T|��o~���m��n���k��wGg���:����3�[i�6�^m'M�y�뮁 n�r%�bX�����r%�bX�{���Kı>�}�cȖ%�b{޾��\!I
HRB}zAjʙ�*�j˽M�"X�%����NC�Q�DȖ'���iȖ%�b_�ND�,K�{~�ND�,K��'�!���0�5���kFӑ,K�����"X�%��z��ӑ,�dL���o�m9ı,N�p�r%�bX�����kZ֮e�5�K�h�r%�bX����m9ı,N���m9ı,O��p�r%�`i8��� �;��M�"X�%���	��5�5f�um˭ND�,K�{~�ND�,K�#�������Kı;���ND�,K����"X�%����2\�[�!�*�nn�3[;L9��:�>��A�h;Z;3[e�,��������{��7���p�r%�bX�{���Kı=�_p�r%�bX�����r%�bX��w3�ֵ�̷̚0��ND�,K�w�6��bX�'���ND�,K�{~�ND�,K�{�6��bX�{���ߟ�Zb�T�|�}oq���X����m9ı,N���m9ı,O��p�r%�bX�{���Kı=���kԆ�&�˫sFӑ,K���ߦӑ,K�����"X�%����ND�,������~6�!I
HRB׾Aj�f�	�.��\�bX�'���m9ı,O��p�r%�bX����m9ı,N���m9ı,MބI
2��`ƃFRH���B0�i*�F!U�J(w=��Y�Z�5.a5���[v�����N�T�m+�US2�nuPv ��n´��;�����.<{m����n��9��|�[s��I��cL����X�nӔ��&�B��m{ck;83�������'k�';ou��ōǴGm��	]�bG��'����)t��{Gvr�˹;X�]����g����9��m ��<���<��w��t��Sv���\�ۃ�{�,kl��ghx�ɚ�nwW���iC��1�m����ֳZ>Nı,K�����"X�%��z��ӑ,K���ߦӑ,K�����"X�%��:{=f��j\�F�iu�ND�,K����"X�%�߽�M�"X�%����ND�,K�{�6���Q*dK���n��M\��r�Fӑ,K�����6��bX�'���6��bX�'���m9ı,O{��6��bX�'��ϟ��z%e�=��=�[�oq���}�o�iȖ%�b}�{�ӑ,K���}�iȖ%�bw�ߦӑ,KǏϿ���3�¢�������{��7���p�r%�bX����m9ı,N����r%�bX�{���r%�bY������덶�.�3u�7]��vX�@�lۜw]N��ջ�^;q�B�g��75Q��5u�kZ6��bX�'���ND�,K���6��bX�'���6��bX�'���m9ı,Oxץ�a�&���.��ND�,K���6��:��B2�H���!aZ�"�!H�'�3[����8�D�K�����r%�bX����6��bX�'���ND�,K�z�����VV]ِ�B�������m9ı,O��p�r%�bX����m9ı,N����r%�bX��Ş�5u4f�3Z���r%�bX�{���r%�bX����m9ı,N����r%�bX�����Kı?gOg�ֵ�L�h֭.f�ӑ,K�����iȖ%�bw�ߦӑ,K�ｿM�"X�%����M�"X�%��?>m�yɌ��Ձx��y���s���WP��n4mQ=��������ۚ��t&��ٚѴ�Kı;�o�iȖ%�bw�ߦӑ,K���ߦӑ,K�����iȖ%�b~�w�C.���fk50˭M�"X�%���~�ND�,K���6��bX�'�=�ND�,K���6��bX�'��ny��e���̹��jm9ı,N����r%�bX����m9�Ή��I)�A(EZEZ�R3ł � JD��9�9���iȖ%�b~�w��Kı:������3u�U6�����{���w�%D/i�}��B������x�\!I
bX����Kı;�o�iȖ%�b{��/���MMչu.kiȖ%�bw�ߦӑ,K��}�M�"X�%��{~�ND�,Kݞ�6��b]�7�������3������m�q�����!��r�����6����y�׵�v�%�e֧�Kı=���M�"X�%��{~�ND�,Kݞ�6�~��,K�����ND�,K��,��&���������jm9ı,N����r!%�Jb�!{Oz�`������H�>���n'�K����Y�ֵ.�Z���ND�,Kݞ�6��bX�'}��m9ı,N����r%�bX����iȖ%�b~��p�F�k&���[3Z�r%�bX�����Kı;�o�iȖ%�bw���"X��?���"&�D�O��ND�,K�~�?m�t�6y+|�}oq���;�o�iȖ%�bw���"X�%���{�ӑ,K�ｿM�"X�%?e��do#�I�$��ǆ,3ɋmB[:��v��U��7�ۀ���xa�M�X�p��M�"X�%��{�6��bX�'�=�ND�,K���6��bX�'{��m9ı,N��kV��.�f��ֵ�h�r%�bX����m9ı,N����r%�bX����Kı=�{�ӑ,K���6{3Z5��ՓW&�֍�"X�%��{~�ND�,K���6��bX�'��p�r%�bX����m9ı,O}�I�RY��d֤�����r%�bX����Kı=���ӑ,K��g��iȖ%�b{�ߦӑ,K���/�$�ֵ3	sY��u���Kı=���ӑ,K��g��iȖ%�b{�ߦӑ,K��u�]�"X�%�什���ݽ�{l�]ˢJPR�:@��h�,H�<����l����]&�ȉ� �\�5)�Pw]v��E��r���##�˵]A2\�� ��������c����G�[�I�:7nS͎q�{X����8�4�ْ�o��6�}qf�</\˖�g�q���Y2v΄,����Or�vͭ��9-fn"x���w������Levh!�'��r��[Z^���;���r�.Y�EnX�V�@j������{��7���p�r%�bX��w��Kı;�{�iȖ%�b{���"X�%�����u�-՚�u5��֍�"X�%��w~�ND�,K��{6��bX�'��p�r%�bX����m9ı,O����p]U��%o���7���{����iȖ%�b{���"X�%���{�ӑ,K����M�"X�%�}�{���6ybUz)�����{��7�{���Kı=��p�r%�bX��w��Kı;���iȖ%�g������A]713]�������D�g��iȖ%�b{�ߦӑ,K��w�ͧ"X�%��w�6��bX����ߚ`�HL1�fc�moF�<.1s�+I���6�骏9zj��Af�MK�ND�,K���6��bX�'s��m9ı,O{���Kı=��p�r%�bX�������E�ɭ�u���Kı;���i�mMpC�<(�D���{�6��bX�'�O{�ӑ,K����M�"�Os���~�q�}m��{,��~{��X�%�����ND�,Kݞ��"X�%��w~�ND�,K��{6���{��7������Ĕ�Hf���%�bX���m9ı,O{���r%�bX�Ͻ��r%�bX����i����$/���7j�.�l��.�d�bX�'���m9ı,?��w��6��X�%������iȖ%�b{����\!I
HRB�I�}��jBH&ɻ	ڵ�����m
78y�v��J��Ʋ<[����p�tPA7jOǻ�=�{��Y������m9ı,O{���Kı=��p�r%�bX�����Kı?���|͞]J/K?=�[�oq���{���"X�%�����ӑ,K����M�"X�%����ͧ"
eL��{�_�߿։���&��{�����%�����ND�,K���6��c�z
�<&�\ J9��*e�F�q��o����m&�� ��a�j$H��Z��sI5��afk|� p�� @B������L�W	�����D�q�1�@dd@r4�b��d�!	b��7�2HF�JL�m�ɡ1	&����Q�9�@�@��o4n.bT�1b���s���Ljg���� �$A FHP�~�]hӪ����!!���W �@�d!	@����FF� v.�N�_�M �A�N��`��b+��A(�Q6/G��w��R�D����t.�<n'"fw�siȖ%�b{���"X�%��l�kZ5I�[f�˩�Ѵ�Kı=�o�iȖ%�bw>��iȖ%�b{���"X�%�����ӑ,K��{�8h��Y5��e֦ӑ,K��}�fӑ,K����ND�,Kݝ��"X�%��{~�ND�,K�C=��;�����:��-�x3�P9���䰺��>�t�_i{1#a��8��U��Y]}{�D�,K����iȖ%�bw����Kı=�o�iȖ%�b~�뷾����{���?}���#�)���,K��g}�iȖ%�b{�ߦӑ,K���{�iȖ%�b{�ߦӑ,K������4L&�jk-�֍�"X�%��{~�ND�,K�u�]�"X�%��{~�ND�,K���;��{��7�������n�UZ��Z�ND�,K�u�]�"X�%��{~�ND�,K����"X�~V�'��zm9ı,O����5���5�˙f�WiȖ%�b{�ߦӑ,K��#�O~6��X�%�������Kı?w^��r%�bX��{2v��&ڻv4��CX��=����8�q�wA����8]��T3�M6����bX�'{;�ND�,K���6��bX�'��޻ND�,K���6�!I
HRB}k�ݫ�]��rT�uk�,K����M�!����,O�����Kı?����6��bX�'{;�ND�,K���[�]d�5�Z�ND�,K�u�]�"X�%��{~�ND�,K����"X�%��{~�ND�,K��}xCZѫ�fk3&��v��bX�'���m9ı,N�w�6��bX�'���m9ı,O�׽v��bX�'���x���I���Yl���r%�bX���m9ı,O{���r%�bX���z�9ı,O{���r%�bX��BL�?_�Y�q8��S�n�UR�� ��� Z�	ۢ:�s�5�6�Aە��8�y�[�]��")�Oe����9�eW�f�Ӹ��f�������0Bi;&�L<Sɤz8`�<]�
��������q��;L��'&�֡۹�ۢ�7�c�v֍<Mn�fn�^���jn@�F�]�*۫�m�z�ے�mf0��v�u�ݑ-��n�JM\֌��-�S2� 8'�5�Xx ݎ\�j�a{�gP���m��)�]ɗm���{!zl�sSI�:���ؖ%�b}���M�"X�%�����ӑ,K����M�"X�%�����ӑ,K����-�.�kZ�ֵ0˭M�"X�%�����ӑ,K����M�"X�%�����ӑ,K����ND�,K�}۞n��]j�̳Y���Kı=�o�iȖ%�bw����Kı=�o�iȖ%�b~w�9�)!I
HN�Ol������Ssy�f�ӑ,K��g}�iȖ%�b{�ߦӑ,K���{�iȖ%�b{�ߦӑ,K���6{5��֭�Ve��h�r%�bX�����Kı?w^��r%�bX�����Kı;��p�r%�bX�ӽ0��r�����ڵ���.Ţ�� �t786�z�i�>�6*Y#��`���J�=�[�oq��'��޻ND�,K���6��bX�'{;���"X�'�����"X�%������Rk��fM]j�9ı,O{���0�mC��o蟢X��w�6��bX�'���6��bX�'��޻ND���,O���Y��3D���fkFӑ,K�����m9ı,O{���r%���"dO�����Kı?����m9ı,O߽���1��k���w�w���o�n�'���?�ӑ,K������ND�,K���m9ı,N�w�6��bX������qV�<��=�[�oq�X���z�9ı,O{���Kı;��p�r%�bX�����K�؏��>��	&�	#0�2$d�g��Xf�m�5��vV�zo*%&'���t���љ�5��ND�,K���m9ı,N�w�6��bX�'���m9ı,O�׽v��bX�'s�ﵫuu��\�uu��h�r%�bX���m9�H�L�b{��iȖ%�b}�]�"X�%����6�����L�b{�6f��T��۫2�k4m9ı,O�p�r%�bX���z�9�H	�" yDb�D4r'"o^��"X�%��Ӿ��Kı=��N%�%�MasYsFӑ,K?� dO�����Kı?����iȖ%�bt�}�iȖ%���L������ӑ,K$'�#��+�	�j�ꋛ��\!I
D�=�{�ӑ,K�����ӑ,K��}�ND�,K���]�"X��$/D%��z.iT��J�W`+cgv�:�.� P<=X6s���SX8��K�mv[�35&h�55n]h�~�bX�'�{��ӑ,K��}�ND�,K���]��
O�2%�b{���ӑ,K�˫���ʹSwk!p�$)!I��p�r���,O����v��bX�'����m9ı,N��m9ĳ�ow������j���������,O�׽v��bX�'��p�r%�bX�;�p�r%�bX���iȖ%�b~��3�.��]e�s2k5v��bX�'��p�r%�bX�;�p�r%�bX���iȖ%�����k���������ow������&a��kFӑ,K�����ӑ,K��}�ND�,K���]�"X�%����6��bX�'�z���I5Lɣd� �G��5��Z�;��&y;!p��������ſ���a�ִML�%��)�f�'�%�b{���ӑ,K���{�iȖ%�b{���"X�%�ӽ��"X�%��w�p�-�.���˚6��bX�'�k޻ND�,K���m9ı,N��m9ı,Ow���Kı���ߧ�n�E��G�w���oq����m9ı,N��m9ı,Ow���Kı?{^��r%�bX������fk&h�55n]h�r%�bX�;�p�r%�bX���iȖ%�b~����K�� ,ȟ����m9$)!I�^�.�WtJ-U�ܩ����%�bX���iȖ%�b~����Kı=�{�ӑ,K�����ӛ�oq���~?g~~����YLj��j��%�#m&T��e��`�q���;~F��nv���뢞L\x�#-�R�;%I����������.�f6ev�vz�9��Ϊ��8u7V^΁:�S��{QNpA�d���u7@�ȷm]�vʖi�㮮�;cg'h����Hx�[���t\u�:���]��v$�.���Kv0T�΍�]��흎���=���.�.�V��f�w8�QVN�c�J�ۤꌈU��:��5lBZ�Z֮�)�4q?D�,K��]�"X�%����6��bX�'N��6��bX�'��p�r%�bX�����l��ˬ�.fMf�ӑ,K����ND�,K�{�ND�,K���m9ı,O�׽v��bX�'s�ﵫuu��\�uu�ִm9ı,N��m9ı,O{���Kı?{^��r%�bX����iȖ%�bw�=�֤��Y-ՙMk4m9ı,O{���Kı?{^��r%�bX����iȖ%�bt�}�iȖ%�b{���4K���&�����iȖ%�b~����Kı=�{�ӑ,K�����ӑ,K����ND�,K�k�Ҧ��ً��v���/-�:�Në�f�ϛ*R;�9��IY�q��v���.�6��bX�'��p�r%�bX�;�p�r%�bX����iȖ%�b~�����{��7�����߯�YH�fѴ�Kı:w���"W�F018/�:<D�����m9ı,O}���9ı,O{���Kı?x��u�T�dњ��]kFӑ,K����m9ı,O�׽v��c�!�2'�����"X�%������Kı?g��Iur�]kY3%2涜�bX�'�k޻ND�,K���m9ı,N��m9ı,O{��ӑ,K����g�d֦SY�.Y���r%�bX����iȖ%�bt�}�iȖ%�b{��6��bX�'�k޻N��$)!w�����TYVTڻ�-k��I���:_�N��V1��ێ:�=�1��"f+5]�������ow�~~~�vӑ,K����m9ı,O�׽vB�H�����A;�M�kRMf�K���ִlI�;��I���bX���z�9ı,O{���KĒM�B�
HRB����ꤛU�35�5��Kı?{^��r%�bX����iȖ:�$���E�D"�B��t�Ȝ��{�ӑ,K�����"X�%�����!�՗Y���d�֮ӑ,K����ND�,K�{�ND�,K���m9İ?�dO����v��bX��o�?�@�&+��w�w���d�:w���Kı=�{�ӑ,K���{�iȖ%�b{�{�ӑ,K�����~v����Ny�*���lBZ�zM���ÍN��B�ڞeS�����;n�mu�Fj�u�ND�,K��m9ı,O�׽v��bX�'���m9ı,N�w�6��bX�'s�����5n��MkS��iȖ%�b~���Kı=���iȖ%�bw����Kı>�}�iȖ%�b~��3ͲkS.�h��5��ND�,K�{�6��bX�'{;�ND��!�2'���iȖ%�b}�]�"X�%������mT�ȒU�=�[�oq���~~N��ӑ,K�����"X�%�����ӑ,KH�h����W��ud.��$)!n���wb.�J*�[��h�r%�bX�����Kı?w^��r%�bX�����Kı;��p�r%�bX��w�,��)�:�v^|q����֔���H�H�H�[m�����;�ڶҘ��[�{�����x�?w^��r%�bX�����Kı;��p�r%�bX�����Kı;�ׄ5���\��d�֮ӑ,K�����"X�%�����ӑ,K�����"X�%�����ӑ,K���=�.��[�-֋n]h�r%�bX���m9ı,O}�p�r%�bX���z�9ı,O}�p�r%�bX��{ܸf�V\�f��֍�"X�%���ND�,K����ӑ,K�����"X��2'����߻�{��7�������؍F��c�ݴ�Kı?}�z�9ı,O}�p�r%�bX��o�m9ı,O}�p�r%�bX����?��6)�$X`a0 鐮."�e4�4\��V���%��c)`apJ�D�V�!l��TƔkhP�H�*�D �cUR�V��сJR���F�`ˀk BB!(�+,g4A)�,�#��u
Hi�`Dd�ȁ��0�IH�"@�d	$�HBB0b�@"F$`H�$H�E�$��jB2�ė�T48~�hj9
Hb@%�0�1�%B�Rd!D��P�D�XA���l$�&`S�cH�"�@�0�Q#`FYe%!l*B���iV�ߟ?U��p֏Y�gvmX5���:�7[ld�L�y��y��s���iӶ���F�A�C,��7KUUV�a&     ��6�  ��>�_��>�` m� ��� �     S��Ō]��֤r�t&���;q[��e5m��}��\�T����,n��N�ύ��Nmi玫k	�zO[*�F�p���R��Tݧr�-v������]ps
p���y�8h6$e�=\�ӎԛ��ە6�T\a��n��\K���z;�:��װ>)���q�ՙ�˸ӹ�{�d�g�y��y���q�2�������{�d��5��B�Wm�m�G^�M� v�Z��ƪ�(��9~e1��mN�U*�+m�M�ͻ=�ARq5� �U52���֪ן$�-T��]��ζ*ZW�0cg�;� 4�pގ��1<�Uui
�Ժ6������Ĳ#�<�v�;P�٭�����Id��-v��m�F�l�b
]�@��*p����f��y:K!�Ō�<�c���&���{[P����l\�7gk)#�a닛�/nS-�/;�6�q�/����;O]�"�qg��]e;'�Ǯ��ezǒ�dYQ��΍�U�r�U�|s��BGYM�Hm�'�f� 9VĘn�\�nH;b݂� ps�]��\�ڝ;&�s���v`;>���T�n4Oc#�����{��n�G 2nwinlڜ񌁻���m�����t�M��;7F:��6�n6ӝ�IƱ�P�^+":�qmmn���&���MV�pg��X[��i]r���Z��{s�S�������N[W#���q�x�g�v��s���B�rA��.�=
�ˮvJ�l]s&RP�#m��f���H)R�l��]��8�x�+�) E����@�*ѵ�Uȳ�� �*�M����pv�k��7#��{As۫�YZ���I��`��;��u��uƍY��hɬ��D8"�@�P���@x�QN�F�
|����7���%����x��3U)-u[R�� UT�j���;��t턍�2��츇U��Ѷ��`�:31�׫qg3&(����Õ�������6-�\Ř ϶][�M7]�6�+ܻ�����n��k.#���pn��ݰf�N%�y�4�<�ΎӧOa6��mpn�!��o^ݮ�۞�/!�cv`P�ګR���� e� :7\�����;+�iAN�O )��3�$��V\ԓYF�68��oQ�mr����+;[�u��v����ڮ&B쩲�*����/��$)!}��ND�,K����"X�%���ND�,K�u�]�"X�%��z'��SV���.n���B�
HRB�g}�iȖ%�b{���ӑ,K���{�iȖ%�b{���ӑ,K����=�֡.�Bfn���iȖ%�b{���ӑ,K���{�iȖ%�b{���ӑ,K��g}�iȖ%�b����ꤺ*�W7V�RB�����ͧ"X�%���ND�,Kݝ��"X�%���ND�,K��}xCY�)��Z�Ժ�m9ı,O}�p�r%�bX�#�������Kı?���ND�,K����ND�,K���a����3.�j��]SooN���ٲ�m�lQ�l�JjW9砹�����0X[�ܺѴ�Kı=��p�r%�bX�����Kı;�{ٰ�PP��dK��￸m9ı,O�{��55ME�֮��֍�"X�%���NCa��,N���m9ı,Ow���Kı=��p�r'�S"������܊�˻��UZ�\!I
D�=���ͧ"X�%���ND�,Kݝ��"X�%���ND�)
H_v�.ʛ.�h�������K�w�6��bX�'�;�ND�,K�w�6��bX�'s�{6��c���������anF�U�=�[�d�,Ovw�6��bX�'��m9ı,N���m9ı,O}�p�r%!I
HS����P!H�hR])��q7n��j�Sy2rr[B�����n sM'y�oc30�u5�ND�,K�w�6��bX�'s�{6��bX�'��m9ı,Ovw�6��bX�'���椚̳Y3XK���ND�,K����ND�,K�{�6��bX�'�;�ND�,K��m9���,O{��ׄ5����u��K�fӑ,K������"X�%���{�ӑ,y���!��(�
�����b�rX�@�!)H�AH�l�ND���ND�,K��}�ND�,K�t�x��5n�����h�r%�bX����m9ı,Ow���Kı;���iȖ%�b{�{�ӑ,K���'��dѣ4ff�rٚѴ�Kı=���ӑ,K��B>׿��i�%�bX������Kı=��p�r%�bX�{��񱽋��km�n����G�)�<m��J��7��}S���m:���3R^�;iȖ%�bw;�fӑ,K�����"X�%���{�ӑ,K��{�,�����$.���Ҩ.®n�h��fӑ,K�����"X�%���{�ӑ,K��{�ND�,K��{6��bX�'�z��r�˚ֵn��h�r%�bX����m9ı,Ow���Kı;���iȖ%�b{�{�ӑ,K��ݻ=��2�-�e��h�r%�bX��}�iȖ%�bw;�fӑ,K�����"X����`�U�I��5���Y�)!I
HM�,.j��*�WuX������?t��b��ލ0���s��GcBf�7;'^�`{J+lM\�WF����(��ΥlV�Eۦ��J\*��di��i�;�L��l�]�%$Ɯ�&��˖�h�4�����#L	��Y��̲�Uv�޼Xg�u��J!L�wq`��}��r����Ƥ4�h]��di��i�;�L�U-�D8��z���ۖ�h�4���-���:?��Y��/�yMU��j]tu�
S�H �(U4��*�x�ewY6>���nz�m�؀9���a�����n�w�gW�m��s�ۗ 7lf�h[\�vm���l�u �x��ם�nFM�  u���mPi�[ka�g\#�+���9l���,�v��q�V�d'gk�{0�#�;�i�vg��r`�ny9��l��ms�佭*X���9�F�&M�mۥ���u��;w/&'���w����-4�;��W3�#5�����;�w �׋ ����B\���ۚ}TϜs�O&$�8�ɚ�#��X�w�M��͆X\�dc��nf�˭z���ۖ�h��hu­���Fԍ�H�	�4�ؤi�;�L?}�J����\���J���U5h���Xo����p�����`Wz�R �m�=���-���Z�v��.�]@(e۳>��o_��LxI#&Ls�X���]���Sl�0=�07�2��̚�e֥2��>�>���D� ����M��4���`N��v�eȢRc�-�n���w4�31/��s@�ߖ�س�d"y1�EeVf&����0;��0&�ց��2���ڈM���^빠w_J`M�����T:ժR���eں6��t���5�D1��]m=L�u�]<g���btF�q8�Z[�m��߿��7�LEѦލ07�%4*�UK.�2�*�)�7�LEѦލ0;��o��ϟѡ�I2)'�����;������T�Q�B
!BX%
.�����X�C˺-b��3,��f&ލ0;o�0&�k@��]� ���$#�H,��w��aB�����j{� }�ŀj�{�ߛ������OG&�7&˫!�]��n�q��)'#[ç�cy�IpGhrXz#2�I�$^�}���λ�z���Y�p$��NL�<��SwF��Ҙdi��Պ^^}V�����f&�0:���&��˝w4��)����7s4>��K�{�� �]x�>K�N!%
,�w4z�V�X��(��q��w05׋ }�ŀv~�R��ع�S���l�۝������msq�H=]�
!Td�r��kF��I��L`Jכֿ���z4��ޖ��Ѧ��c�1FI�	3@����=^�z������hyz�$jHG$q����ޖ������wF�鉪'���$ܒ=�n����h�w4W�^��,��8�$�&��wF�[���4���������Maz��En�UA���	i0j�w����g�q�0YK͎��k;��]qۛ���he-�᫷!�4��т9이L�̝2���wI�Enp�1���N7]]��b�Cv�4�4a4����؍�[����r�q�#�������n�e*�m�γܴZ�<�-�6[�o"��2�ۣ.�u��p>�{mrm��]v�\�t�B��}���|��v�ˮx��:��7�N/[76�&���j�
�w��ק�����m�����Z��������0=8�0;��S#m�1@nF�h�z��׋ ���`��Y�Q#z��S*��f]�W�����LN#L�`z���W�]�	"�Bn9�����F�[��:4���X�����+��푦���΍h^.怳���7�M�I��#Ύ��gwfc�拠B��g�B��qe�6Wh�j�I ��Ʊ�3�=]T���4;��|���/Y�Q<���dM�#�>}x��%
���*���ŀs���=^�zbζ@�bC��rf���4�푦���΍0=:�K�Ϧ�Y3@U՗kb!(R��ŀvz���w4/s@�i�dm�����x�[���4���4��#L����l��b���lx��U]l�];�3����ҏ��k��Bi��{%�͓�I-Y���Ѧ���l�0:���5{����,��$㙠ys��}��V���0'DD�+/.���)fb`M��V��m����E�!|}#
EP��]�? i�2虭$)��������p �P N~�e�B� l���Y@�#a!c`X������A��
D�����F�@�D"BA�������&�2l��)a��4�		.$����j$�a)�1��ba�S	�|�U�����c�� A0$@�#A����f���7ɚ����~( 2 h���)P���C$�$��$���M��?�g�`V r��
!��*?iЇ�P���"��O��*lU6(��|;����nI��������$��)�����^�{�LEѦ�`{f+�]��UyY�Uw��l	�`z.�0&���z��mǸ�!��r
8�Ɋa�7�O^u�ՀTۭmuQ�����8,1��q�Z���^feU�&���l�0:���/u��<��V�A��&�$��_li�ս-�;�LEѦ�X��10nD�h����w4.u��/��h�­��D�%����4��]`M��	��H�|$$���	�*�:)�虏3?g��[�נr��cC�H�G�����]`M��V���0?{�￿ϝ�o�1����^,n��G7A�[`����e���<ʧd�g��[:�U�9�樒Uݮ�{� ���X���DB��e�s@3�~�)"s$�H�4�h[��z4��]`M�����F��M|6H�qH�nI��_�4.u��/�w4^�z ��H���$J��ti�7�L��l	�`z�Zq�JLI���&h޻�/z[oF���L���NeK��u�꓅�gF`m[Kh�d���u�#����ۋF� �ra�y[�����\���E��-�_]���#���T5l1\�����I��cv�����K�)����L9���N;��3�6�=��n�C;;�"/�I��Y�����O9Оqv�Lfh�]$��%��M�;�����۾j-t܁��vX���dm�`(͵�#[�u������C8M�<;�����lc>끍:xm˶Ռ��q^��=�E�w2'M52&	�������޻����oF������t��̺³-�7�LEѦލ0:���<^�v<O��bN9��:�hލ0:���&�i�:"'��Yyu�vQK3oF�[��z4��]h^��I�#���$�h���	�`z.�0&�i������aG�@���ܼn�U��#��ܜvv�'t{G7q�v�R�<��9�N$��G�_z�hU׋ u��	rA�^� �;�vwXfjY3V�nIΟwf�A��PI �Ab� �@v�-_W��'8�k��ލ0=:�V�b��ǒL�/�w4^�z}�}���߲���^-58�&�10o2��z[oF���L	�`{�
�yX�dj
G�_m��<�Ѧ�0:���7��T�]"���:.}��yh|�9�L��o5����J�g�:��E�7#C��c�1'�˝w4�`�1�6F����>�°�(����;�L��0&���tk@2�\�9y�ưNf�w�f�������	A�FB��	! �$��F�$���#B��B	�M'�����n�`n�i���Y�Yu�'$�h�w4/s@��sC����]��r��0�(7$��ӈ�wF��L`M���t���M�ڻx�]�8nTz�9x�&ܻ��>f�� ni�����RW�f��0N�� ��	�4���4��H�9i�1��9��f���fbG��� �S�X�x�aL�z��ST�jT�dk"�h_�Ɓ�λ��w4��4Wev4�Ԃ#�I�˝w0��`~��$H���� b�� D�.B�! �XD ��t]{Y�M�;�x��f�7��$��^�s@;޳@�e4lQ�΍fZ��Ⱜ©� ���a�v�x�X˻�ܱ�L7��\q��m<ȇUt��r&���� �޳@�e4=�w4��hu�����8�rI&�:dأL	�4�7zc�&L$���7�n]�����f�z�h^S+QD"Lj �-`jP�u��`z���l�9�Ox�Rp���1�N
L�}�4� ���`N��*I	IS��v����4�%�
S���r�m�@��/i���1[gZr�9{=;H0ɳ����i:�pӦ%��;(%K�h�+��ҐĻ�����s ��ys���c8�!�Ѽ�c���ݩ0nŶ�� Y�$\�r�(zN�i��9-�t��/\��sۿ�����/�
%F�Ev^D���N��[k��Z��N��� іݳ�X�5��?����o{���q��GcBf�%����]l�k\ծ����3g�S�]�t4V�;E��'�:*��}~~ߣ�i�:F��L`oY.e��u�Q��U^flQ��`�1�z�h��I��PhDy&hH� ��	&A��4�qA�9Qcnf��g��w_����O��n]��w4:��d�<#QL��� ���`I#Lw�04ߟ��;`�pfC�J�nz�g^w/W=�0���y�O��u�ˊn�=dLD�,�Uw��i�$�0ޘ��d^S+QS�9&I���n���/�"Gs�u���>i��/�N���,iĤ� �޳@�dأL	:4��]���+$��swx�%;�4�>�ŀ7׋ =���;�WcO$�NHhz�ŀn��. u����0)��5���s˶�}��c��D�Zw��N�N�3�{g��!zl�v���ͣz�����Lw�0$��i�)�eU��G"j,i��{��-�Mιw4z�hu�'��0xF��I�7�fδ�`B]��!D BK�
��Ed��, �z� �C�ݪ��G$�4:���-빠�Y�[Қ������F8�d��IѦ��vA��4��R_wἝ���`�}h�i�
ǯV{kclz�nzx�����t��"�X�bn����	; ��E`IѦ����D�Dk$rh����\���w4��4������G ���(�N�0�����v]&LNG1$�I��w4��6I����ɯ���㘬CKu�k �h0!��HHF~G����!���%$��G"1�3@=�@��4:���-빠y�Ҵ4��&��(8:�S��Z8�L҂�j��B����yRP'�܉�2L
(�#�h����\���w4��4Pu�cREU��Y�s�<Y�!B�7wq`[����5%
�>ݛZR�sr���&����7wq`���np6<X�n���7��XӉI�%�~��?�XG�T(���,��+�E�$ܗR�n� n���(_j{��ݵd��?}��?�_���@U`���舀��DW�A_�" *�� *��ʂ�@W��DW�TDW�Ȉ
��Z���@Uꈀ���"��TDW�Ȉ
��� *�����@U�1AY&SYBG�e ��_�rYg��?�������`n_|S��$ .Ҷ绾    ���$�|�>�� {3ڕ*f׭u��P�t������R�����@���օ�(��Y]i��B�h�44McE(Z���tQ��5�Nb�r��D�(�F�ιF�tQ�{�Tfb�F�{:)I�iN�ފy��F�,�Jtջ��3e����;h4;�j��4u<�i���j��y(�DJ*�%H�	M I*�#0& &� �Og��%J�	�&M��d�i��`�0��j���S@4`&� ���4̪A%S� h�  d   �L*zl�B���i�	�h�HB��d�L�5C��M=#�bMH�����M��@�W���Is��Щ�iEDA����?����+�PP+^����>�����,wX��aY����OG����v��hߗ>L��1��Y���BA<l7�I	9m�z���h8��t��ݛE@�R��(Y��GT}�m%vZ�pR�ů�t� ��E !DQ$ ��_�,<ρ���d���m�r�!D~�,^<~#���#��/Ǐ�x��<xǇ�/<x���x���x^��x^<9�x����x^<x�Ǉ��ǉ���x�����x����G��x^��ǈ������Ǐ<x�Ǐ�x���Ǐ<x�<x���xsǇ�/��/Ǐ�x���x��</Ǉ�����/����/Ǉ���x^9+�rNNJ99(v@Q@�@E��i���ǉ!(���&}����(0�k6�����gTww�$9�%�vb	uL?��Jq������͊���DaHs"!L�՘�Ӗ�8�r_��bs�����P����_���"5�A�l�K�L�"������J%$i!,JX������ۉ���Z��0a\M��F��kM���	��h�|*�Ȓ�X@	�e���T\sc�6J�[I��[SK	�M8ʙ��(���c�'3*��&���I2dՉ�p�nY=Ԉ��g�(.0t(�up'��;	��Kc^>�V��F]Kᆉ����q�<2xNU�iH��ɕýI��X@�e�Ď͗��xR	�OZA�4c�գY�:�zk�Q\Ʉ�PX�A����񌻸���1]K���q2�Y<H�ĔX@��)3�|� g��W�c(�Qu319��KԌ��~Wg"��dcQ���RH�0j$���S*�hY�RB��i%,Ȅ"����^��X�K�� f�xd:��dp�e�䰇�k84��q=jn�	�Κ�ʖz��e��ضXL\�D$aB��|T�߅ٽmr��}L�2Dkf�xiv"b1<3���<K��03Pд�gdѵ�3Z6f���0�+&��Ed�b�)d��jSjBd̙��$�N�1J��4�r�z7ific4p�S���J6�鱳f4��f�q��nYHB �ċ�$�-"��IY=/'S��-�l%'w9���(E����l)m�SZ7:T�h�� ad����:�C�dЍl�G����mP�y	�;	����I"%*�nF�n�"iC�A�qÜIb$�4��`�4�Q���I ���F�"�,�Ic�@Ye���4��Ag!a!�0���M44��$���@�8��(��4�C�Qaă�qd�aC�q��P�",��w�@�FV�Y5��I��+�u��mK+��i[sS�����	�'rዐ�D(��#D@��IGe��>4߻���n������v�׷�}�9�i��?��_;_��E|(s	��^nfffd    �             �    hj                                    ��r                                                                             9@                                                               /��$7H�@	     �&'��7�7��N�4$bp����p�I�n�Skf� PP�p�-P���H�.��u$/���.BFm݁��L��ŀe.F�l�ٶ 	�,T�ͫk0��B�2�\g���f�
���,�m� m��A�UP;)n���"�Ēd�ْI,�@7@  [d��n��	�U]����YlK�QT�L��ʹb)$[d�mH$�BH�M0c�,k�U�R�-U�퐵�m��y��V0X�����mW�;f�s���eҶ��U@@T�S6T��l��F;qCk ����Kb��U�4��R��1+�ʠ�ms�le�&�W������nX�kK@ �m�%(�Z�D]F�(  ��2cR�K�kl8nt
�(�!i�R�378z��U\Y�@ ��RmWjI�m]Z���sm�˨D˶�k�[��U]�eU��kA\J��f.�i�����Jj f;.���I�ݝ,�m�
�9rk)���sL�f�@�����12Fh٘+����/��ͷ%�]���Tm��J�)\�T�f��5m��e���.��H8�W+HqA�U��V�V�@$�HIIZ�kp� ��H��aCz��<�7srM�I�7I��(#"Z����,���h�FUܑ
�e�vڋ����^M�h�D�,(�
�@�tJI$��$�%�1OoN�:�[u�,��߸@S��������:�U�������D��OT�=�ow��7��tH*
=�/���o�w�?������������ǯ:
<���H�R��4'
�c[ �HjʅZ�~4�ʸC��Kd�-�k�b��q���ة�B����"�(���4HH'�q�(!�(ݛ�bw'�ț z��m��+�D��P�@@��y��)��ݵ���en��.Tx��0���i8�d[!�$/\"oZ��%f�)�S��@0��Z�#��\Hj�23Q�N[N9�ȑ�h-�.�.��f1����7�qc���5��B@��-Qm�A�Fr!Q��I��\.v$J�I	�hӭ��4l�n���-���U�����<�ٹ�k���m��   $�      m               ��            �,�
��՗��A�8����B�[�$F�4^+���� bv�����ŵ�z4��K�ې�VQ����q5��-�i�evf�MZYU�.!�ݬ^6�k�1P���e��m �nV�E˩���R
�f�b��ٙB��X�8{�|���<��Ƀz��p�"� �c\�J�}[O _��g�<�_$�w����  � &5�ܖ�-M�r\�An�ns��bU�[�0�\ {�#:f;� %�.1n���������Y�d����Xddn�s�dg��;�/os������J���k�.��n�ި��!@���}蛭�>���w�<�ޮ��fs�?_�H.���-����<���w�y�{>��w�\.fk7 �M��:wnb��8�a�}9����ɪ۹�KJ�9���z'�'z��&ى�ik�KG�q$Ja��9��6\�k�{�⺪ffffKim����;�����ԽN��s�^��:����󨛤\\gWD�NG#H��I�[l�      �n3n�$�͙���Qֹ̬і�α�v��n�t��<|UZ��a�W��+z%Y~	ͨ;Ֆ�E;�+��P���9�����g[��3��.{��2��(@<D�Nv�T����V��Xsfd�"�
�f��ޜ��OD�W��蛈y�Le>��a��g4@x�y [uwJ�$�^�w<������=��ɂ;n.:�D�fI4P��>����y����Ul��i�*D�������
r�*�{ִ�'v�Ӕ�GSݬ��8�޽�;��ٞ���XI�2p�Y���Y�u��+��y�J����3/ݷ�>��1���rz�f72�Ч��3���T?D��������     �0ٵ��8\7F�����.%WcZ͌����x�*2���n���o=u̙��q�9����>c�(�G���ɷ��������y��������d����y��=>��rd�$H|����R�U�-��R�c3�{Ֆ�"Ws`Au�����&I�<L�qDD���OTW'�������{�;0�����3��Z>�:!.a�
�@�+�n�X��a��K�\t�3Si����IŵQ"d8�2��UJ�2VVK!�6�KuVq��͝�L�9�|�D�Np�L`m	8@�̈́+:���P
�!���������Y59n׽^�8�w�#3���;�;����i���/
v������y/G������w2eN�g��p���r	)��[�g��;��}u�θ����? nnJ�f�H�>C��N��{��˞�oޯ�wv�>�٤eU�"~�����Ѻx����6c;�ϒF��      1�Jɺ���ŵ�3,���p]vG�] �a��?���3��&g� l+]�)�x�w渟M~�g���Sθ~�+>x��w����%��5��}�3�+Z��s���e�Y,\�����g}g��?o�rB��xω�N1���37�kҸ�鯜_V[�#8��:���?&{�����<�w���%n\�2��ނ�?�۟}�'�>>���ߢo<i�Ft�A�A�=��\O��w��0\׫�6n&h��>��陙�w����O1$���ӧ�K�Ֆ��M=P��g��|)��J��:�s����vQC����{����}�����t �f�MV�bbv�M�ߧ��/jz=����������a����;g����Jη'���>���=��Ͷ�     -�17��_3ns��m��m�
չ�Е,4��qln�g�p�y��y�6��&^"��;�~\���e�2������F����D��2������������ʓ%E�f����;�;�v�w�i���A�����<3[ȉ[��Yn�4��d������ÜŞ�����;����>��� ٔ��Y=�<�k���5�O��;���ʃ\��ڞ�D�i�����c��1��9_>�
p��꩷�kK����k��~̙�����&P����J��|fؘ6���zvL+o����xO���}��?==�ӿ(mb�3!����{�W�޻�g���=��77u��lC�wy���݁y=~�S�hڭ�R�[:n�zr��1�2B���;���?�0��.���;0o�������8!EH4/�J$$�KU2�8v���%����B-5'��)�K��H��%�+�W�.3[�����(�q5u4�VJd�k"f�hճ5�i��MFD$9"��r	 �� ��L$��^���/K-���7�<]�ڪ�� �@                                 ��0,�aVL�Յ�&�&��R,�Lh0jfTC6y�E�a�?�¹<�k�P	K�z�n�ض%����L�4��5h݂�k��h;��yz���6�l��gcA�b��GR髴ٖ�[52�{`�����F�p�m��e�3R�b��[��͠�i?Z��]N�;D��W4	2�r&D����?f<����w����=Pª��    
�j��`X�ۦu�yw�u�vl��\�v��2�����G�Ҡ���%6G�g�����y���M9N���h˝�h�W���7oλ�g>���\����y�ίY������T��3�Tʢ�\��]��������aKQ��S@�d��n�s̷}>󿽄���N'}1�u�݋������~�����s�����RČ�9̶��s�\���1���~��#��\�F��mU}o�X�"E�D��D����ߵ|߆���~r�|��Ͽ^���&�����333)�H�%'��wx�w�vY,��#ﲬN�vc��8��#3���ٞڂtn���5�bt*d��7�8�:/HYx�_���9���{��~����3332�bb^$�S/
|u��1v�{�.(�v���e30}���|�x�4�j;ӈf��{���z�}�j�0Ň�k~ט��D@ �Ð   U��֍!�6�3m�z�ֺ���E�R �f�ܳt���	����,;��c>��N�6�_���`4��7���ѻ����܉�Ц�0�2CSM7�~��\|���l+]�^���s�Ra�:r����wۿ[�TgO�(��7��N�l����6�8l��y�<z����U�C���Q�%����.�ʈ�UW�sߜfq��}��3�c����e�Z�ӄ�4��јb����z��c�Q5���>w�����I�y�����Q��ѧ����<E9TLw�Ӧ����/�2Fl��"x۝�(�/��v�P�y}�	�	�G,� f�	���B��Yۮ�~��ֱ[UuO8�2��9͞.Q����q���YW��7�W|�F�|�^cK}�d�z:vLw^���v��n�񺀎a&+%�_e���     UUb��NU��T��-YZ:�(��V�]�&�e���#��6�j����W�k�1g�9|b���hF���f4�2
���t)��m��{���';��a0y��{���*w��s3>��t T7e��_ *f��(ܭ���?��;ќ316a�*h,\%�+��D����c�f;����蜂�ܸ�s�6�y���{�q�{�����ۚ�mK$w��ᅬL�Uo�d�k�N��KՖ�'j���&�&c�?x�������b�ti����d�335�f�b�&ML�d�J�\V6ri���i$�9��a �$�D�z�1���S9ѝ5q�]V�����4vf�����,w��,���{�;�s��۟���e�F�v�cL�ԩ�r�
��#1%'FU��9b�e�����Ͼ{�(� ]�B�;.E��W�
h���b��1��&�1ـl�U�6]�G�.��t�{���]t �Vm���W2u�n��sT�7=�ᷟ&�C[��`���w�SM��/s�$~�:�&J0C�i��E�d���h��eA��hO�=��^�%�B���a�UP     "�	v�a��63:�s�竒�0�,% Q4�Eқ ��..p�!M�<�{�K���_�{�ĺ}Ц�Z0���<z��ku��:�n��G�?��&����X$t4N\��g�t��!��j�K�$�zfeT��en�K=�;��V|لf9�^�nMuN�A�f�Q�DS��a5�5`���h�s�#���L�,������y�6~�w�4�Cx3���x�ɗ�?{� ����1�2�#U��n�BX�G�]�54N�$`�W������9�DVˌ�Ls�#SG��"�a�v�S���nB�D�~ٻ���i~����K�~*��(�$�,%��水eA�0��|��k݈fX�FӖ��`r�=������,�8���/�˘kƢ�V����8���,/ۚ�r�QB�q�n\�'? �[��Y%��&g��w��;�-Tc��M��28���^�q�E��8פe_�eQ���njlEtǢa���j-1ų)��j�(      J؄�7vы�� U��[N�a�l5)+��@&)�ܱ�*��rf��ߎ�"���A���E;n���G��c��4��`��^S��H���B53a��S<{<����!��Mv�z�fffWM���͚��~}Г��~y~fڽ�Mb�_S��`<�S�H����ǵ�L|#��G����3h��)�\���Mdc����nF˶떛�3��ʫr�X�b|��|����ǚ{�}�ZE��1�*\#�������F��GN`�N	�$`�9@��=�
�Z�Rm5ϱ�&��&�M1���D�g�N��ee�K�W.ny�η;�?Cbo��w�9�F#S\�9�3�0l�W9(����ն�GͣtX�w'�R� 戻c�`��G˰�xn݃�?���9�������m#nJ�ގS����jl�>څ�C�F��3+M��jl��D�b5e=���l�3���g���p��-Hnvͮ�SF��ãP⶷�s[ �϶5<#:��&L�2@��H�a��aeAf
�X��Ht�I�$UaUsr��)L��  �                                   �3l�2n��EF�Y`�-��e��k[)�a�e�Hj���X����ړhM�z�Xia�s��ꐽ���+�fS��k֕q��-�f�WJf�3U�Mk6��@�^��,5�lLvYqKKskf&�Q6�b��^�U�Ьq*V�\�3�Ҧ+\��|ہS���3��(zw�O���9�$�m��UUUT    ��r�^2���k-îuI\�5Z�-��͹-���V�L��QS�6�&�h���=�:z54˛�ׯ��@�W�;���^P*M��;�����t5��f\e��!�K��L�f��}?x �f�D�G�o<����m�_�Z�v/誦�x����"��g"h5��F�~�)�Zх��ܾ�/���❻��X��6�F&"\��H+��33332�(y�0�3h�rSb<�M�m�w�V�#S\���w��Ⰱ�	�(�,B$th��N��Tf0��؛q|�9K)��-F���2ۮ]�vY�����U[-��S~��|<٩��oB��I�0֭R�k��^���D��
�s�ם�\�؊��A�ff8|֏^�w���H��o?S���g���UV4"�ء�8s�5��	�wI17����G&�}Z����D�f9i��w�!M�������-���6똚[��f� �n��S      +�c ԅ���4�((�9�LS1�)u�J�;��'�Ӽg���UUkP�*������/ߘs�W����ʓj�Zk�'��I�j�Թ�]��|wlF&�s�0×q����|�����%�C�P��U-pl����,E����SF.�g)����Mr�^Ao0٣���r�=ud����M9��S�������F&�����a$m,���u�og3<\��<vJ����6떇V���4bk�+�l�Ql�`���a)PL�&HL(c��������0~���Y�܌�'ަ���ѩ��7�3�_�@b�Z����9�^<�&�r�w�-�ј�T�&�I�7��ՎJlE&����F&�b�)�����B��������Aɰ뾌���L���������55˚����G�0ۮ!���֢��Х�9xE�/&�r2�Iy��Jl͂�v���z14K������^䭶P    m d��n����6-��l��GQ3A�G��	:]�A�UW,X6�`txc-�F�Qi��.]�ш�p壓f9�Y,E&�r�ނ\�Ng8�=�����a�\�؊G
���3332�QP����+��~|���{׭<�����L8L��t�jl��w�SD�X�4#�g;��]�Ynڃw��;щ��fv�u�˞N~ L�!+fIua��3-3�5�f��sSR���J���rќ|����{�w����<��=Hqs%�e�QYX�UL\�"%��,*�D�Is$�V���$��4��O���V�l3 ���`���Xu{p�	���2щ�z�%��o�&�r��E����<�g[ſ��aYZ�d��.�F"D��Mp�)�;������bo}��ީbjF&�[���/�)����	@�:Ν͉��Qu�7:��̓�.�ˣl���}��6#�v���4bjF#Ev��Ao0ؤ��X�NZm��x�3�z[5�"Ũ�Ns�6��S���ztL!�0�����=�n�h      �k�d�Ȼ�mᚺֹ�5vf m��kCaP���!�⪫J78��s�ɥ��κ����َRj�މ�\���v�^�tL6�bmE\5�U'��Y���w�zN�~
���`0Ȑ�;�/0H�8�6g���17{+��鑸���Ʒ*�֌Q~w��rSb)P�z+��Q��s�q���wN=q3�g����[v�j���M���/0"1�ˏD�n;��b)5w�!M�8�#�AG83)�����<S��[��ո�Bqn;KMA��s�3s��� Cw"�r�-��\��;���}��ǣ�J15S�_eļCb0�g�)5D�t�F(E���<����3͢g#�n�-6K�ɰ����3+z�bU��Af��>�,�=�ϻ����s3�c�6�
�27\�`��ړS<?��Z�W��;/
���&������Q���sF��ȑ���3x�;�w�'[�O@     m�r���cY�[XW�*ʩ!u�d�]�:��)��e��= 6�$&��*f^!��u�MQ=�4bk�15)mGD�V9����ޭ�4|ͮ�oKR����߮w�w�ys����] )l#̓0�bf]Q��M9���9�1�8�Y��Co&�B���z��HE#]��Q�؈M��&���17��|�Ϸ�����U�ʪIivbba��؊M>����HŢ3���N3mNU�t�q�fD1JQ��sWUk����4�!
��/���<��x�s��c�� ���!lH�N�b	F��v�R˔�ؾ`e)�\��2k��h��.j���GD��];bn�q�`-����SF㵡�U9���ض����\�{��x�2��uR�ؚsSZ�\�<��\�c-E���bw�&�b>Y�w�%;����x������>!y>=(^JdM��ɕe�U�v�46���$]��*�J�B�i��X��VVJ��
��%]ܝ����	�Y�Yg����e������-�  [h�P                                   �tfŴ���S5����j�����Ũ
���4���2[�-����:9��W%�s�*	a6�3���+.��=��u����t��L#��37[fX�0t�ZZ�Y��*P�yj�T��ҍ�hڵ�-40��ű$��ʱ���eS9�[suy�#Ca���ĳUvnfeϼ��g���9m��     њ�ۑxHŪ�׭nf��r��M�t�v�P��O�燥U�fQ����y����\���^�s�ȅ��&�R����4jjF��s��d(lD���Rmꥒ���Nbj��Ι����u`5vc�|һ�i���}���ڌ[�Bh`� ��M��*��N�#QT�� �d�tM���D������UI��r5ۑi����&ffff;�L��yS
l�ԍMT�z�Pؼ*M��ފZQ��^�F��5�nA�N�c0��9I�/�o��|xz�\���?/{��ܟ����֪���ڈM��#¹���1x��榵��"��0ۮZ�cQ���]
h�ԏk�I$��16�G�2e�b0�g�-7yQO�� ej�fֳ���Ù�onyE��	c�ZmF*�{nӽ��Q������;�-D���y�v�XUy14u�N<��nw�d����=��P      0e�l���"��2��im���p�6�h�ޝ!6��UX�a��Q;��_w�Y���~VB�3���rl��qB��Jm�)7z�aF&�sR�j��x9n9I����|����]��P���=�l�o�&��q*�B��c%�ň�L�Ia��M�stOdM���jkE�a��u�M��ݪ=X��MH��㚸��@m��k���V�Jl�0�m뵥�hisR9E���=3!��FØ�����^`�hF��s���%�u�G��_��1%��mm�]g��;�g����E��bT6��E��z�щ��V(r����qNۮc�2ce���\^{�T��x�s���^�n�]X�2����b�ە��LQ������N���r�\M�M�)e�������U�y1�w�͜s���3��m�      �cS�)3uK��ީ�x�\be���� +�R�r*�z�LE)��z���y�>�=��t�h�b�iꥎ���.b�	����ZmA��.�����S��E��{�@Z۱���o�7��p����b�8 ��7��n��L5c��JP��"h�և1ک�ꋅ8�|��s��ɝﹹߗ���YYjf&!IG��49��Q~w��rSb)Q�>鿺bb�\��|�����>�/g�W�i7$ �mdu�F45R�V�K1sIY21�N��W�m0�4l�d���6rR�.�]\�e^w\a�����f�4QRU���h�'2�;��f9�n�5�D��]<�{�����Ul����)�DN��Ai��V��)�Qb�jk��.��D<h��M��&���bh�娥�iyZ�a��n��|AI�Ȃn�fffdb��	�]�z��O��'�Gﻔ�ؼ0H�6���5뉣�}��_�=T����M��s����SF��f��3%���3���9���       cY����2�I�50�""%	F[I�&țR���>n�o��J������x��/	�Q)�l��o]�(��.bjF��t�ٝ�F�Y=�AF�R15ۛ�r���{��,M/�~*����&��dG����Ow씵*���0�o>)� f'Sr-6^V�&�Z;��S]�}Q����1�)6��Y�ޛ����s�x�ň�>���̨VV�]$�2^<�cx��2g��y��^�\2=nrlǶ`nJwmX���X��\�bl��D��nv�sQ!C{C�G�a�}^ӡ��M�s�������&�	_'��Y���=z������1�T��v��D��)���1�M����Hd��V�׶��Qɩ����y9�&�V����8�r�w��Lvʿz&�v�o	9R�j+j�\)��r���bI����F;Z1fe��q�'mG��u�L��w�Q      
�SBѫu�l�.Ь�-r6����u�V�(�
�l1q�%k��=��sy�g[�Zr��xc1�M���vV'z14�U9��*b�M�D�淢h��.bjEk[6�⪫qp£Le*w�zz���~&���)��yO�xEو��O�Ǩ�N؉G�떛�_v�M9	���=~lw�z7����'�<����\SC˻��/F&�b��ofJ����|#�sW�t�/�h�J�|���� �]���Cz�a��ٵ��Tf:�@�\5w�aM��y+�>�L��ʈrd�u$�;��'mD���M�v���,���wݟ0m�������L�a%��|�7�{����fffIw�����b|e��o��/*{�!M�e�o[]���[�w��J�f����7��f`�6s9ƨ�����h`P*�j1��mad���f���\�d��j*�F$b1��j7�H�b-��V���R�`����L��bF�x�L(��G�|��6����X_~���=m�*�� ��4�                          ��      *�df@UXXŖ�.
��5�(�m���K45���(�B�@��ܤmn���ق�4n��S]LJ���1�6-p���kL���TP�&�7#J��+-#��^ �[��ˮ�,՚��n�'���頎�b�6րlX�mh�s��u�Ŕ�S//	�r�g�H ��&a��1�P�Tz=�n�y�J""fff@     [X0+���m�#n���UNèq	V� �('w~JA�U ��YKEI�W��ߺ�u�z_�d�'�㺩��ueWN�N���*}��񸺻0�b�]x��<��|��|��t^c�c�>Oz/��{v��z���uz;�}׿ bԖ�ܴ��#v��ނp�em�~ ��G�Qݎ��B,U�$�X�xk�|�_w��������<�/����YYB-�5�%�;�3�kɼw��k4�̘ʴ���dh1;�{�����0O���;��;��;����*�n�vR�y�ޯ|_A��Qp;���";:��|�VA$M�.Es�	��|К���Ŧ�� �#�@y�uu�16a|R�H;�9�8���67�
rl�Q�����K�ꪳ6�@     ���76]F%5+%a5e����e6�+f��2�W��OUF,�����ow����rE9��U�(�D��qy\�Z�� � ��#�����o�6�w�[CQqC�R�9�;��w61�A��3���fq�>�콀&Ե��f�Za��rNH�"� �A�\��M�A�[��A%�-T��	x��X��ͷ�� �t�x�@"bm�[�� ""� �4�$kY�U���)�qx�O���?4����;��=���0�5+,UZ׵�������"7~��z��H:��q��R��qi| pD$�G�����͐0�"�H6/��v�A�S�����c�\�:��$qwqr^3��? �VV�֜�2u�go6�;��D�A����L �.!x������Z�R���#h���x�{s�6��� � �(s���r6�:�:ݯ�AM�P7s�������zUUn(�R؀��'|��f � �T��q��A�Z8�� $�x��9�фD�GDCDG1|g|�`G��h���)�����=�?�k5����w�舉�     �8�T�fe�)[l�.��m^�u�YH�jl�b�|d��| L��d���:�w���us�x�=�*�p���N�Gz:�\�k�t̄��X�V��qӿ/^�ן��ψ8��<N��T;x�Ƀi�����*���o����g܀6ܕ�U�XS�ψ�.��lNM��O�N30FN�s�#J/��R)va�ňF��`Bh&^�Lֱ�kjݙ*���Un��u����Ƶ�$fh���,Y)�g�&B�Yf�F���H$��� �4e���Q�K�1��&xX�Pѳ��y/��o�6s��k��H�(��#2�fffff%LLB���wx��Ό����:X����%�q���x^@Ԑ����{�zl��6e���6نYd��y�:�3�+�p���S^w�����{{�s���s���8˗����O/�l�      b�n��@WK��m-J�K�s-�V��a�Vf�<��UX�J���:�ʺ�u����﫝C�^�O�b�d,���}��>)�N��333!Sf�]!'s�ٜy���}g}y��L��*�my=�0�\�`���Sӽ��a��>���֌"�>�=�c=P��>3m�}*N+)���K)���}q\��/�bz=C��h�=33331�dj�:�^�}�q׹{V�=��L��ꉶ��9��Zy�_��(��~�K����Sf��~Ǽ������<�^�����T{�3`9-��M��α���s��3=����m�      kSm�Č���)�=V���Sl���VZ��;�'\������P��Ĩ������oI�2�����~��}�J�;�22��ެ�u��|�s��332�1�Yr������D��y��{��t�E9K��'�67�~1��ۚ]>��{�ǿu>�,I���IWzu|��VvND�Mӽ�x��c4�W���o�K��̿> �&J�Vkd���{���"n�I�窉��H�ތ�Mswfs\+��a���eR�K�[��8���$��w��;K��Ϡ6Җ���]�%�ߤ�\����|��������Y�\���8��<�6�a��j����>o�y{Ҽ�2��m��O��"�KU�^=�Z��~APQ�����6>��/��m��m���"�E�m4�97�x��3�J�h(b�VN5&#J�Y�SI����(,�B+I"�
�A�R$¤�bD��1rHM(��,��u��H�I4X�9��B[�(�j�]P�-i�MV�(fʔ�T�ؒ�(Z�@� �b((�EA��/�u�uU@xf�bu�82R�*��׺%�6�Ua@QE!�y��:�o����5ݏ��7�>��
�?������w_�71�7���t�d��F�V[�3����'��U!N�7E�c=sE�A

��r`��7}=~s�}O��3��^A@;��_�z��>�?{�Q�>���S�������TE����"D��dY`�z�: ��#Y�Z~~�̈́�<A�y� ��╸��)�z|���-�erv�Gi�_"����̪
<�z>�]��X����/�~����,{�/&}���5���xh�R��qrђ')3�D��|� 1�%���X��g����#��o��:`��~�����Ǵ���^���yߖ�zp�۞��l���獠z��(ߍy'�=�g�jXq@[�IdBDY�{�/L��FXăE�$RAc aHDP�DHEQ�U�"K)��e���I*�(,RYd���
�eE�B�J��d�REYV$U�XE,IJ,�[VBʑe��H�l�e%XYH���ЫeAJ)d�dZ��|��
�P��[VIVB�UbU���,�)-Yd���*����XUR��H���"�F�`#"�m��U%�jZ��P�-H�2,�"I"Ȑ�",$�*h �**/Ř)����g�V�l�{�s��a���n���=c��2��������<L���s�1!�0��!��*BԅT��R�+_��8����>������g����`�
_A�c��@~^��<�|I���<&Q�����C�w��������}?���z�&�?��n�D�������r�j�d��|��_���:����6^��W7</�Z`Z\��1&\z�N������e��g�>3`s��Ϗ�߯_��i�d���m~�6/�Oyw��g�W��,��$����OE:,"0�+�>����6~Ϗ���{u,qGo�#�ůe�,��S�I	�c�?@���Mϭ��T�<�C��r"�p���摣a;O����*��}29G��|���rjۑ����ϻ�Ǝ��$I����������r�gW��#�񊣣��6�mJ���함FT
 �H�)�(9�8\��{�\��['�am;���`l��쬎����m�Z�_�\���6��|�!5Ѽ1��$$���|P���~��q��X;��� (���_���gɟ'������������eZq뇿�=�?w��d����3��|�E���v���iz�t���|O�:��	��Ԑ�3�綏M�=����l�['�5%dd�k��O����! a>��s����~��͟	��z>[�������������/��tS���~>�~��ƛ��1;u���E�����z_5&z�=��g(�o�M�� ^�s��`屠.������g��&�A@8���ڼ���Z�F�t�x�*j's�̱�]l��n#���.�����r3�^�U��(#�uj�6�='�Mz�s6zl�����rȡ�<����A�Ab�"�;��l�����"=�"���ߗ�?.4t=}�QDW�OQ�w�TP���}���_?�}Niw���/��{O��X�g�C�
�K0�Q�`�ϭ���H����)�2 