BZh91AY&SY�
=E y_�Px���������`�=`pt_x��` � 
    � 1�-�Tl��MRo��R��&��  � �@���1112�@0��4�挘� ���F	� �i�Q�5@  4 �@H��jy��!�A��ɡ��= D�4m4�&��&�Fii�#�K"N�J*��
�b*	D��J?�-�A<�T R���ګC�6BN�!90��A`�A�>f�����|�G9���1�����9��P� �2]E$�CAB�I3R]IuE��B��I"�K�B�� �1EEQB�B^ �t����Iab�Ab�,T*  HH��&�B��B�!B!����h���vn����wy���������W��̫?:��Wnn&!YzkUX*���S�dIqw�v��eT0�{ǉ����D�ʳj%�n���a/�R-���-������s��_8�&��mi��J2@fl�B�����i٧�|��A��^�����O2��fM���x��XN�ɖ���$J_�=o@�s%\32��niJ\-�֙�.Z�ж�t���Y��]�F���R�\wqV��&|u�w�$��?�ynۥ�#"�6鼻s�:;��D�����ӌ�.������Ѯh]��q�wT��t��R�ݸa]1�fe���f�m.f�37I�r�ij���+Ku�]�9L�H����S[�(�uVTYB�R�vx��ѽUu�ܗSM4���m�    ��m� ]�  ��l 9�r    wcm��    m���w�iF�פ�4X�r'AQ�0�(�m��*�S�r�t#r���EE�#�c�T�9�Sc��Nw'	ק]��;��w>.�{��B$N~�봠�R�R�
t֩M�۩ƥ�S��*�޶���`BaZR�N� A	05���BøU?bff��<6"#bv6���8����#����>���a�gC��nw`V���.�J�{oN��݆�z��  ���:��/��m�L�n��Bݪ��A�`sT���G`8�TfO�	��I��M�n��j �G�o��E�#/!�%�=<K7�-���Y3�38�UV~8��,����:Y��!��N���}��"(�eE�2�&��m�M�]X��Pf@�	��[:��fS�`�U����݈,�sȸbp� �~f`���k6J���8_�����!(#@�jS�~D󟇃�8�,�����4ZL�1���&�U��5(r��`�%0[KY���K��`��9�	�l��L0b����uK�������#���ѹ��	Y��&1
��IL��DD�S�&�cfgީ�'^\`z���Zk����L9$�C
��\�q$��'Ba��r���@�n� ���;��'�g ��	�a�$e�3�ۧ453���;�H
, �� �B�M����(�R$0Y�.�"w ;��>^'Ʌ�+"��*�̀���X,� ��*2�[�r7��/�?��Af ���=��-	-\�v�pn��h�(덌�׊�0���ꪧwz��ʶ��DCZ����N��#A��r!��	 m&�ی/P��w��#v�6y�q��$*������XC}���VT�@sB�!˝^V��ت�qz��q��1���f&S�ҝ(ո��1>�ݑ�$� �q�sOn/��ּ=n�m���oxV;��R��6���f���>+�+т�:�/X  ��I����;�jniF�������ճ�UT��U[�����c�4<���#���9�Nd���=��3��L &�P�(J� �����@n�fsѴ�>'�����zg�#��E�lH�ǽ��qҶP;�I���e'�D����a��j�<�@��AL^\�N�8�;8B�D_9����l�C��VǊ>�V`Sѩw��}����˺�J���V�J���d˚����Q��OEht��"��
e#��Jb��;*� zS<��f�LU<Ȍ++
��(d_K�Ո�Q�.ٮ���N���T���h(R��Qz0=ٮ��m�޼�ݞ|��=׋&�y����G*��0�}@�!���!��@�NHQ ��<f«��J#5��I;�5�E�V�w�5[Nc	89���#Wkו���T5����t`�w�%�a�<���1����@�#�S�}ohۍ���>7�*��vUCE�m��pq�8���u3rA3�-�QV�v��5��w�0�)F�w�",�L�<�S�z ���#UX��}Y]�*�lNL�˒���U����d�K�T�P��	�.z���6^�c��)��P�t��������}Ȏ6�{��&1����S��XQ�;n�9`">3��I`��~e�BpC����ۜ!5mmd 	��;��p�"g��D���	0I ���~z"���i�BPp^�寒 ^%f���b��"�����%���ǩ�P"3j_�T`��g���V�vF��	�I�CJ�K0E\J�gjU�XNVӖ�8S�{�X#U������"�� �A!��xE)>�WO��y�r�aY�ਟ� ���X�~w�z��}�Mc�Y��f�pyګ���d�ID��4�H���z6k
wѦe�L'<DF�=Wk	�0�hڝ~��\�EE`�	Q�x�$m���U4{�s��_K���"kh�[��T�W_ [�Fqx~#�"�_���2I R��u�|R�/T����U0��^�l qUC<!Y��	�f@1t$�C���-(QEQX�]��QEb�*����>F�aA@B�I������Ŋ�X��E(���
J���"��R��,U�X��"��U����R�t105 	5�VRN8 n@P]�Nt(&��03$�*l`��&�HO#3��ƓL/@�c���Y $C9�:%hM~�{����t����%��}�~��ʸ�t���J��w�=����ZSA�P�B�;���W"�v%���D�T2�zc���Oj9?���	J�&włRCh����|����$2H�������H/�S؝��؊�� <x���eH\��<�	Uh��l�z˅T�B,�)�f9'��H����>.��!������v���V�X�k�U�&>�ɏ�l��^
�=2�H�X��b(FF""��!((
E"+"���F"�EUQQ`���$Q���Y5%QQ�"��`, 	�> ��)�1 Z�-�{~d�d���dIk ���Ze�TR��و@@�+!%H
@R0�"@��r���r;
r���!���;܊&)a*8�!��a�ޏJQ7'����UBM�\����1�3�9����3"����,[�t=�N�����K�~�I��Oi��)ͫ	a�����o�$ZnL~���f�׍ E`rEP��h03�����h`:�:��M��Q��`��0ɬ���<:�踂%@� �qӀY\�FfY�ZQ� ��8 `)V�ӱ�\��U-1|X�+Y���j�0!d��|٨Fl�r*��F~��E��N���ۮ���;%2��*P���J8Km��c�fI#��a���@�T �D�H`m#��uP��ͷ?�zڍ��i$*���擔PN O[ΉL�#s�<�ӯx�;z�{�D�*��H�`��ؘ��`�zYC�u��H���@�� pp��fgAg0�Ɋ�x[��@�ҟ���ɐ]��@�|�x�>q��Ȉ�UC�����b�&�P
{yP��}dI��Pb�>���ie�1p0�\�Z��H�
aG��