BZh91AY&SY�Cx��_�pp���g� ����ap@>�   
       �@ >�J 
     o|    � (�        PB* UT�EP!
$�J
J$�$PE
� ��R�D %        �� !  �1�@ijV{t��*X�����Vv�f�{���ZQ��)�� QޔŽ��  � ��) � � 	  ,* � � � � >� �;�9  ��P( �XT` �ޅ��x���w]U����_z��Ӗ����oR�^;=�����J��U��֜�ͫ�ɯ �{�}��m�zu{�
�=���-���^N�5�˯]�������>�O^�<����Mzo�>J DD  �
�}��7|����j���]��N�����>���=��x�yoj�o-��	@=�q��k�v� ;/}���_zl�� ��9o�Ξ[����zܚU��(�}����r�6�g�{�=����^� =�  !@P
 ch���������z�&��o7�U��P>�}>�ܞ�^.����m{ŕ/�T��m�n��������*��^׾�*���>��m��ޞ���k�M�w �oz���&���9��כǳ��� �� @-*v=ʾܞ�g'�m]�}=|���R�z�[��[��,wW[q����3y[�E@���w�j���� ��&��{�� �����X������������K�=��nO/x^=��-��8 P       �	��U*��@ h � �"���T�H �     D��R��OA4�F14�4�M��T�����h�h�ba ��E?Т=����F &# bh�D�FIT�1LԘ�z��#'���x�Q>?��+�����Q��po����D �s��T � @�(* ����  ��������W�B" �T�O��" {�D@���A@ 5������J�(��("�?��[���������ڼ������oG��V�x��266r�{��y�t�:���<i�5���ݍ?��_h��(�HTRQ�	
�+Z�zi!q�Th��C�(#�nF����	!.��Y4Ce�OO5l3N�<�L5L�%f�8j�v��h�V�M�*F�x᪳hٸ瞜���,�h��<0��Xg���xg��߼�^M��=����Uƛ��I���B��y^��߸쇵��G+5��\�cϾ}yı͘���f��}Ǔ�@�^K6x�*��4�\4\����D�5�GR����+~��7Z�.7/��/늲+v��O�nw2|�=�g�X3��g{A%!f9�R�7.��ʕ��܅PT�K�*%�^�Ѱ�(�	#R�4G%�m2Y�\C�eU�����A$�i2Y(	R�]ʀT��T��U��$�aP
���I!P����B�q�Sa�5~_*�7�>_7�~7G��GW�8k8�E�+[XT
4*�]㡹O��8n�}��ˆu�`�TZ�A��с.	 �	�E�5#auC����h�l
�T������^<�����^\7P�&�y�T��q�fl����BIM�r��۸�^��·HdʽofL�ryS����n�O52���/�sͅJ(��*�TjRoE!������Mh񭄷ԅK
�5�S�O�r8��ۆ�=4x��=2BY�����G�����aIr,xK1nxm�[l�3HUK�(Q���s��cW�����A%�"U%%Lt7
����^���fh�����\}n%%B�IP(�*QiE��˘����&����B�t�*�¡`T�*��Ph�Ia����*S�I
�YQ)*���d�^��{#e��M�5�8��tO=5o!��Ç��_��Qq�����мy���d9!�� �&�n7�Rs&;���ގ����^W��_Eҙ�#c�J���"Qfa7p��3I���F����HT*c�Cff��
���3Z�᠆�j��T�F�3P���ݚ�ȵ���ޥ�J��Y�M(�n"�&��s��ܲ�5�ׅ&B�+=��x�r	"Se��o��^�Sٻ���^ro<ֵP�ܢ�ؓ`U!U�*�ea=K�
�i���XC�B� T
4a��i.	 �TB�cX��f���8n~��i֠��P�0���g�H^�m�xYMʯ|��n�e�P-��H5-aV�!
�F4JK�mJ"�q��c�K�MCf�L�be��J-$����rQA����y���<w��\��L߆��$�̆��景/P���5�4y�	�5���&�&J`�}1.R@�z�e>��5����a!Q�X]/���QAw�l�� ���4Ӓ	 `�$�k���SG��̚�h��M�����)$j�P��#KP��~Ԥ�.��l�yLԭy{^��둫#���>�Ph��{�����i�7����Q�*^f��ɭ�kP�^Hz�
-�nx��tMx��e�5�M����Q�Va���~�����B��eY���F�٪(����Q��ZF���2Qpn`�nмB�8��oy�y�^���B\*�oXo�����,ߤ�eʋ���d_\�]Gt��ux�Xl�-5)��Kr�S{ߥ�5�皨K4�Z.�J��k��^kCE�.I.�!q�Y�n*Ĩ�{pI<B����kACQou�c�PPar��L�Fl��ܩ�[�֦���Tl1�v�dt�َ����"US {p*<, X�eP�<Z"Ō!$`�Ke¤7!s��%�X�����Tp�K#a�H$�H��T|k�6�d457�4��dij��Q!PI����{�%]���zsp�a�!E�aBH�pI���
�%!Uu5iD�F�JB�a$j�Z���$�T�QoZ��:<�jH��BI(�U�0��8D��Ie�PԠ�P��Q��A$8P��P*-5�Ш�Tʈj�H@��A	Ʀ,*��A$@<*P�s��g��y��ᒋ\�o+Z�^BH4r�0�_�IY����&��B�ߤ�=<#W�\l�¬����Cۡ���RШ�L��F5U6J-ITR`J�SPI�I�P$jRT�D�4J�-�E��Tj�u!$%UBD���IHTmi��A.\�(,�wAxQ�(�A$A$JJ*����(,.[tY�����d��y5	qi��*�,�H_(��3%������toP�rndBؕ�����fI>���"&�"���Yee(ɏvN�ed�T���T!q���E�L%�) U�&g��&K�&�kea�jQ$��J���&�*�,�,���XB���j�eTe���oVkO�U��'ie��q�K~�*=A�J%K��͞!"B���4�'��Vc�u�_�����5��R�}�����sFyZ�®���xl*�љ(����s��HQj�
��z\
.4��Sg�����Z���V:ӛcd�I!w�5��Y����r�%f��Y����75 ������P< ndBѿ<�u��.4B4Cmk�#{�j5����2y��:�^��W��\,6*-$�0�IhjSd	�Q�i�����,(d��@�R,�0��EX\
�+Ur2L�
	#$��HITP�$2T��e�'�[]�%�J�*�[�뚦���e�2q���vd.�˅7��P��1�:ݗ�g��lg;�-�ɻ�\L�H7��	ȗ�T`T�Q�5o�Sl$˥�����p�.�"TRyBKJ3��&C$�aR�w���[�~�����jQB�-�I
.\K��$t�iȗ�[5���Yg�P"�;�a��:=(͋4���
,��E�� �w���q���PHU���
�z4L�nf�gdTG�&�$ELLT�E�,��3;��!yj⬈*H�ꭁqI��	����^h�ܣZ5�4]54�Y�=9�
���0��5u�uFh�
����r�$'��jں4�tX���O(�A7 �VzSx5T���&�pn>�q6J�P*	 ��PM����&��	pK�H'�p���ʐ�\��*�5����j	�M�����|�p�4��7Ve���=�y3��\����J�H$��
�H�5Ȥ�n	�A$�I�I�Iʎ���F5*I!21�D� po�����FGM�,��|n���2�f˛��.�5��*kx���Dj�
=���I!	cMA�E��p
�ʥ�(����$j�/���y����zK��rj��e{�L�	���$��j	S��7�7�ʽJ7Z�j�1���M��o�>p�ט�&�-��7*Y$n����^���K��ˁ.q#*p�����%0�Qp*�RF��d֡!�q����Ee[)�RL.�t�ʧ%��~U��Z�vg�����Z��W(��7����VNy�>ѳ^^jI������C������7�J�7��m$��\mj4�F�]��+*5�����	 �TA$B�!��B	!Id���}P��7h*4�L(aT$�B	!R4��Y�2%^9l.!U�TZj��h*	$�H$�E@���ˑ�R�B��	 �	(I��4A$J!��Ja#TTZ���A$jME�TJ#PI�I�I �(��ĩ�*��$���%B�\���6�\jI�H���{G5VJ�ݘeI^a��^���\(%��J�wfaP#S6�K�������w�]�`QQ*F�!Pn5�m��U���hܛ�f�%����Q�Ie�$tFJ�P����H�j7%�H��z�2�,�5&D5Q�5-d����p�k����NUUF�To1 T�d���R�ZT
*%B�[�/F^{���'�f��r��L�+aAe��Ori􌺣�3^{�e�<����%J��B��T@��|ud�*�]�U{�p�yN�|���f�������"{~�*^��,��m��f�jd֨�x�B��F��^j��Jc,�c7�{�!z��WTU˕7+27ʩ���ۣۗ`���$��n݋k.�n����U����u~��?�p�����F�������             ��                 �   ��               8 ��   6�     �  8  �>               -�                              �>                                                                䄎-���      m  -��      m�m�m� ��Z��4�@T �M��;Z�Ŧ�   mm��p�6��l�� t��ldY�Zf�$�(6u6 6�Ue���8� H $� �I�]�X[�:F���� l���!�m ���(���   $�6�O[7k[�6�l 8  H ��m�-�I3kn  Y���e�m���p4^  kZ��fʇGT�P�v�[���    �  u�ISN��$m���i���z�-�$Ӯ6�Wh╼9�e�Mһ5v��V*�U�
�U�\-���5����    @R��zАm�m�F�H[G     �۶�t6�ͳl���           ~��  �J  d �� 2 R���� )@A��   -� d �� 2 R���� )@A���� (0 8�� -�         ��J  d �� 2 R���� )@A����� �p �@
P`8 p (               ��       [@A����� �p �@
P`8 p (0 8���b$�         � �p �@
P`8 p (0 8�    d    8�  6�R��                      -�       �>�                                           �     �>                                                            �     $ ���Ƀ�Alh��H�4��[*ʪ�+����mpm�   [x۲�     ��m�Mn    l�kt����/P �l�@p  6��[� �   �[�m%k��    I[ �g9�p  m Z��-�@�v��
�j� 
Ft	fkRt�h^���Z�-�m �i �[��f�h�e�mm� �l�k�R��p�y�h`
���Tq,��u���܄�-O������5�Z�HMP�WM���X�I�� N�H���5t �X�i�|lqm�� m��N��� 2 R����l R���� )Cm�)@A����� �p �@
P`8 p (0 8��  �J>��� )@A����� ��m���L�m� Q�Q����۪^o�w�|n�shj��lbv��A.��I���B��"���,mK&Β���m���[l��v��]��H����!2%��zk�*��[|q�@��
BiV�ګ� :@rAc�i$��δ�+J�mU:*�6�hи����Ցd �v�hh���  ��l e6�U����L�Q���  �f�Y� KV�m����1���kH'M�� h�@l��� �@m��J�-T��+T�F�h    ��m�I˦Ā}��o� [x[M۴� A�a���A�Ö�V�U�W��-�`5�`m�mm�Uj�6�Z���b����m	 kRT�'$H�.� kn� �"��2J+�p$u�6�v�[n�6� ж�   ����[V�H��a5P4��!4�l�a��$�6���5� �  �g��+v�m�m��v� n���8���� z̗-6��%rpOa�3Tp,��5�G
Դm�"R�Tրn�k6]n�M����&���I�E������6Ӧl�5n�[לp�� $ p�;�1[-T�UG	�P��l����<��i�y$���N�z:i�\��B��r*��i��[Mp�"Izd��պ��C���qR�m<�8�T��ąl�F�ٜ@\ps�����H]�T�U��e� 4J�[p�d��n�l 6�e���ZU�T���^��V�-Aƫ)WVS��j��,��z�mf_,�kn�8H� m�t6�Yt��l$4�-R�l l�V�8�$���],��aV�!ڀj�,`v��Wo^�ai��ZR�@6Z�Z��E�J�QeUuJ�l�*��(�T�Nh��:�	<K�lU�EKUv����8B�UIm����9���P�G��K�8h	vZ�Z���QT�UTG�]���d�lUq�mG
�I-��@,�z���$�;mT���e1�ef�+[!m�mU,pU@6ۀ<�mٴ�X�u�V�ʹ� h��mHM�1�yz�v�u;�H۫ �;E��cm�d��8 �� � �C�ݶ�7e��r�p�Q�K��UT��tQUS�d̮˷U�
B�`�ki� ���a��I  p[]�K �^������`k�eN��B\m9��uf��/m����UJ��	�.UۛR��n)�ڕ�'GP�K�׶��y7`S�����S9����		ey�A	�0f�l.ʫ*�8����[e��.�` ݧN�v��Ll�IAlN�T�>��}m�n�	����V1{(�ۖ������˃�MN�hU�B����z�j�x��';t��v�8iV��7cLM�8A�S�,�r�υ������g=�\�k]m@J��Z��GA!4�Sj��	�U�yU�W�j���6��8�`��!� � vܴ���u��$�$���ִ�[# t�J���5m�k`6�wm)�Kh[�   ��c�$��m&�sf�+���(��	 M�;Y��Vi�8`��"�uUT@ �k��Zި�yv�����U@T�J��lJڭ@[D��jA��<m�d���e�nm'm��� �N�8^�\8�vH t��hݶm�-��[��#��>����� m�8�@�	 :�v�h��*�I� ᴼ� M�ɉ��[v݂F�      $���m��O��}��6ͲM�M�� ��888���#�Vm�"nY&Ā6��,]P�6`%T��vk�^��f��Wh�,��Nw��ϟ���Y*1k�+*/gR�( I�al5 �Rco�gz��]68�WF����ȴY�vk����(AT�8.�[Amm��%�����ӌ��ڶ�9m^M��s�F�m����\b�X6�rxtT�[UWV,-�T�U�
UUZ�k��b������6�p:[�ƒ!z˱��6��֖����`:�ȵ*��G*���o0q�UElT���et#[s���p-�zM���j2��V��Ⱥ+�lq.��
��N�J��.�ģM/��O��Tl\��܁�pX(�ђЪ�=�)j���9�'(-��[v��;U�ͼ�ܭ:o�m���p�5���p �4����dj+ļ��UXw��ኪ�z�R[ic��V�l�Un�|<R}���knږ��`� ���-MNR��  �2�m�bF� ��i��:@�fհ��C���p8�	l��	e�Ft�%��m$pϯ�>� [@6�m ��i�m m��l F��`�[Hn�� �Kl볫"�*��4��g5�ؒx�Ӻs3�VU��圠@%+���Z� ��ɮ 6��HMMK�r�ܑ��E�V��YV��Z^�3R���M���\�IE�	�����z��*��Y��?��`'�z��#��R?���'�
!���w��?�L2�*C�"lW������E
b -�Uݧ� ;P�S�=@�"��K� 9�8 x�<Oit%@`8b�@���A4� s�'��H��"�ȡ@��ҝ��_�qt F*Fb"Dm�lG�8*;O=�A�<W���A�f&0�Q<<�
@_��� ����W@��G^��q@3��i�^p<A�E=��m k�W�Lت:QtE`���z
��B�(�| ���1"���H�(H�"Fc,XĄb�a0�B��@�� ����$Y$`0�J���0A��@`������H�e �Ta� $�2c!"$YJ�H� �`���p��1dV,Hd�@ AA�A�	!=�4'�d=���J�HăR@H	��B� �e
D@(�R&���$E4���P҄ �)�.�CJdTN]�=4�-3\v�1J�W�T�0T6$�< ��4���j��P�������H�<%4����J!�
����rP
��*P����U,6���AS�Q�Av` z�;<?������ �O���K��F����9��"���$�H$�H$�H 
��$�H�I*�
� ��,�H$�H$�H$�H�0�� �ȨH$�H$�H$�� $�� H$��$�H$�H$ � �
��	"$�H$�H$�B	 ��"͐I�J�A$A$A$A$A*�I�I�H#pK�@I�HE�I�I�Y�I �aAD�A$A$A$�hA$A$A$A$A$I�* ȀȈȩ  Ȅ�� �	 �	"`�	 �	 �"H$�@2	 �	 ��H$�H$�H$�� �	 �A!�I�I�I�I�HA$A$A$A$A$I�`�$A$A!�I�I�I�I�HA$A$A$A$A$I�I�I�I�I�A$A$B,A$A$A$A$	�I�I�HH�D �	 �	 �	 �	 �	$�H$�H$�H$�H$�B	 �	 �	 �	 �	 ��H$�H$�H$�H$�H$ �	 �	 �	 �	 �	$�H$�H$�H$�H$�B	 �	 �	 �	 �	 ��H$�H$�H$�DdDi�I�I��i�gw�zN���� ��� m��   m�� -�l �	      6�            aC � 6�g�@kf��R���g�6-.�J��@��u�;%�U"��:,��q�3v	��5 :Q�گQ���-�d�l��$  �  �J-�G 2 R��l `(0 8��� ��� 
P`8 s�p   )@C[Ŧ�h  �   A� ��    ���`       �   ���6���i&6�6�.5�iz�;]0z�m��UW��d�Tq��P;Al�\v��͵�=k���0M/]�%rlH�� 6�`A���� �p �m����߃�]�j���ѣ*T�4�nn���g��;���/�á�(63�y]�VV�,�ej���Dh����J��X6�j���Va�yh
�a��Q�V��E[�Y8�+����U�����*^e��j�M����q�)�f��(\:x��h��u�%㥊�;�;m[=ґ2���w<uZ6iH�)4o3�����ѱ�v\B���閲�n�֞rܷH���R�ksRKFkC�� H�$�*�<����'m�
yu�%t&wWe�8�S�vt�rulZ��|��_0��f��LF \���{NݤŹ�3	����n�]���ջ%��4���9hA���/\�� =��Z�*�Y�h��2F%�Wk�\�Ϋr�Rk��.�j��ܪ�Og�dߵ��m�Ft���F�wM�EK���tz�R�O��v�FS:�m��؝�L�v�^]���������{�����gZ��>i����H��w2�Y�Mũg�*��;N��,�����������v���`��j�iJ/e��7S(
dZ�UU���<a�y+j
!��v�z&�yǆ(�!2�j�C W�	��Ъ�ex�������˺�v�	`6� m��F�s׮�+i�ZȥmmH 4P�� 7n�J�@۶q���ے ְm�l����k�`N5e�׮#v.�;j�ԫ�+n;n�0&k����	���u�9,8,�i�m]����t������vm+�/n9�g8v����n�l��51-��`���c���g��j�ᆰy�ދPi�آ��	��9�h(!j:/+Wwmʻ����6��`;=�q��� 8���������U�VMݑgz���� ��^ޯ�p��-X�	�x܋�j�u�.W�.V�*�8qJSd�6���swX �W�.V�*Jp*UrU�.:/�7ėEXM������ J��O%X �QxQЃ"K�.&���&���� S�V $���i�?}��V��dC�B'�QpJ۪���H�HF͒
�ONݔŌv�9uI���sj9s&9"�m�����o�4��up03�F�nD�L�8���	%x���>���菠�� n��Wۯ� ڰ��cs&6��' ��0�)��U�	%x�)ʩ��*����˚� J��O%X �W���+���n���,D���<nE��U�	%x��*Jp�R}��4�>u�����EZ���X�N�ڡF]�S�u�[W������Xt�K�:๻� I+�+G�A*�8�J���'��$!Ly1D���o�4��T��)���s"P��D�R\M��sݘt���)����"��n��n�8�߱��j9��I�I8*Jp$� �T��w�܉��<j7 7wg �vi�7^��������5�G��ǎ7�-�I�W���3��6nm��]O&��u��g�6���bs&&��' �wy�*JpT��I^�Jr�l�
�&�����0�)�#�%8 �W�r[����|ib&I�x܋�}�up$�2�yt���*&�?)�	��qp�#vl�n�3�n����^g������O5LHDcɊ$���YT���)� I+�<��iI���m�l��+n��+-�l�dog3����'Y�erT�v�u�Ɠ\W��7T���)���F�&�F�.�ˍ��Q�D�$��}�upwvp���os�Un� g��܉��T�U� $������� �INp���	19���9$�n�3ޠR�Vʒ� I+�;�NUM�UM_�v\�� �%X*Jp$� ���p�y�/}ݒ$�RH	x���   �f�u�gV����r���6˪���|!�Ji� ��p	8^�:�ݳlH  m�7m�%�E��eiI�I\�m���W:K�+cG7b5I�1������5�� ttE�Uɕ	,�bۃqm�δ�|&E���2D�����@��ݐ[VS����<�Ǒ't$;NY��޷73���gk���z��n�w���wV��4��kCg��;dU=F&��?M`�@<sp8��Ԁv��43s�B��,DɎ8����׵s 7wU�����*�;��0���f�蛻������_L������ �IN~�<0�.���S�b�)' �^F �%X$�# J���A�%ԗwW0Mـ)IV�,� I+�n�8�߱��j9s&I#��������`
RU�zA�?u=���3q��v��!�#�]��Оtv�]���c��� Ν�ŉ6�ל��������`
RT�ﾈ��M����^+�$��Lc�p�f���C��BF�`&"E�r�`�dd $���*�ʀ��o�.j� �� �F $�����{���񥈐q?��/��m�� m��V�JJ��J�SD�3qtM���\`I^ ��`
RU�-��pF��{�D�qǏY�ɶl���f��v��w���܌7�1�<�.tM����� ��`
RU�$�F $���Ѓ"K�����	�0)*�K# J����}��'H�\mG"��$����� n�����A����ԓ��r�$�=��A�"k&L��Ng.y��[l��LJJ�Id`�Q*(.�j��*�� �IN �6�@M�� I+Ͷ���j��p̾�����"�ֻD��N�=)s=��g��Î���̡F��JY헉����� R���9%��	%o�����>�X���9 �ud`I^ʒ�JJ��J�SD�3qtMݕ5q�	%x*Jp)*�>��g �O�y�bF(�D���|�!�}S�np-��9%������2>�Y�x�t Ȓ�&���B�� R���#�[ �+�9RS�gи;w����O�a��.Km�@e�i2�vb���fulW�h�HL]��WnvՐ%����y,� K���)��� 3s�܉��<q�3����}�)��� �FʠU���*�/驫���9RS�)IV�,� IB���6��ħ�8���j���>Id`I^�����9B�NT�Ivuu_M]��,� I+�9RS�s��V���y�pUB�uz̻���̓.݉��  m��[�y-�YXmuD=����
����86�8�-��l-�knH  mmVGl	 ��kMk��:���� )\�곴Kí�Ƙ��΍�cDn�j�MZl��]��e+����Wl�+�S�zw%��uی��7�Dc^kn�wm�ʏ�/�|s��!�v�ډ��]��kR���C�ݨ�{��{ӽ���t��9ʠa���jZ��+9���^����5v�Է.��٪�:x.�U����~~���)��
c �F �t_�n%�RN������g��W ��F $����D�Q7��rW8%IN�,� I+�9RS�zE��q�$�s�p.y��m�� Z���)��� !G AUWsS�]M�`)*�9RS�wW)�9%��߯��}��K������%6S�J�Z��{VI�n.��t�u�4��^.v�j�������9RS�wW)�9%���5�������x�2Gqp��yZ碠�V��_5�s����sF�
ʙ$�������w,�U�/%��<���L)�~���&�ʚ��U�/%��<��]�"W���M��tM��UU�ܹ,�}��~��dh���Ѓʡ\���<��fs�hv��W٤4&�m��헙�د��u��x�W��o������\�F�*��%���*UM՗e����]��˒��%_r�;����>��p�PmȚɓ�s��m~}�n�y�������N�w˪x$��.�D2����e����.��f�^X�B��X�P���N�!�)���"U�9f\Z-%1����@��!с��ƥ�U�!�f�S�vcd��S�R�z�E�=��N�R��Z� ��Tlug�M�F��X7E"�.�����N ��#i�
u�� �T� �E�-yh��խT�򋚺*��&��a%�5�4j� �	�6D�W�q�"j��(��yHBd�2\�(�$% �B>ͧ��d�h�A�	��b�H(�I Y	B�0�}K@�K�)l���w��e�$¦�(p|�S�U�!�_,g��QlA�i ^��H"a��؁�ꖨl<AS�EL�+b�QN{{�iI�7�9��)��;et�3�1�*�/JH���;��$S��v���H��;��
y]�oJH���;���d�3
��2�.��5c�����֔�I��߻��"�)�}�ץ$RD�k�{}��v��}���~��r�����+�n�X�����q�H3�.���Uw��燵5�r�fL˼�n�+`Ȥ�߻���$S��{zRE$Nv���~F�!�E>���zRE$O�~���W)��.VfK���)�w���@���߫�}c���v�߯JH�������
�}���
�V\�����/JH��߫�}k���r��ޔ��?Dd� }��~��"��߿^��I�=;'J�ea/!yRkY��$>�����RE$N�߾��)"�W{�Ғ	�?+hP�~pPT@	t4������lw�NT�����ə�U^w�RE$Nw��qI�H~��Da��y�?~��~,�}�(���ܝ���zB;Bۧ�E���9X��BѲ��\3�������;�7����o���1������H����^��I��w�;�H�9��C�	���߻��{"�)_Y>��.L��*K�/JH����;���QN��kJH��߻���$S��{z��BTD�߾���&���V�����X�) ��}�߷�$RD������E'���Ғ)"w���X�)"�zN��]UVd̻����JH/��w����qI�s�JH����;�]�$�~�]��Ғ)"|s��>��T�3%fd����)"�����$RC� �D�>�_~�c�E?}��iI�9�w��$S8���_��]5��věl UUR�v1�=��\��qa�ݶ�A9Am�R��Gݰ��Z��}��  ���\iM���E�v}z�lF�6�����4$���,�T^�2�g��.���K��v�;\ݹfy�A�uӍ�!�B;c�:ƫ]; ��m`� h7U�v[v��m�w;gQg�1�dǍ=v��
bl��d�����{����|>u���Z���]cV��;>����|I.��[�[V��m�;wѻ麊�wU�d���)"�'߫�~��RE;\�oJH��������O��٥$RD������V1��5�Վ�)��;z� �?$$R�2'߾��C���O���4��H�;\�lw� TSڟ|Y�wYy30ʫ�32���H���}��RE'}�sJH�@HAj'~�����)�w�^��IӼ���.�2��1�����)"���iI�9��{�;�H�k���I > ϻ���$S�Y>��.L��*\���)"�';\�lw�G�
b���zRE$N�߾��)"�����$RG���v�~o��~T�"rK7<��*��A���}7+q�n;%m�b�N]v�7|�������nP*����d�3�/ye�o3V>�$S���ޔ�I��{��RE'}�sJ(|*) ����X�)"��O�.��2]e�cW�zRE$Nw��p�"���� �i �X(0�E'����$RD����c������ޔ� @C�T�'�O�~��T�3%fd����)"��~�D�����9������߯JH��߹���dS��P��U.�I�.�4��~@�#P$N�]���$S��~�)"�';��C������{�E$N���:T�+	��T��j�qI�s��)"�
A������ؤ�O��s@Ȥ���;��$}��~#�'F��ֆ�6q��L�f�զ�Rd��Mv���TODPc�{�����E�	��U^���$RD�y��w�I�{�Ғ)"s�����RE;\�oJH����v����w�WY&7�W�"�	쯯�@|j)"w���X�)"�W{��I�y�w��dS�t����.�¥ˬ�Ғ)"s����qI�s��)#��ը!H# ����x�=[J$b�H� ���z�E��wZ��;�H���iI�;�{]���¦aZ�f^V�5c��� ���}������}��ߴ;�H���}�RA>D?��O�W߿X�)"���~���U�.���/JH������) ���}�RE$�W~��p|�QN�3��$RD�'�r����]\��fs�N��*�v�N�����J䓰�ך��/�z�3/*P�b6f���\��d���2]fh|�H���}�RE$Nv����)"��s��_��! H�QI�w�;�H�ܝ1����fK�ʻ��)"�';\�lw�,1D )�����ץ$RD��߿hw�I�{�ҟ�!� �1@�qI��O�~*e���o*Mk5c�������zRE$Nw��pO�"�X��J��f��}�Q;�g�X�)"�T�K�uw��3��33/JH��@#�w����qI�s�JH����;��$wh����{�Ғ) ﳝ��e�f^VI����qI����)"���1{�w�|�H����zRE$Nw���{ݷ����{���y�n8yn�NʽmTќ��a�sc��z]t�熺�n����n�xhݕ���*���ˬ�ڒ)"w���X�)"��s��$RD�y��=F'��"����Ғ)"}��W�td�9�h�����f��qI�s��|�+)J�߾���$R}߻�E$Nv����$H/�@�j)��ҵr��%�^V5y��$RD�����);�{�RG���n'߫�߬w�O��߯JH����N�ں�R�̕���3C�����`J��}�RE$N�]��]�$S��v���~����,���~���RE?v|c�����Y��%]�iI�9��{k���?@X0HbA��߯JH��߻���$Rw��4����ow��~����� ��8��h  �͹z�u�7=�.�b-v�cn���a���p �a&+v�:��6Ā  �g�0���j�
��v�v�t�[,�R��2��N΀��� ���f{p��Gv�-�u��\�4���nێ9�7d���)�2k��y�\n7��g�$+���ɑ�r ��n�䝋��"#;/Knŋ�ĕ���o�w���wwS��:;=Am��͒x%m�see�z�i��v�q
-��erV]J<�E�
B!,�rl��VYE�I�f�|�ȧ���ץ$RD�y��w�I�{��}"$F X1B ���B)"�B��'~�����)���|]]�eJɓ*���Ғ"s��t;���P�Db! 1���}�iI�;�w�w�N�9��?EV!",D��ϧ~��2�/+$����C���O��٥$R@y��{c� ���*�w�^��I�w�;�H�(���wrfxcwWY��$~H�%D��߾��RE>���Ғ)"s��t;�H���V"EJ��}�RE$O�����0�\���ֳV;�H�k���I��0"����h|�H���}�RE$Nv�מ{���<°���D�D�����"�ֶ&�� ��7e"}6�ڹu'�g�w����oFV�n�UfK���j�/JH��߻���$Rw��4��H��s��@�!�RE>���Ғ)"{�;>�꺩RVr�2]fhw�I�{�� 4�%�C ႕�5�k�w�O������H��;��'� �������U�.�U�f��I�����;�H�k���I~X�Ċ� �D�����)>��f��I�=;'J�eau�^T��j�qI~ " �H1 v}�}�Ғ)"w����qI����) )�A`� `D������;�H����uwY�0��Uxff^��I��{��RD~ ��H�_s�JH��߫�}c���v��ޔ�I=߯��{���y�n8�.�:�ɗ��V��#�m��D���E]�̙F3/
��Kɛ�re�f^V3/4>E$R}Ͼ�)"�'��w�;�H�k���U>B"TRD��}��qI����0������JH���+���� �� \S�}��Ғ)"s�߿hw�I�{��)�����{�}wFMc�V�je�kXj�qI��߯JH���;��w��0:,]��`�'����RE$O�\���qI�ӕ�Z�*�&e�^5y��$E�H5�����$R}Ͼ�)"�'��w�;�H!���߯JH����Ϩ��QR�̕����{Ȥ�N��)"���� w����b�)�����I�<�{��)ڝ�ʿ�v��4qYԵ깲��&-F٭ۧg��s"]u�d��1�;�����;羋�4]C*d��ͩ"�/;]���$S��v���H>s��qI�W}�sJH����G�r��]��&����RE;\�o@~+�`�RD�߿~��)"��~�)"���w�;�?E�����uWY�.�eUᙙzRE$O{��hw�I�{�Ғ|@j';]���$S߯�V��I��vNɗu�yXLl̼��)'�)������iI�;�}����2)�o��) �Ꙍ�0�$Z�H)E�	��|��)"��Ý����*��3JH���+���(?1k߻�h�=��}��RE'=�sJH�"z	�*v���XU����hl�Ӌm�T�]�Y��z��x�b�8)����.�*��Xj����5�aZ�����f�|�H�����RE$O9��C���N{���X�b����G0� 9��Oh&nȻ������Ғ) �����>`�@ �ȍE'y߳JH����~��qI�w��"��b�*) ��g�}W(�XfJ��^f�qI��~�)"�'9\�lw�I�y��2)"y����$S�Θ����U�2�J��Ғ� �B�w�߾��RE'�w�����'��RAS�@*��w�Ғ)"w�H��T��嗔M^�c���O;�攑I�O�@^�����ؤ�O����2)"s����qI���}�o��a֊>��������*��wY{���!,�0�.���� ĳF����@��

�%�.��*�۲�1�]���<��{;]�?�in�����M#!a�
J�g�R@�%0�nou*����aE׉��!�F�$K`6]�*�$@�bݚ$# �68!�.6�x�@.V�L�͊m��)h��)�a����3�. f	g�c37��;�$�I$  	� 6�     H�m  6��                ?H> P�6� �������mE6l�k�ק,�U�k�rM�Q�KU,�Z��[�j�yư�<i����JP��4v1c���=��\��f����s� � d ��-��@A����� �  �J�    �� )Ii� `8 p��m�M��  �  @  �               � p [@��m���JIq��������n��@�� $%[Fݤg��@2�V�f���vyi�[&���4�u�a⹸�rڥ���6؃�> �@
P`8�jg]��b5�h��Qͥt {gqm�;�1�����ᗕJZڥ�/Zd�Z\�z�]m �I���ī-v�a
7#uN��m5V��e�
�� X`��^��ڍ#L�RU\��pn��&����â������٭�F���f6��{+��ҽq.�[s�i@�HD��
�N]�qE���l�K�/<� ��z��z��y�W��Rs�9�^��alPB�cD[���͕��u�l�Y˽l�u�l�-g�;B�>c6M���1zڢ1�(\�{P\8ڲn��^zԌ��[b��	����|��{s�?8W�ڪʴ�$E�kV����
b��qS���;Z����w����@ઋ��,��GS�����U�d���϶�y-������N�.�Z�g��$�m�n0�7W��j��[dcp�B [v�7C\uu���lN�v��&�6P����黓E��/4��:�;�6V9^��U�Z��\۴�Ja�r<��0�T9bsk�(�n)%l�v+f�.���|�v
�\�[U�������w=��w����B��<`�����~�&����������w������ V��
�  m���e�K~��*Ѷ���k��t� 
J`�kh`�T��v�Զ�   UT��(p6�X�xn�=�L���p!!,�M{1��
�7	��Nzvs��JL�����l]�qמ�v\N6�c[.88���l�G���;`����CrR1�R<\�bk9�)�f��'d���l��C��κ�W8���w��tl�R���f�p[l
/3I��j�>�7�>����]i�;����l���uWY���Uy�Y��$RD���~��)"���$RA�+��D<�H�����RE$O{;��I�u�yXeB����)9�;��EO��H�}_�~��E'?}�4��H����qI���w&aW�7uu��RE$Nr����Ĩ��攐�Q9���C���O��٥$RD��v�0�\���Z��X�) <�;�E$O{�wC���N{�攑 �9��{V;�H�������UfL˼�++34�H����qI>�]�~�)"�'{_w��$Ry�w4��C��_�?$��F�co��8H��b��+Y(�Y�-�/�nke�-;�{f�����;��XfJ�˕Y�"�);���RE$cvV��a�@s�|�_b"	m<���XQS.ꌩ���5$�/����G�W��0R�!rI�`2(k2�*�A�4�-%��Lh��� r�/H����
�Ϸ����� o�_b92j�q.\ėW1W0m^V�sn�m=�">rw�%]k��.4ڑ
LPq�$�y�������*��Bf>���N�G0�R8�Ic���@7��3nϒ��=䮻!�Z� |���:���o������%6S���k�PYu�Xe*�b㉶}u�N%��w�����>\���u����ku��W�>KV>DD�DG���@^N]Tř|���.���k =��G���y��@�����n�t)��7$�㓀{n��>����-�R�HO�`��1��RQ�$dF2H2$#��d!$$	!A��P%��߼��	�}�jp��;;W(�X\��&for~(S��0�~�I9����^��{�ԛ"H�@/߾�F����ՅT2�ʙwuyz�{���ԓ�O�	 #ȭ��y�߳ ��*��鍩�s��wY��5���\'f��&�A������v�,s��c�8�d�y9�X��8��} ���ԓ�����׽��O��AbԐ;��ߟ@�?~��mH�$9$rpm��"#�� �Hn�}*�� =䯱��30���A�7�~ڑ����ށ���B�����#�$7[���i� fe3sl��I��$mH���<��8DSt����~���j�
��1�	V����`�Eb�L��7����6��I���99����s~D��A�O~����v����s��:�m���r�I�E�&�pښ%t��U�s���k�6�5j�A�v]���j��q;�Q�ԓ�N`������@տ�>������9��u��
=��4LI7s7w����U��G9 �l'X���Um�L���7'�LHȚ2"$�|���@;���5��@��� O����Q��q�3<=�g �{�5}��<��0�m}ܷ%ƛR!I�uSwx���D)�� J�:�n������ϳ7�F�I�7�rm�  �m�I��q=8#�ONExڪ���6����@۶ж�  ~`�F��٫i%r֬Q��Y�j�[d::��9۠j��*l�I4Y'[���F�{]1%�]��ٚ������ 1�rm�<q�aMN{�r��
㜜���"�gn��M�Ex;\��	���.�I�:�v������{�{�v���:3�Z<�v��U�E8�z,�+yj��<�N�Ć�mH�h�Ǒ��@��π%\�h�w��� ki��
�����<m�#������l��=��u�/'.�bͿ��g0����+ >Z��bZ�܈��H�S���jo�{����H�jI�)'��ö����u���u�}�ǚw�(�*b�FH��	'z���<��v}����p۷�߁�Ӳ?x�d�y�öZ�ƨ1�����g:.�h$9��d�y�1#&6ddI����k�4�m=���O'X|7��S.��D�kW�$��k��� X܈.,Ř�J��{Uc�'�'�����ԉ)1��ԓ����_�������%\�o�BZw�{�G0auSwW0�Ǒ�ޘ~��^�πZ��} ���0�{�>Y��cl$��O�R> �ru�}�FO�w�y�{�)�� ���}��J���Y��嬓�/]�ʷ�rspll��3֨�W]��ݔ���W�3�//2��;�5��@S��G�G�Fx#^�Ϡ}�_��`��F����jI����� R	�@s��߯D�ﯿ~} ���u����ɋ"RL$����ݽI'9^�Jn,�h���2� �t��P?�u=��Nv����ryTČ�k#"M����s��9��J�)�����_@�$� ��u��>o똛��������4� ""8�"8B�O� �S���^�X��~.�#���+�s��͜G��l�YqD��f
����@c�'4Pc�������w˾���ԉ)1��ԓ�~����z����j�܎} y�}��.�nl��䊒�� ����G9����s�� y�}$��w�Ȕ	S�t��w&aYr�uwX�I�� �N���
y:�;֪ڀvy"\ᑓ��}��۶p����$�{�ޤ��"xШX��9_@��R5�b�I�7۷��N�u�րy�x{��S������zt�T�;h'X�N�ڥs���1�����,��u���O���hZ�~ )�� �\�o�BZw� ���p�e0Y�FD���}_־��<��4�-i���U��� �ա��s
&�xE�d�����p���@����>��_@�<�%ƛR$��RN�՘m{U`U�V�DO'�;�����P�Ɖ'z����Zn� �N��%�DW9��w��9�߮��~~T��lpV��_*�T  m����iӷ4�Y�gN^6���kjC�(pm��0�ā�l���6Ā6� H�ۋ��L���qz�F�\�� ���u[�V�A�ŷY7�y�{N�i� �#HKzNs��rIz�'�n'�2�psF- %��Px�&6�,5ub:�r�X�sm���$�4X���wc�tf�8�SW=�����wy��>T��2��-�I�W���3�mћW=H��lWR��x����<�L���I�0�R>����} ��sot<�`�˪�o�s�/�}� �j���"��<��u�>��_����x��m���I1Ewx5���O'X:��@sҝ�A���J���%$����̯o��5ַX��}�"V�� Z8�a7�1���7 3>��_@�۶p���@����=�ͫZv5�`�D�
2�6I���U͕�5l%do<:v�$��W<,�J��bL<�<�M���I��n��7�0�j���[�Т�	�����/%��ff�U9�{����"m`��"X��!�2��^�';}�or�l�wO�P��P�ƈ�z�j���KUa�G�w������cl$�1��jD�їl����7V��q*�:����M��˲{�.�ʼ�4� I���N� �M���VݍIO��NFFJ�Z�k����_�-l��,�m��ѭ����X���q�I�)'@����������_���8����"RH';�6y:��6�@<Ӽ&����b�Y1A7X}]��۶p�s��y=5~R>a��P!��5)i(��4�R��t�6FJID���#ES��t��TU����
BS)eABM!("H ;ҁ^ �qaj�H$HsHl��Oh�@$�#��a%�dI"0�n�$H!FT�!QP�y�`Q#�	o!��*�˷d<�h	D����BS*H�#.RJ�P����)�**RP��JؽNh�� <^�<8���W�N&�T9��S��\���"���o4�Fs�P҉#U����{ܐ�w��I=���\������.`ʾ��G93���y�FϵW@�	V�lV�����9�mI8�05}����_@=�g0}
f�dY�x��㘱Ljv��!m��L�nڠ^l&�:*��Y�h�Nt�ʐU7use�%�� 㐫S�]ku�-V�2AkO0�P��U�M\_*���u�րy�x��
y:��,�[����j��As�I�\Rq�@>��^�{�R�N�t��܉ee �l�b�I�7뷽W�_ ��������̂�z`����PUJ�K��h ���yEZ�4��[)�߉�.��D��C�l��ys5$��}>��T˙�7wd����4�4�;�{{�>�*6ݍa�H�HN%�A�Ij�l���Z��n�T��Ovq%���3�[e�cY1�7 ����۶p۷���V�ρ�?~�,Q7��N>�y%}s"֞NL�N��jU�}h&Ԋ')RN~�<K����
��� �����n����
�#�˒*K��O'X:��@<Ӽ��߮����f���	152y#jG�>��� �N��=��u�w���"b	� B��,U���Oj�w��s{���� ��<V�UU@ �6��,��k�:�)4lC2��*��
�Ym&�9�$HCu�Զ�b@  Eg��i=�T���nt�^��A�崒G�'ͧټ[@ �&�<��&��C�ۣ�:��\-�>+��N���qd�(x:�s��fq�]�Q�*�v���;s�d.֦i���B��u��綗�I[\$V+א����[|W���u���N-�ES��K>�y+=/�8+`R^+0�s���t|�|m@9<�\��q���s����@�����d�����DDǵ��K�6I1E$�_��癁��}_־�{v�?3�΂��1���)S"2I���n�@R���su�i� ��ށ�&PS�cY1�7<������<ӼsOt S��˃����������n��;���\���k�g�}k��ڳ�I��<q9��\����vi<�V�}lgt>��t<�ZqC�LrmH�&8ڒp���@��u�s�n��4� �sU7usfT.�^od���;z(��R���1`��! l�6�$
��$`đ�`BH�YB�u=hw9����$�{�検���c|��L8}���������T��@�Z�h�w�����
y:�;�˪�/�d�:]�۾����r�E4�-i��j�U�>��_@��W�q�%#���&����=�!O'X:��@<Ӝ�~(�cv4cx�M�bp���(�����u�[Fлnk#�=%Ӻ�j�pl�p���)$�������k�{v��]���re0X�117 �*�U�ܪ	i�@Z�� 6}�����E≸�E�d���l���ޏ��2�q\���٩';}�op�Å�&Ԉ�aRN�v��j�k���k�~K��������P��j*��6}���':�|��[�0�\���0<�2��m������NHJl
�WJ�Z�{qx�1�3<.�\�]�8�:9䑶bjd�Fԏ�;_���nف����l��N����M����9�]��yZ��|&��O'Xu������f�.0#��LQI8�՘�*�� #�ηX��}c�
TČP$$�Iށ��f������orI�y�ԑ�#yIR"ÿv~��~�����Ʋc�9 ���h6��	��@n��0�SN�i�γ3�kC���(��j4�۰��v�)<q�x���-�ގ!b�;?W��l6��	��@n����۝LjDG0���'���׵p�KW@-�8t��ڑŒ5���� O���Ӽ4��1��6�LML�H6��~�3W��ߗ@N��՘U�z�����2�vNae�^N�6��i<�)�NtvZ���\��#m$��Ӑ  ��i�޷�"��]�l�55t۬� 
����86�8��6�Զ�   �6��0r�6�:�t���N�k��@
S���4kovn8�-N�B�q\��E����t��jJ�B�X댑nn�g���9�>r�ڭ�^Q�v���&�V��l��v�T;K�c�k��l�,l���[u�OI��juqv���V4ZM�/4㇖�Wik�F�Ʉ�7U�8ۢ�\���h{v��$����&(���v��@��\k���v����J�Id��$�);�-{W�e_[��[_ �����ߋ�()���b�9 ���x���@/�V`~�9ݧ=-7ȑ�"";'9:Uv�}ݽ�����3����@���	�"#�A�SwX�Otn��ϒw�9i������W�N����zB;B۪����z9���ct��X�Vw<��ی��JSH�Nw�Z�� S��:Wl�����@՗-���S'���^s���J���m���v�$�9��p-{W?ffx�����n0��H.C$�����N�ԅ�8�7I�@s���/٪��(�$�ԏ�]�{�-{W ��l�Uv�st4���F8�$$�����U��t
���.��f}�[v91���A���ӶQ��54h%�s�:�ҧ]CҘ��fw�p�9�0X�LR'"�}m�����oz�j�߃�|�n(w�z��`&�@n���6�a�,�{A6�Ds"�R>wm�����ԽJP!d	�)1�Wk�k��>V��=���#�&O��V��
|��J�]-&��6aBwM��� dcn.U�g@��|ݷ�����y���+RH�k��q��Y'`^�1�x�x�Nc�$n}u�+��f�m���D��2I�9��*�k���}��
��:ܪ��H����n�>6����u��J����\�T��$��w�P�:����y:�M���&����b�n����X�w�9��%��{��*�bA��]���RO9����ʫ��*����Ut���;>W���7�;Ȱp��D�������M�+.(�Z6�Mq2�8�M��e�b�#��R"9�(�|��ށW�_ ��l��=��{M�*#jGH�T�W��j��L�u�x�N�ݷ�四cl$�9��Ĥ|����7I� �ot-:�=���]�I!���'#�'@��\��ށU��_[g@��Qq���I2&��u,�s��u�9���	V�����l��RO}�n�(��j�h�b9�(H
�"B
�,)�0��JQ���	X�����,���� 
�&n� B*�cHv�(FE�D�Mn}�2��J�wI�|    � m�p    p [@  �                   0`l �RY.;-�LRԭV�72po]\��mR����/a��wQ׶l�����ti���I��ۖ�u��s/��T�O38�����  (0 8�4P8 p (k@  �J �    �g 2 R���  p �Am�����    � H   ��    m�        �  �8mqf�]��lk]�-�6�WU��m� -�l����K+fܕ�K��ږɂ�F��n�Ul'n|�U���)ѫm���2 �g  d �� X��9�B��ژ�I�T܌��]��Ha9����-�n�cQ����pd���M��ɶ�� m[Q�brަ6�m&��mmi6-��Y�� izD�V�$�� j��2���"3'�m�+5��5�+%U;����;&�q����6��n̒ƞwɚ��u��.9�6������ma�N�泭`��t��a��\�A:�FC��:^Ҝu�K`]�IT����M�����OJ�#>{g�u��5J� -¢3�+�`6�[��g����^������݋��v�Tmջۋn�^Hγ�͈� ��pk,��NӲ��N��e���RR5�u��V��[�����i8�;��8K�'.�n��'�I�t67N�J�%�ӡ��������/�ֺ6�g�d�GF�,�s�+VJ���-�[�x��Yy�/#%��2G`7j�<3�:�QS^^
��x�s�\����&�k!��פ.�|��j�ܺbs��F݋�zGl��ڡ���h��&�ZH-:��S9���[�R �&Uٮ�����L�ˡ�p㊆����{�< �m��eZ�xX��<E��yG.��W.��0�nؓm�  �[��8��N8���JN�Jr�[[hd��Hv���i�  6[%q�^��Z����t�5�m� ���9���l�J��3h���m����N{WA�+�Q���ΖnrQZ�7o#�r�9��\v�����C�v��=�/Q��y�u#���Y����lcƫn��
bl��d���{�m+�n��δ6y�ӶES�m�(��P��vQdHθ�Qۈ�2η�D]��e�5���� r�w�7I� �otE��S�PLR8��m�t^��.�{�*�_?������Ad�F]���7I�@Z�,��W�ꄯ�}���R(� �ģ���3�1~��� �}N��LʭS�>F�
KmH�B���l��<�Ŀ+~�]'=y%��2K����������[����Z*��]��6N���c��euaU��9�dǒ4�1�������9�s�>M�.n�#�n�U�eę��d�֦k5��{��kV�B�c)	 ��z�%[*�"�D(�ǽ�w@97x�Mށ��1���I2&��� ߭�����>�j��6�4�F8�$$���.n�<���'8�����ʦ��b���p
��g@����_����l�v��k&,y �q�y��[u]\�������뎧�P�7=L�J�؄I�A��Dvs�����~������U�l�e�h&Ԉ�yU��\��c�DL���9I��=^��>���#�&O���lԓ��w��^ؼBB,`/��0�+��n��@�gٹcM��!<�W}.�n�t���`�+�{k�����$�����W�p�`�+�
wR��"9�����u7P���6y�ӶES�v�gÿ��?,<Z2ٷ/Y�����fn�y�N��-t,|������W��x�j���CJ�B"Ds$Rw�����1#��������u,�=��⛂y7D������@S��U�z>re��`������ɋ*�l.M�̽�'8��{��'=�sRy�����/�Ij��b�<���}��z|_>���2�^E�U��\�&�@7x�mށζ��3�?fЦ~jH����1b�˶l�Re�ۚ����s�������v���DFԎ,�<i'=���ӀU��t�ڸݷ� ��>��mD�	�h���$� �S��9și7� �~\�n��aو�\�I9�NN��{W@[�fdZ��s$�n�P�I��HD��qp�oz�[8_[gO�U�\��T�"9"�tsw�9����9�M�?}�C�H��2W{�U%ffITQ&�   �mνRN�nx��tE��+[[���a���p �Ă�j㭭�lH  m�7m�U�u-��çm�n�iҹl�AJXA��m��5��J�����I��s/]@Xă���՜*�w^+�����u�f쎞���n���p���=mD��<nqL��#Û�n�m�e���^1�tX�V^^U�L*B�2ͣ�C�7S{�w{���D8��jZ��+-c�c�N����'�7\tҵ�ݹ�1�<�.ǉ�\BU��r�;�<�T���r0|�����$R4DL����W�s����߻���NW���>ˎ�M�ȼq'W8I������.y��:y:�=��Ɔ�6�ƒ|�}ݜW��tO�WA�9��`0�C������]Iuw�9���<�`&�@=��m�??f�W�K���͞zqm�*��%���l\M6�k#vx�B�7<�,��x���U�w��tO'XI��sw�9�l�nZ��	"D�#R>wm�y ^�<��YRs��ԓ��{�ܓ������hS�i�q���_o�נ9\��<�`&�@\8���Ɋ1d���U��t��_ �����l����|��7#B�����j��ަ�����>ԯ |�G�ߟþ���|��qr[l
/)٤!v�D+�tn`Ϯ�[��e������5��[�nnn� z�� ��_@S�J�O�W@��nЍ��JdD$JN�߭����Sw�l�u��,�=1�����nf������� sɻ�:y:�Ǡ��>����H��4BPE��1a	HB�(Z-�5x��F1�"�u������#Uη}�j�U�e�n��.����o��ju���D϶��"]{S�T7Ru��B%$�Ԙ�����[8^��t��_ ��T�ݍ��4�s6�̱E͕���֫9����n��ؙuӺ{5]� dM!"9"�� ��g �ߵ^���|����O0��㛘�n�����n� s�N��N��Ot�[9�8���g��Ad��DuI�s�T���7ܞ���������6MH��Ŏ(�|����߭��~����@hPn��v�$�g��wYWs7%�s7y�y
��9,��V�π_~�ށ~Ҷ������N=!)�*���V�ѫv5聸�f{pmqOg4�K��<�#M��QO#Drp
��l�/�W@_{V>r"#"#�����*uWA�7eg�wyYyzO'Q�?r{��� �߶΁��xc	��$R> �������s.}�����@Q�*i�q����[8^��tO�WA�9��� hؾ9��&蘸��&�������֧X�������m������ V��
��� �m�Yzލu������КL��� ]�(m�����5�7�gR۶m�   -��k�8
��,��;l�p]UUWP-�@�˝���^���'�I��$��݄�8�1�7n�Z�����ή]�n���؍��<�p.̤�s۳���t�l�9��b;���א�h�%w	.�;��k��E�/6{�����̓�~G���Y��5����GC��Z�˻m����sGo�-���-��U]ԓrl���<�`ܞ����*��}����R"71c�)+ ��Ov����7x�Bw�t�u�v�mڎD�DBD��@=��p
��ށ��� ����
;��������������������� �7x�ҝ]i�ݕ�]��e��<�`�j� ��_@S��^ �,s4U;�s��&�p��J�v�n�Kj����5[/b�7/"jv�5{];gf��)�����������n��N��J�B"$qĤ�@=���s�<���Q���l�,������_�<���y�E�Q�&,���
������%�S���S���U�3��E�SWe�ܛ7�zO'X�OtO7X�ss�}���R"78�����{�=<�`}�ށ��� ��uT�.J��6y��nk�&.�p�Z��V�\��xX���ғAtkPW����~۬Ϲ��:y:�r{�t�i��QO#�|�~�t��_ �}����[���l�WAXrn��.��]�o@��� }��l\MT�}�D�B�
֬%�.�l�H���1X�H�k ��]l�T��P�$��@R����,!z�"��l�cCP�Y@L�Uˢ]؎)��ҧ�,�h����4�!�-�(�҄�lg��Jղ��D�d	 � � HH�H$�H$��vd����I#(�==v�[��7G�~8�d�-X
�]��X��
f�);��"@^���+&����=耜 �pC|�R"$�_ShqN"��7��N�k[�I=�;��F��J�ǀ0s"�I��_~�ށ��� s�n��;�{��jd�䫉�������� ����rw����|4VݎF�?c�G�R����9{u��@�jsč����t�y�LI7\MTT�� ����rw�>���=_Z�~�3r�YrGT�'@��Uu󜉑�y�zu��
~�W�d�?c��jE�$QH���������U��΁��k���B6��)����� �7x�sw�ʙ���>0հ
�gw�䜣�N���eT̘��uw�9�7zܝ��=�sw��_�����*��NIf㇖�Nʽv�c9{uخG[������k��]v�7l����Y����Vf^�w'x�Ot�����{���l���rc�I�ԫ�op��W@S����{U�̎5��Y�(�N�����^�l��m�������O*��17�H�^��B�C��'����{�2ɋ����nL��o =�W�G8�S��=:�t?y+�&9�s�`���UL�$m�6�  ٲ�l25�v)AX��l��� i�m��pm�p�d�ami�  6N�W[%s��t��������j��q�Hu�f���7(���E� 䥲V�Mؚ��5���kPU�Dc+��;س�(t�ݼ�lkU�xI��&8 ���0�m��b5H�������[x����d5V����q�������w����;Y��t6y�����M�+.(�76n��v�s��6�,��A�=�m�(�+j�������� s�n�G�z}2$�^����F�r%2#��;�=_Z��se�<�`ܞ�0�C�����쿮�n��>��@��� }���䫠����S����Mŕ�]���������r{�zy������Q�rd�G�>�������j��:��{���5�c���d"s<���"��\D���=OK�r���cF6��TmS��"i%�b�'�@�}k���ށ����'�������$��.&�̽I9^����*`hіKH4D�bb# �N������U�2}�(�s���LqS����p��{�=_Z�^�l�yq�	�"�HF���OtO7X�sw����s�QȔȌ�5'z��_ �߭� ��_��ހzS5�$y�<x�q�p�l�!MFWm�Փ� 68�/��/b��f5�H�j$HL�8��~o�Ӡ	?׀>��@��X�But��vWyww��{x�j��s��A�_��*��gy�������dQɎ+��?$�n����QD.Sͽ ��p�����D9�9"��ٙ���)��x�ګ�|��0�|�,B�d��5#�����>_m|����W�k�m�;ȁ��<�ԭ��l����m�l�<�w#�L��Rc��"���s&8���N���k�߶��z���_[g@�ˎ�M�J@�����9��@��u�mށ�ʾ�7hF�r%2#$QIށ�����n��N�i��:aB�u5Ss%�qeAuu�)���rw�sM��oP*(����>��$��v���K�s뻼̼� �N�i��=<�`��΁�>
ۨh�F�D���t�T�q��3��b-�k������3vg5��N�Ùrc�I�7������+���΀o�g ����4�ȇ1G$Rw�{<�`
y�zܝ��{����C����x�Hm�5}m� ��p�g�y�_]����ߟ ��U��!1�vs��ܝ��{�zy��r�[w�w���R(��Ɯ|���z���<۽���r3��ό����fh�X��H�$bJ!)Y���~qt���%�I6�   m��M�oo^x�k�9x�,��IR0h����� G݈[[-8m����rI]xѨ��O%�ݵ����5��T�.�V���5�a	J�=p��٫�^0���:y��j��\i|3ɋ���	tR�qI�ZG�ݘ�6�k�&�\�0�b�ۜY�n���I��-]:�*^��%�Y�9ߝ����'�;���3q��m�([dj�+�nk�k�����y4�ֻLݜVғAth�����t�u�)���<�`i��,�ܱ��H���q�_m��z}���R���U��G&O�a�.�p�n����2�/@R���<�{�zy��5}�΁�Ҷq��̊92E#�~ȎDr|�`�n�ϵ+�=>�]F�iSI,����E'z���|����*�����m�۶��j6����� a���v������n�5֫m�:��g��D4y�I�C��X�0ɉ�jG�5}�΀w'x�otO7X�&�1u3XayR����I=���i0">��,��f����o�R�|�r9ɓx�0M�I�Hԓ�}�������|~{k��m��nЍ��JA,�E'p��W@|��������|�,�=9��cM��!2����_C�ګ�|�,�>�%]�c��u7SwS����N-�ES��K=e�8��T[h�u��W<uj$F6�8��zx�8w��'_8�����R���T�AN�� ��Tv�`�E�"��n����H�o�πU���=>�]q�D�� C�����������0N�w�6}�^_G#���9E��҈�\��oRM����$糬�
a�xԏ�j��:��}v��W־߾.,�#I�#�������u�kM���� Sͻ�=��{~���b���n8�-������v"筰Q�z�r��{j⇷�n��
��nn� ֛���U�6|����}M���H%�(��@�}k��N�� ���yjY�zcca]MT��v\YP]]`
y�zܩ�4���n���	��2"��3//@�V��otO7X�興�À�����C^k[�nI�;;w5d.K�+/0��΁�f ���� S���=�wm���7�9$��ylpڗ2�]�lMt�56�y�V�XvZr�Wn�KS	$�N�W־��l���U�>�oz��'�E�S��Ƥ|W���=�ـsM���� ���Û&.�j�*�����=�ـsM���� ���t���PiȢNbr����� ��w[!�V�X����)�E�������l������f8�;c`��O9��1�:�J%��H]S��(�.��!Q���,��E�
���G0�Y5a�T��U��,��H���aI��̠��C�(^!!�L��R1�1$�$a!J���*of�����f�H�B�H)B�}]�Z :��T$�a$�h*��I�T2��^�@$b B��uRvFV��p��!-�J DH�da�3��甄���@��,����0�RU&z�>!+{��~J	L�1!�۷�x���Ƿw�a�UUUU@ /Z  �    h   [@                  8  l �lN���]�\�l�]9K���W=m�mP D�εuyz����B�d�UG���d�F�8�h9��s0��2�SU<�l�h2N�:\ �����"���@
P`8 pm� H)@A�����$    ���Jр �J-��-[\  8 � �  m     �         h  h��UҒW"A��Y�7 �i6β�[vͶ
P4�#�h�:�MysI�pV����b4� p=�U���Ye�� @�A�m�J  d �4uU�j�)՚fךƺ�@�8�d^���n������\lF5�z|�Wj^�ɡm�����Y���J�C�9�٥b���.�m�#l�[�m&����[d�k�����d 5m�]f�����������kae@(Ʋ��c�1���#=n ��ue.pv�F�4 Ϯݱ�zq�Ҽ�/��
q�t�{=���Ě���v\g��Zi��X��w����sל�M3���;(��sUʀK�l�n��S�kX�l.��ok�l&�7un(��s�۞����#��=��\�FNCo&,��V6lr;mZ��V0]�\[:��Ż �m$(-��=���R��K]��^VTV��j��u�N�Z�b�P9s6ېء���ws��>@;4m�\�Ƨ�pN�k���u�l��h�;&��=��%����)��*��z�7'A��.I�v'���i�v�VR"=p;�iηN��Z�	�Y�J��:�ƶUՔF�cT- ��B\	nӡI��@<܇9+*���r]�fffeUeLɔg�3�
�CBiU���z�� �C��� �]X�3�W��UUU�Io�%�   m�m��n��m�\�DsUC0�mV7 Vj�i7 0a��L�볩6�l�   [v�֬٬�jA���- �b��6�SU]c��QÓEtl��{&�uj\[�ێ��!V�=�Wg���:�T��\�öζ�����\uҜ����7X-�=���$뮅���ʎ���֘��飥�	�k��5�~���v�w���|V���kCg����#��%Z���H7M`��GX�9��]ώy�H��ˋ*���sw�{�� �������t��vg�Uy�yz�[0i��=<�`	�n�LuFV�̊9<�C�m�{�=_m|;�y�%�������nj�I,����I����� �&�@�+f}�Ji�h�_'�E�S��Ƥ|k�_@~}��0^K0�ګ�8�9�D|�fM#�y�����VlC��n�N�nyKe�i�捘���:,t�[1�����ڭ�V����T�9�z9s�0��?~}s�?��r%p����;������U�D�*jOk����_�_C�߷����ڎD��\�����UtU�V�}���M� eϲ֛P^HL��8�׶�����5jY������:�D}��t��vg�Uu�yZ�[0�{�z~��׶���2�'$~17�(�a��Q+���H7{%�]v�m�n�ع�T�m�od6��`�E�G!�6�����ݳe@���sPmIdmL%�������0�7Z�[0�{�/��yTX�0ɉ�jG�6���}[
z[���<�s��r,M?� �Z�g��{XJ2�2���j�'�"׼��Z��o0�ګ�j�J�(�*j�f6�"	"�v��W�_ ���Ӊ{�ڸٟ�m��D<�,�NGh-�sŵk����EV�c�M�&7=Upv2�QȔ�Y2(��@�}���m}ߞ��6����㭧��<%]tU�V8�DG92{i9�	�� �|�`��t��vg�Uu�yZ���V��8���u���`�*��AW5W|��������`�N�����&��j+� �C|���P�~-$�F��I"������?fffBv�����s�5jY�{�I�T���o�:��y��v��Q�:����K�w%�����uŬ#�3?'�E�S��Ƥ|k�k@�Rs�&�������n	������/;}��V�눉�4�`�M��m}뎅��F�$A$\V����U���t���I�@�nЍ��J@D�);���f/��π_ηXޭS�r�o� �:��'�w%��� �&�@�Rs�&����}���~w���g�� [���U@ ��i�޷�p�̸���fںm�^��%0m���p	87nKn�ے   P�Q�^[�T��V�q�$�V:�ۀ	��5�ՁqmkJ�vӍHz3+�/U.6���ɬ<�M��Fۆ6&�g�N#��jGn��s��O�5��uۦ���s�����/h9� �)��:z=$ؤ�p�N� ���آE����̰��.��n8yk$�+�e2�n+�� ���.��PJ��%�20^�)xۘ��9:����-K0�ګ�9�	�n�P�I��s"nO$�p�oz��nW�Y�=��\���g�$~�)S	$�^�)��:P�i�}�L�Rs�.m�~/�ʢ�)�LM�R>�{k��Z��o�Y�㜟V�]��S7w%\^��h�Npͽ�=<�`����֝�dX8A@"px��x��ee�y��v��j�;�S�0���n]�4�J6�"	"�g��b����z�o��>�m}ߞ��6��#j9�"33{�y^�>���D�	,�[�_���!��`�R���O vU#,���"�]��@�D��Q;/w�^�{}�jI�[{���$U�����p^9��|]&� �ժz>Dreko0N�u�3}�t��vg�Uu�yZ�� k������9�i��5Cu'h
��.j�����sotO'X:Mց�������������zt�T�Kr�N��h�x`�f ۫��3;��f�4��we����� �I��=Ԝ��oz��O*��17�H���L��Nz��`O�Wn"dͅ�7�ܗw%\^��h�9�6�L�G�آ�1 ���W\���Ԓ��������?�iȔm�DE��rV���=:�t*ԫ �ժz��B"I�<R2Iށ��k�^���=��_������Y#�I���a��ݲHt�4�]��VNc�ciݥ��Z�ئƲc�N��E���^���=S��X���}!���|���'Nd�wu��j�$���k^ )��#�����>�N��n�@�ѻRv��*���ws�5�� �}��8�D�T����������B#&�I;�=�y�ԓ��w��'��;5&΢X�E�[�z�|�U!9�&� ����=Ԝ��{�zy:�:!uT�:6{7fg�l�jV�W6V[�يRۊ��g&p��K+����}c�uF�����=Ԝ��{�zy:���h�ܠ�R%p��p�����������ߟ@��pM���L�)t]��t��R��u'8���\�.Vӂ�HG��p�m}z�9�6�@�� ���A:}7f}USy���.�� |��Γ��V������ܛd����@o��ۀ  �[�������p��K��s86��*��mm��6�8h�ݰ��Zp  �۵̒�� �5Wh�Ƶ���U�':npK�;�9��!��$��Y`�����;�G��-�M��ݚ�ld��۴k�����qۮ=�W@l��Z|n+�x�gM��;v�<�읎���]q�:�1��@d����{��*�Fb_mhl�ӧl�����|;�ܨ7�|qmu\=g�$6�3vg5�/h��L��<�E���?��׵p�m}~{W �6�S	.˻�Γ��Mր����ow�"9ɑ��|ssM�UUs���h�9�L�m��I��/��\]ܕvgo���V�s����!�I� �]���r�ܠ�R%p��pͽ�<�9���h�9�<È�O�;���3q��m�([dj�+�n��Ѵ	�m8��XΊ���ѤvՋ\�4]��I� �&�@]I� ���>�[N�2�Ɯ �����^a
D��R2�Pd@�RJ
XI!���H�T(���� ѡ����_;Z�y�y��I�� ���A:}7f}USy���.�� |��Γ��N���n���S#nO$�p�oz��\��_@ߞ��-�M�ĄF��I	'z��O@q�DC�m��-��-Գ |�wq�������* a���v���6͖s�:^�;qg�5��y�Tc���Jq�*.&�&�� s���7ժz�K0kڸw.o�L"d�N�s��o�T��K0�j����U㈈�<�0M���H��p�~�@��������,�a	�;�h�3\��Z�	�A/+˲T=@<a��I(�F�.�	F��֏	HK4#G�Q�&��yͥtP؁@(T�S�6'�9�4ބ�	{P�UE�"R�h�T�P�^���
�����:�ڸ�����r%2x�d���'8�iހ����ot��R�Ƥ\����o�j�v��kڸ�J۱���D�y�ŶȪuqԭu���h�ʴ����m���,�����.�)x�\���~{W i7��'8�mށ��L�**nʩ����p�{�y�s�9����j��4�<HDmF(�$��׵`y�z�Np�{�>�:��&<����\����o�j�v����v �E�	ZH��$J��XX�	#�*�����;�?f��L"d�N�NN��=��-Գ �V��
|��q'�'Qۛ���>a��73�������b�/=n&�f�+p��nظ��sml�-�ح�a��`U�z�$� �+G@Q�@��n��n/�wE���Z���ș�n���\����A����ͧ␏T��@s���7�h�u,�>U�z���	��3ꪜ�̽r�`+{�=�j�}m�߲���)*n���0�{�y�s�9������&���&���.I$h�x�~[��(Il��m� ��Yz�m�+y\�A���m� h����p �Ă�j㭭�lH  m�6�a�6A�A+r���n��K$�%�%�ξ;I��&P۴[�v�4k�l�%��\,�=c��\X;3.yv�n��D�Q�՞^|Ȼ݈%������8*���6d���`g3�0Qƛ�B�)2�l��u��;�����;��w���}��M�W���s,Qsek#����]�lj#<�Ų��٪��f�$"6�HI�z��\����7��~���_&2��LM�n. �w�.V����t������9�1��I��7��v���ڸ_[g@�q�PiȒ����p�{�>�� s�;�Rs�8ݡq��L�)$�@�=��U��_���Էe����)Z��)	���HF��H	J���t��PN;&Ѻ��擊�׋&�lx�<�������~~_U2/V��|�~��"#������te�[�^n�f������B����0��=O�W���A!���ƉԞI"��������y��}2�<w�.�� }*	�.�n�����#��;Nz�m���SОb����/��c+i1���&��|ӽr�`s{�y�s�oL:�q�<��fs��N�J8�4q�ۭW=��ΰ&�kز&�%���t�fq�?>��o����,�>U�_9��:Ӽ���~ڑ
&�"!�.�oz�Ꞁ��U��u�r928I���������n諼ə<�9�
|��/9�9^�>�""-R�`���>��j��n˨�������9.��x�l�u,�<�9�5t7E�N�M\g�U9u�z�l�M��I� �w�w1�����N8yj%vV�i�M�٣K��k��:rS��7�g�<���飠-�Y�|�T�>Z�� �[:�����F��I	'z��\���y�$9֝�U��-�Y�/�*��.��j�j�p<ӽr�`s{�y���wr��T�b���'9:���5���I�|�>�" �"�!0T,I|�{����ܠ�R!F� r�m�@��s�9���� �(U;��⬼u��͜Gh[u\��h��sg�D�i������q�mr�AuƣW__[o���� s�;�+f �7�9����~���**n� s�;�+f �7���\�wQ.�'3�6q���7�h�|�`�gΓ���Zw�}�)�3��	�<�C�]���kڸ^Z��G9+WY�5�&T]T�we���S��i��-V΀��g����?;�ws���� ��<V�T   �u�gV����d���$r껭� ť�� P�8�/]�Knٶ$  ��^^����j�u9n��Yӭ�8 qnΒ�n��.u	��Ӑ�c�����<Ղ���$C��N����d1��p��Y:L�7lu������q=��.��O'nsvNEg��"��'\'�v:r�����\
��s�{��w~��m�cWoh��y�;`U��u���ӌŉWJ��^'.�h��;��ۙ4�������?����_@r�� i7��j���
7�n	�*�&�r�/@|��\��t��}m�ۏr�mH���� i7��'8�mހ�[0�8mG"S"DI;�=�j�}m�}�����`8��j�����TT�� �w�$��I��<��G~��?*{�9�Y��嬓��[J1�x�b�������nk��W]���ٍ;[�w�J��̽%l�M��M���>��d?-������I��$191�wR�Q��~��"9�;'{M�@�u�x��;�d{*	�.�n���� ��)�J�|�DL�����`*\!(�
17�ȸ_[g@��Nwk���j����*�,�7	'y'/@I[0�{�y�s�9����G�N��P[hl�d�	[tٲ��O7Vn�4�G�̝g���T��r�l��ڮ��,�M��M����Q�ﺂ���\�߃�6��)��#$����=2j��Z䭘�Ot0uSW2D��QQ3W8�Iր��`�ﾉ��!�,�HG�@��]��{���������'M\v(����X��:��� �v��:I��j��<l���RC�o����}�~������@��N��c���B&�=:vȪz�-�G���.֑xJ� v��U���xA���0�BIށ�v��I:�V�y'���9��&�.
����]$�@I[0��t���s|�`�5! ��|���)�7�՘8���|�'X�V�
��Dl��� �woz�ڸkݯ���|'�Z+�4��'��#G�ة�������t�������ʬ1��.�0�%=���u�	+g@߷Va��o��i�S�y����n�$:p�&Wm�Փ�ĩ۫v�tv�����phҌ���"�f�pt��%l��{��Hy�s�>[r]�U�bʉ�o��n�&E�`t��U�� ��L�ǆ$K������@��W �{��ݔ��|Z<"6�E$*�0��s�>t��wm~�Y�_�|2�/0�7�ɋ�v�����0��t���������z9�E׷Z�t�iN��� �@�7���*�/"8��\XD���T��D�$��J,�B!4)#	�"��% �*�`Xc�؁�F"RPy���6R�U�B�j�#"���		#Dު:���HT�J�.�<M�+�m�h����$+%7U_���   h      ��� ��                  � h�l�e�M�H�-�^5@kvU)ԉƘ%�
^�v�����q�V�7a0s��,JhV�C�'A�㿻���:����F ]��5VIԒ�  )@A���>q �H0 8��6� $p �@
P`8 s� �  ���%��  mpm���,     m   m�     m�         ����rƎe�uY�� Fט@inD�� �����:[�	��PK�x��f�ں,�W�Z����5Gnj]3�bI �G 1��p �@
P`8 qp���z�+� �����ZGZl�;[�۲��ƃ,>nƧ�y��i&^jJƪZ�%-ڥ�%��-T6.��/@�@�պ]���t�m����vu�n���a�2�5�2zS���w��riN�7QYҩ������d�1ʜ*�y֑fx��x��W�Z<��z]+�Y��mN�.|�7c;�ƍ��֠��q�Q;��g[JN˟\s�=���gg`6���N����Uy�=���7L1�L�Y݌m��Me�Nzu�����^{*z[�$�zkv�R���oS��ێ5��N�I�+q�8k����Ш�҉1��-m�N�u�؞#�Z�8�W,��Hκb��˲��",t����wc�Zk�#5Tλ��N,��!�ݝm�s��Ɠ�5��n�oj�:㖝��������m�{v{��������k�7>!�HLIc�KT��[�Ώ'iݶ�Ƃ�b���ے�Up[�1)��{][��Ts;!Ke��Ԭ��Ҡ�� d���v֮]��?O�{դN�S�#h��^?�Ki��`sa∼N
�]-ml_}�5�f]�U^fI�m�d��   m��-�/mĬ��*Ň���USj4����86�8h�ݰ��   Um-��nWf� diGV��V�i A���9*C�uy,��6�����]q��`Yvڨ�OVvt]�n�bt3[nҜQnv�k����!m���Z��aD ���֮s�v�����bK ~8Cc�ȇ.K�������� ���J���:��fy��v�m�f���Qdvꌐݹʜ1��KêLx�>��	Z��?>?����/$�@�� �I:�9� �ӑ� r}ݽ��j��v�����sۡq��L�)%��M���u�$�����>o��~���N$1ȑ1' �{��݌��{�y�s�.��PN�%\dYQ=���ݴt�uf�3�M�@�տ�@��ͿѨ�o��NFG�ES�v�gû��2|qms]�OC.;f3vg5�% �n6Hcp�C�?m���@�]��v����6������ĄA�2) ��I<�������P��{��_^��s�7�ՙ��ș��C�'�dTM]�@��N�n�:��� �i)���/O��VR��&d������OU�w��j�O0������r'�i:�5�(a-��8�r}ݽ����׻_@�vS�\���jȳ���0���^f�/>�J����AJ땈�5Z��M��cj9�<R2Iށ��_ �{���eq��{��>�[N$1Ȥ�&�t���[0�OtJN���U<��N�SE�Z�K�FK+Z�^����ԓ~���s�4�B-Ah`����]����<�~�_ ��o��=�jI����nI�����I��L���ՠsw����h�!�2)19;�=[����]hJـor{�f��u0EUJ8��jZ��+9�u震$M�����]��]�{!!?��&�c��w׻_@�v��3�Վ9�D}!�I�C��l.9��!�Lb�z���>�S���H�v��@�[����k��ܡ�mH��AŃ�`ܞ���`�Iց䭘�]���Jd�I��ށ�ݯ���_'o׹'��}5&_0��(DA
��2ƀ����w$���Q���C$�&
G�;�ݯ�<���~0�S���U�DDD{�uT��jnM��zB6Ȫuqԭt�[��J*t[mf뎨�t��F���n3wεs�?��%l��j���U<�����֓�v�I><0x�!��I߾ͽ���X�M$�@�V�(8l��$���.��j�tJN��$�@�V�{��@߇pʠ�PȁɒH�}{��%l�7�=�=):���󛉒J�.������<�� ���@��� �V�}��xe��&4�9$�H�   ������t�f���xqի%H ����(m�pdq m؅��Ӏ6� H�-�]��jf�컯�%X�� �*�<���@0��^�/U�ṟ�so3+S��x{f����K�����Ɠ(:N����ղ)�.sv��hMF�m���v���K�|)��ٓ.�Q�8)��ЯZw��n���|z��b���g<���
^3�HG<��VlY�:�s�s�ۭ:��]�Ɍ&&����pq`�>���w�z�Ut��UD}!䭝G�Suw3qM�]]��I����hJـo}���y�A����C$�&
G�=��ց䭘�'��'X��\�('H��2,�����<�� ���@�wUt9�DO޴�`��f�PAQT]�Ue�ـor{;!�I��";���x����T�ݍ��4�pX�$�+\ʱ���Jع�x���q(�L���f�۱�<,Dc����������������;����oøeP^(d@��|�uVN�����w��l��y�};����o�LHC��R>�q�we:{�f�"d���$� ��Ԉ��X9߾��ն��v���� ��иڎD���&G'zөW@q�=޷��J��3�K0��ߊ���=�6�6y���6IJ���e��n[���:;s̳c���/&�`ή�.	��ϭ��9+f ���ҭ|�Qq��s9�i�s��}�)�.��@��� ��nw��'���ʃ���$������z���ޘ�y�����܎���MK�npճ�/@�G��F9�ɉ�ށ��_ ��-]��`�����6O�d]��]t��)�?F��`u��>�J���o��=��:��y����GD�'���S�g��Ié��Slg�E��֝7s[y?hrV�w7��7_����A�퟿/s��.~bjD4�,� i~���7X�[s�rV��aq��L�I�Iށ��_ ��-]��`��� ���M\�EݒXM]�Dr9u���?%l�wV`{����`)"Ă��rG9 J����'蠜"J��YSS��tJـ.��@<��ϭ��?��;������j|�y	�<��*���p�3�U��c�v��sL���a��@g�g�QV]ݘ�o0�J��֔�>s���]g@{*	�.����&�� <�/ ��nt%l�s{�.)�Ax������ߥ��}�)�7��@=�g ��f�TČNA�H�g��[0����wy!�����P�&�C��,� ߾���f/��x��s�{v��?r=̍�q�����hIo�%�   l����vvz�v���uRmcn���f@�I��pd7]�I��fؐ  ۶n�:��lQ/T���n���mZ�Z�$v^�ݔ^�e�zC���h���K�4[��vLn�ź���c����v�m�ۓ��0uۛm�=u���������;�V��Ñ�șsA�\Y�Y:�{\�$�5���w��������v��__]�G����6y�����OL�ծ%6H*�=v\���皣:]�Ri'0�1�;�����ߥ��}�)�7��@3~*+iĆI@NN��7:%l�s{�M�)��D���ٚ�Ȳ��3*�Jـ$�� �J�s����np��3=����.������s{�M��y��:��`�)h�X��919;�wl�߭)�>ݴt�����N���]��>u����v��V�4�9�T)�{n��h0�u�Z�3;���E��vj�_�������@�V���`�+�����$�̗r�*�����y�gf��]�.1�(!)�U>���$���f�=�KW�y���~��9���8c�!�4�~� �N�>��@�V��m���r$�&9'z�����t%l�s{���:���(��K	������8�G��0��`۪��o��~�}��Op<�,�p��d��z�Q����6�G`ۃfv�\��0��l3pv�.v{雹������̝�[0���y'|���]߶����fG	$8�7���}m΁䭘���X�"QG&''z�����t���\�Y��"�xhMw���!
�%JIA+��P�)!Cv�6�ܼ�IE���*BIA`IP���TI��HlJ� ��m�cRBH̻�`���a���1i�IP�B+�����E���U��HCJj�@��4��D�D�x	� �ѷ��ЀƉ@��}O7�2qBT�K�<H��<��,��cU�*����̓�y���"ҴRJ�1�xB��H�iB�-��yO�@L�R Y��M��- @I�ht�1UM��#���q��y��P ���!T4�1�p����Ѻ6�M�G�6*/����`<@_O�"�]H��(⧍��B�V��٩'�m��)A
l�M�\we��@ϕ� �u� ��{�i� �t/��L�5vUsu�h�� ��{�i���N�������% ���Q�J۪��ˮm����K;b;J�2u�^]S��mp��<���>H���ހ{v��l������e8�/����9�I�]�y�x��0�Z0y��3!>�[N$2H"�p�e8��4��}�`�w���%EFU�b�I���7�h�|�c�>�<Ӿ��B� P&˲ȒC�� ������5!��~\mA�6��Hp}�m�@=���F|��=��N������G9�����|�Cg��;dU=F
��󂭇�1���1� ۫�b^����X�4�Mt��p��^�v��֌�i���*��C	��I�;����e8߶��@=�g ��e���x��m��l�<�=�4� �;F��D���Q7U�Uـ���o7@=v��l��߷�����~��r%$�U��y�x��0�\# ������>�;�߾�� Ul+���  6�m=-���ߚ�����ٛ]rk�M� p�������"G�ém�[r@  J��U�j��)u�׷�I�:�� d$r��ײ]�:3`3���#����gv7-�N-�<덌�l�����{zv�wngq;�;��E^��rv��G��F��C�"ѺlXl�y,�l�Lre�¼������������Z���U=���3q��ݲHt�L�ݹ��q;Z;a�m(WU�T�1b�N$2H"�t����}zt���?�Ds���4�5q.(*4��2.���4�ـ{�=�4� �V���1#߶�6��̎E$:�O0��9���}����gE��X��&G''z��8}���֌�i���9�~� �*�˻�|�{������	��W�N�泶fy��v��U͕�)2�ת��n�q�۫��1�<�.ǆ���[f��[0�Ot�;�7�ـj�F�bK�.&������g�Vc�ȏܳ���#�H>���k��@�޽:�����"N#$���l��up��r&w�h��DL�Zy��X:�������,&��T���`���w�%q.(*4��2&�k3'@\�����������*�WE�2�kCg��;dU:�h�|;��7|R�{]V�Gi�ٌܓ��.�R�l��uQV�����������;�h�7Х^%��"G���l��up��i�߮�����G����P�`䄓5$��kRO|�954k[%�5�!����0��/�B⛂bJ�.����΀�[0i=�4���#�߭��:��b#D�� r>��{�8��^򤧠{޽:�!Ի��.���n8�-�������*�t�:�e����a��������&��j���m�����5�S�wu� �� ���M\�L]���������4���'��p=V��+�tC��Q'�qt�l�9��@<ۼ]%8��r�l����$RC�}woz�p׺�&
��$*�ӪJDs0��� ����"2d�?�� �n�t���h�9��`"��'nT@���KUsem3G<�!Ƚ�I�,��e���c;l�pl=�,x�k�V��]%8wZ0i=�6� ~;/�L"1�Q��.�����{� ��8k�\�ϳC���1I�ٛ2sX�@<ۼ?���gߩ��V����.6��)0$�$�C�b�~|ߩ�¦|�рw�Ots�uSW3S�\�]`�)�<�рsI�_ �g��s7]���rH�o���   m��&�I\��r$:re���i�mm��6�8h�ݰ����  	'Gf��͖�bӪ:��u�k[d�GU������U��.�v�`v�t�g������G;t�=�T�R��F�f}tGq��e�u�p��9'�!F��>�����a��Ŏ������ϐ;n��]q��8)�NL0�30��Ԑ(��	 �S^o��V��)6�6y�	M�T��R��7F��5e�^�����K�k��S��������&�3+�?��� �Ot<�`W*��ڸڃ�o̒E$8۷���u�9\� ��F�(�S1%�qwW_U]����X�Z0�Y�/��6O&�.
�.n��9�D�Z����:��0q*u����㛂bK����6o+@歘m=��U�k��}�9�xG��q�<kC�)���B�Q��݊%�b�L�W���u�&"4LRx�!�6ݽ����
��|~�i�;K�.6��G1d�7�'k���v� �~SL�"H,�	"H� H��$��R��"! R}]��RN���ԓ�woz��P��q&�d�Ĝ|��_ ]\� M���n��N%�F�5q�57y9��5I� �Ot<�`o�����6���3$�r.����#�u�Y�9Z��o��=�ٗ/䛜� -�SD�Qs*�E:W7n���T��92�ݚ�nGiՊ�5�盬��X.�S�&��p�T�19�O�U�k��up�{�9�� ~:�n	�.*�*ͬ��I�_;Z�s��w[�E(JA�U���U���n�١�Dh��1Ņ��A�M?�:�t+�]Ȏs�+oj��?V���9������|J��@��!m�8M<�誫�Sgj��zB;`wM�U��]�`+Y���8ѹ�g�r�6�n�`N����U�.�� I����`@�+�tc�̍>s�}�s�37m��Su�9|�?�����s�Se@U@��B7 ���ށV��W�|~{��w��h�K1�9'��އ����O���U�7ջ=	눁w�A#��D$H-і4�Ƒ���#����쾐�d��I�^Ysw]J��@�V��|��&Ri� �~��t5kN��?c�1�`!T��`3��ՎZ��t��Ltdzz�Slg�E�������.�W ݻ{�*�_ �����49���5�qp۷1��n�u�9kk���g�c�(���G1c�w�U��U�_ ߞ���oz��B�nD�L�8����"9.���i)��V`8�G"#`�wm�@j�\PV���UMw��`i)��ɚ���~�S� ����?�����J�)D@ +��D ����∢?������P�!D�u��P�U`P�@d@$D�E"� a D�l�C  
�
�������
��	xn "
���D�("��*���H�����"�PDp ˠU� ����Ȋ��( Z� �ETL���rEDѿ�^y
�#Z���Ȫ��",�����l*?��5��?��\�������?�������@����s�>����������?��|��o��`�� ��O�����_�����
  QDAɀ� b��?�.���S�a��#��?���'��D ���i���z�����s����5$W�w����P��?�������8�H��j�)TQA��D�Q"� �Q D�Q"�Q# R@�ED�Q""1Q Q �"�Q"TH�D�H�H� 1Q �Q ,TH#
�DH �AH
,H�+ R(�"�H"0Q � ��R!1Q## RAD�ED�ED�H��Q �AD�H�		@��"���D�Q �TH�@�0"+ � �� �ED�� R �THQ �@��H�Q"��D��
� AD��D��AD� @�# H�@�1Q HED��H!
AD�Q H!*�Q"��@��D�
��TH �H$TH�0"D�$HD�H�
@��D����"�B*D B"�!��B( �B*�H(�*D �D"#��B
�H� � �R (� ��B � ��@��H"1��"A��B D ���H�@H�*� �"�"�(E D!$�BBP�� DY U���@H!��!"$P�DdT�H�P�1(B, �P!$$�DE$P4TP
��� 
B*$�)"�H�$��"��(��)Q�)b�@`
Q�cf&����]����" ��EO�?�$�ry���_�;U�Hl?�����=���D ��G�����C� �����6:?���s���D@ 9��F_������R� C�D ���"ab���%�  ���߾
� �p��?���Y���t�DQ�ɬ���G�����z�o��D@ %����?�������" ���?�A������G��?����JQ ?����1  �`����OCL�=?�?�~��4����?�P�q��?��D L�*��!�_�)�����D�A0��?������Ha��D ��O����,���l@ +������e?�o����?��`�������e5����<Ou� ?�s2}p%|(�B��R� P	P��P 

+A�h 4��
� �%      $(�)!QE"�%J(��@J� �BIU@
T H
�U �D��    �@ �@ K��go�r�����{� 0	{���nZr���A�w� w{m8��q5�  Zq�sne�� �꺼�ֽ�o/o8t#��瀽�^�W��6�n�(qخ�;�vԀ�UB� D��
�T.\ ��B��D@� w)JR�h�s�(b�S;�: �
� �J1   h�i@��  :X� �,` "h 3� ��@�΂�� Ҙ���J ���R J    
%�0 ΂���,����>'�ۉһ���W��ﾗ�k����=;��,qT����p #��O�y���� �n�+v��N}gog=��y�� y�;������<��_o ;� P HP �0xs�w��q����mǸu��&��χ����s�n�\@>0 Δ����wo ���ϰ�@
�&�{�����,��<pz�8 �Y�{G��/������v���   H ���: �喝���-^�@t/���\���ӷ��1����;�WyǾ  ���rrz�o����#���>��<������'�{W��ޞ�>��yz<    4���{)J�1 ����T�@ Ǫ�I��=!�FF@b'�T��J�F LES�Д�U)J�  E4S4�@ �x�����K��J?e~����X7J��Nۿ�(���.������
��p(���x(������S���$B���"#d��d�Q�a�� ����g�~���zq�H��z���Y54�o��e{}��H�sP����I$!tk����
i�fx�"�4�X46�K��	P��Wf�r�MU�7��M���kW�ߒ�%U�d��+X@�^U_�gm)�U+PBB!IX��/�Y�L��~^H��j`�u�~=�jA��`�t� � SNl���4f�8�t0
h�;!(h�6p�N���d6���� &IdYy���g�H5�Y�ī)��o�l!�?R��4F�F ���)��H��e5�B1�����эA
��j����!]��ѓ��%92�19��y��V�w҂�^��-�B���73b,�K0�B�Q��3�8G��$��+�z�"��)�CLZ.�"�c �a�bT����;=WL3g)�aCEM2!	 ���*�6h�/�׆�ǓFԅ��ݡ��R�V�:E.�.�Xu(�q`�2E���]9��!�8B��n:���MHEh衭�8�s7�6����ф&�~M�8��$�YA#E�lJ�SHq�$�2:��7h�~H��@�� �2ISX`L6i�f���'�i�Xyo\����x��/,w)`)}����l!��L^�s�։G{K���=�(~#HI"h-�$(�Det>N'?a1%tc�H�XBP!��J�B]��`�ռ�!�5��]�T���$)T�V�d�?,\�x��+����&�o=f�Ժ4R�^G��K�U.�J��=v-�]�e��ZB#�&���V�(jTя�Al PD��^�sQV����U�b^������\���M�]�ϫ�cMgWP͇]<3���y��'-���<4)���4��H���P���JF�2���`l�č48�xp�b�8�
i�6D+�����6q�g6�H�|�!Q���%�e�f���x,+�q�rM�=��ܙ���BPa&$��p�5�GP+��/���4g6-+���$�dE��s���7s?'�" �BF0 E($��+�B�)��F��exaZj�8�$H�M� A2����'�sb��U��5yD��X��$��?B!kr]������ �� 16�*�������
h0��� 4�`�@�`0JD�!)�Ѯy������%4g&~��;��aWD"��pw����՗�.^pM1�J�c�Y�0����?)$ѐ�p����̏��HSA�M�lu��ō5��~�F~�+�B���z㽸�r���Qy~�B%
�#��:[�8D�����O�&�	M/���ƘSZ0<��)0�
�MB�N�[�BBDr�Bإj����C��?�u��%�@ B�0����?&�1|kEM!H$H$ i�� ĺ���Յ5�Hջ<at쌎���5�I��o{5�I��`Uk��(R�7�!$@�Z$a0���#�	 F�		!��cQ�c4g3a7�!N2DF�%u�7�͚��%*�VEo���Q�"&R����Gg瑮�G�x�	4����I��4a�M�9�|No��@��)�����8�4�bo�E�~$dt�]�5ӂ�>�������4�1�=s?N���k�?�1"�F�!��#�8F�6sQ|�_�x�ŉ45J:�~|���U�c]$J:��הz;ڦ#���b=җ�y� -KNݰ(B���)�$BC@c-�2��B��?~�^Z�Q�8;�!�bX ��C�$Oe?������������d�)�g�?���CF;x~�I�Xl��4f���i�a����`A�$���-e/�T��	�	� Cz����xg%�y�D5Á9vT�\ڙ�I��\�XB+5YP��SE#BE`B��$� �c	��Y!��`P�X��E�F��0�+���dtЍ1�.�aZ�,��*h��%p�f�H�A��p$�l��X� �bB��%n%������qڄ���i YВ��R]�U��9�YrY?o6m��<!pȒF41�iXџ���@b06/�`���A܉�q%�ه��!H��;H�4!�:_��K�bK��5����1#p��?�2y�֧vW���)R���t���rT��So#�F>�.�H@��]<~xp�Ѩ�Cm��̳Ț� lcEp ������ȘB�.�1џ�DJ�hYb܊ܾX�P�DҚ^ν��i�K5����F����!B���N�ĘRE
ۜ�y{�������j�_t_�JR$||<w|ѡ�8���MD�B��F<!]��?xxCa	hk6l�~RbD�_�Yl�"�����CP����nxh�.��֝7A�n�0�$�M*��!!A�q��!]�b�^ʔw"u�v�!�<�ߛߏ[�0� E�Ѕ$��IRPa!i$ !@D/@���D����jZ�$)Tf��I��y�k<��3E�б0 I�@��6�v����]�)/߆4m��d`J�"�$�
@�b���B%B��C�\�Bh�%�f: ֌��+��IB���XS� �,�����a$7$�2Ah�*�t�A�]82��K!=&����lq�i�;ׇ<)�F%!R��+�htR X�%u)�]��	�D�! e������v�R����u�;@�V)x<2&)�����nD �f±�d�����ւSY7{�^s�L
]ZK"|�����xCF&����thp����
iH�W@F�
I��M?��~�tE�wixF�#CB���\��� `s����S[�6p�������^	6*@t�ٟ���Xl�˿�4����Z1���� ��!!�i���ч�����O�)�&8��N��7k��q���(�M%��W�7<ۘ�)Ĕ1.~���{���==�hMa�ל�Ca# B�i�Ǆi���h�~�~�L��~�\ șn�=l���Y�YA��Y�j),ܟn�T��*�*�tjHF�(a��/�$盄 ��A��"�`n��L�a$O8���5$k���@"�1 0�.75���Xo�t�B��� �X�q�MS!�HB�c,|U�
Ѝ��!�ច��T��)a1��MZ E+��5�D���i<D�󚹳���t0��G��SC���7Fl���8�?fl�&�2���9Jh�%���}���^N?�h��h	�I.��$�B�B~��R������jĄ�����u�MH�e��h��<0�2\d$���)�"Cэ1�n�o��SF8m<4c<3��W?s�h�hԉ�H�`CIY4ʻ��~�m쪍��V��A+�T��]J0,
j+������������                 m�                                                         ��-^�]�vh�3�ۛ`�km��m���?����    �8mk���qm$�@�a�l��l�P  -�6� 	 �{�[E� :���2��nOU<�N��ة0iT �$��J�"]0���l����7e�:W��*W��yjU�V�/4�����%���kM&�m� ���m�8H�ͪ���ٶ�mV܅0��R�G*���   m�dU�v  ��4RںM��q IJ t�8xId���,�HK(sZݹ-'��                                  [@                                m�                    ?�                 Uv�                       ��         �                                �-�                  ���π                        	                                         � -�                     �|    ��#�k���׮��FX��8��V�W��d� �����@&�]��   $H!&�UR��1H5��v�
��E�qWm�9CS�Յ��f�m   �l�`�����[��N�k�Ä�n�m�ͪ�a���� �U��н:�ۄ@�)C`hia��� m�g^�a�`  -��a�4Iԑ�� Smulŗ���G6��"^T#���mSR�c��;2�q2�ɮ�ں�U�v�I�nö����@ڶ��l 9m&�'}NT*ǲ�p�UTU6�BwU̪���UUlIg�� %ؙUZ��3ª)����� �U*�5�	-�m��\	�F �Z��m�Zl����YvRT'U!�<��<�p�J�TF5t�nj�@�X�U�U�A���^Z���U^�� ��`^�6����j�Rg��j�������z�۱-��ɶ�[@�� ^��5�-p�d�p ҨR� 9iV��l��r��-��m6�g8ڶ�� H�Ѧ7f�m��Hۺ��n�5m��T��CaV�34$���W���qmk+K7� ڶz�M�h��]��g�Ut�V�ʶ�r�WEh347���q��t��"�*���Q�����Mn��$׺*�,"��5�Jh�UUU�XI�v�]U��& ���؛Y۱ �0,״�oZ� �m�l[]��-�8*6�V�)-UJ��@uR����YM�8�/�:��M��%�ڴ��,WT��LUT�3ʮd�l  -��U�٩V�YI���M=�ܲ�:�*0���k%�~�i,����p冗��Px��kh�$.�3�����6�F��w`�TVV��Hw!�;mܳ���m� nݜ� U[V�%=����c9�v��m�3LV���C��6-�AT��r��,�5uUPm�K��]ߪWΐ:���$�&�]b�%$٢���m��8�`L��d	v�P��Tkh�p}�}��}�$��c�lֲջ �Kin��m[�� %�4����8�f���x�	^ۘ�k� -�i.����vH�T&�U`���n� �l�����nʙ`z�X<�:܂�<��%��q���T��ؐ������0��n��Hh��p v�L��ɭ�mݶ2  [iu�[�g6ط[��  �mHi�Xv�·)-��m��$8�x8H 3��ai�H�vm& �l��9:87m�lp  v�%�i
�*��"?}�@��M�P���;�  m[q��d%��6�Z�7Vmإ�R'm�@�d�  m���&À��'q����M�۲�pl����Wv�V�Bh��[A�m�%�@��#�֠U�(���v'����U�mJ������+���݇\�ڪ��U��6Fc��k���x�!� ����7=�묏�r2e��,���RY���h�i��6�ʲ��g�K'}��Rk ����">�שz܃m��}�|-*�yUU��.�3�-UU�8s���lճm�	����w@ uTlRa����� �l�� ����f檪��]�+-�=��j]���l� 3l� ����d-��h�c�� K�i4���٦�l�P[@j��$��$����I���m �z�����%�  �v�Kp�m� � m�� q���7ٖ���r�������m�n
����@�0 �UT�(���&�sz5�  -��z�m� 6�� t�/�� �*��j����[��Vݶ�5����� � h ���F��_���ߒ@��-Z�q� �5�k�5�K��R��7�J��r� ��j���v���KL������6��� q�8���zx��H *�	��la�9pK9�8�(��  $����pٕ�Wf�کr`��&'-� $26�� �T9j�b�(
��(R��]���M\��s�l�Q��@��*psQg����v��M��eݠ�7VޗN��"xN�^X�n��tWj���y�v�έvؘ�<�e^7��Ls�.�yn{x�,�Ta�
�Y݀r�pz�ȵҲ�몫��m%��<3@V�mT.	`N%ٛPp��\a�ҭ�]���ږ�Y*i��۲A`�T�v��ixR�U�UVQ;#ż:;Rj]��2�i��l$ [xhL���UlpR�+rU  �6� -��m�7t��z'j�g@���8 -� [Am ��n�e�r�`	�pzk�F��-�3���Q+�"���1T��sJ�-V�T��1�   6�n���m� �N�׶ ����ֳIt�q#��ڶ [Kn� $ �j�Ŵe��U�7Z��g06�m-�m� oUY#�8�I���a�|� Y�:/8 8�6� l�}����Gv�m� �� �-Fڃ����@$�J�[+� �2��O.�UG�C .���k/$܄Yye� R��h �`�K��m�'�u6kh޴�m�	���l�6�s��F��K�N9m�nx۲C� kd�\Û�$��m��Px�h����mX����w}������a�ۋh�  ����<WL�5i��'��9�xu$��8{lJ�v=,�m][-���0-���.� �$���acZ.�g^�6��� �$m����8Bړm�N��%t����
��4���p�J������\�`.�IBC,�m�T�Jvv9r������ȢCv�I�ױ�4$�0���cm��x�h �mGk�� 6�������}��o��CI�ؐ`8�d��� ����5��L� I�,��iV��Wf9�a�����A�`2khNnduSc�cd2�r���P�fN�f�$d�H[@`m�`  �nCm��  4��"�@���� j�m �V䤲J$�l��Ͷ �H    ����ζ�6شͲl�dhL�����E�A��U���j�΅U�ֻ#�M;@:⮭��XP��e��V����w� q�o�U�� ؓ)-V��\�T�ʕ�F�ݪ��Ԯ��^� $���x� $���u��W �m�	��
 X�K7�v���f�����[Kh���l��E�^�vͱ,�       )A��[@�[k�����j���`	6Z  �  m�gjP(
��QSj�̩5��,i�kGYa�� z�6�  �cm�   �@�4�֬�-R=���br��*թ
ڠ��A��m ����`-�  Um���    -��m�е�m�  6�i3� kR�m�ZU�U�c�ꪨ8��6�m�p�	9��H�d��D�k�H$A�n���S�AЩ����GL� �� ���S�T�|T4E����O�_�(0T��A6*&)� ���P�>���? iG`5��1��!"�B@"�`�`a B!A��"�����;"��J/�@����
,"#���B����(<CK� � R���4D@ Q14� ���R�U �
�� !�� �+�@|�>��.� ��6*~�(x(z�V �'��  ����D��WAb��+�j��"�'$� �`�X�H� ��X��B2B,a&"�B"ā�$X�$V*b#���$���(��
�E��4��H�X0�",���D��iP���ă��@!DU�T����B����@4E*�b	b��x*���Q(z�8�BAI��}6����t*z��S� ��

x!�T?
��O��t��S��iD���*��*�Ph0E�m
(�C�`&��Cb�Z�]���,ȠEhU ?"�ч� ����>���x�#U��Z��ACW���              6i�Gl���@Tp���#L�����{��3٬��ʩ�! qs`�P�d�Y���6�5k8�            	    l  z�   "tm�m�     	�m�  l    �m�      I    �	7�g���.�$p�4�lYz�ZB���.QY�j���!Z����Җl̳m���̩,su:��N�T�9_6��5�[N�$� 9��+��j��b�g��������t�XE�u��0�Ls��w$R-H�97%�w,^�#/\q�6�����!v���\F;V�.��R���+maFОݵ͜v8"�lH���;M���ĉ����F��Y`�G�,�E�!��͡�W<@l�H�nΝ�nn(u]�ڧ9���mm�B �S�������״�h� r^�Ή-u�c�vHc��Ӥ�+oT�٭g��ˇ��y7%Sw<9�n����d��h6[����r�[���V;lt�ģ�s�6�n�݂�So!l��������[-����<qϭ��\v�p- �>�7�]����.�Ws��1�:����܅�u��ו'�Ӕ���Μs#��G���ݕ�������AU�L�������v�]��nd�m���$h�a��8��U*��0�򳲇���ڽA۴iv�RU�)؛�#k
�eݢU�nt�e���6�<��S��{�mH����+���.�ny�1�@r���3�B�j�8�.�]��Scb��6K���'Hq�e���-m�p�4l[��	�z��Ѡ鉵�:�&�kB�*�
e�
�8�k�A��k��٧q�3�T�t�m�L���mj)ЋҚ6K�h���M�M@7P�5�Ԡ�ƪ�q��5ˉ@�R�F���!��˙�3N�0��*��	���T�Q|���p�;CJ`��7�fI�������ݥΚv����H �m��8ڶm�����˼�n�m�U�ݛe�G�NԼ���1�s��8�^�St8��8�z��T/FNs�8�c�zԧd�@���om����L�"ħg$I4��ݥ.m��H����#��܃���N�q�������g���tm�/Z�׃����"uj�y�������{��������~?����@8 χ�	�a򢽔ʂ��v��94��&c@�6g͸�z�h�������Y�}_'���%�L#R��:�[��f�����D,���F)�#����ހ=n�7l�u� �+S��쩊��D�z}l�>�S@�ҚWkz�u�1ɑ5�D�&����h�S@��o@/�����pJF	%�*�7j��s�/n"5$�0��f�����nn��3N��9�����I���M��� ��h[)�}��mq&�#�K��pe�]��)5UHT���T��ɳ�wvi�3ޘp?b���2�L��$o@/����i��/��Ɓ?ߛ�-�^,za0QcDRM�e4��:�[����~��h��x/�� �7!�_t����ހ_u���hޯ�����nV�x�ӗ�ϓ-�$v�/Ru��q��H77,i�$I�X�Ib0��4����;�<ݳ {��V�%SUwR��	����Y�}l��}ҚWkz�z��ȌdQ,��&����޶aJ!:J �Q
&��uX ��p3�^
�J��UIﳟ���� ���0.�U8�d�(�4�4������>�S@��M�ث��x%#q��������٪�i�u˫E=�3�BK-EmN�X�e.��8̃�S �I��@��M��4����+ŏL&�DRM�e4��:�[��@��OG�
nC@�}V���ޛJ�7ٳ�~ݚp�8^[i��K��pt�V >�x��`Db�{-Zg<1\v5��O�o@/u���h�ՠuv��ux�dIH�k�خ�&�:,c�IWn;g*i�2�ǉ,kכ������ͷWW5ѹ�B5����M�ڴ����@~���֬�r3$�dp�/��@�������Қ��p���,�EF��@�������Қ�h�㸇��d(�z{��>�)�_;V���o@��^,za0D ڒh^��/��@��o@/u���� m�GR7C����$��t�g�Āh 6�6 )D�8 ^��9��kv@޽��q���Ăݶ0�C��=..�ux/gp��Xۑ��b�=��f�n��vT�n0ف�^�؞�N�)t�K��ּ�k�O3�9���9{8�:��ݸv��22M��%q7����vg��ex�������=`�vn������w��~��UHȁ��K]�vz�sq2������]�V��ӯ�����({x��ض��x���@��o@/u���hu��K�d`4��:�[��f�����o�#���?�/�(�D�z���@��M�ڴ���޹\ȦD3"�dM94���/��@��o@/u�o,t�!�2L�A'�ڴ����Y�}l���ع�r4&�m��,nBH�<�����=�t������v��=��ˣ���]�&E��"�:�[��f�����RU���|j�L�b�ӊ9&��$��=��BB�"VՉ?"T��cPB�T���Ss�s�[�/�W��L�RM�e4�j�:�[��f��|�
�#�����mS�M��3ov��d�>�S@���F�0���ZWkz{��>�S@�v���K`��T�"�i��q]ˋ�{s���v9ڋ�<�F���nn�<�y��zp�;�<ݳ {M�Λ��֫�ȆdQ,��&������e�]�?{'5UURl7V5z+�2�PPn��7ټ\�y�|"��k�R�B�٠}zS@�;���� �,�9Λ���� �v��<X���q���Ab�7��f�����Jh]��y�� 5LiBs���qpu�P�vdm�=��p��p���a�<8�,p�`� ڒh[)�_t���˽�Iu��͜��]��Դ�F�4��:�[��@��M�#�F�0S#���� {��7l��� մ�<��LYr�Tw.����f��vi�3��B���T� �iի�W%
��U�����h�)�Z�@/��������� 9���卢$D�8���I��� 9@�'����.Nm�F�d2	8h�)�Z�@/���e4{9\1�̋��4�4]���Y�}l��}Қ���&8̍�A"I�_u���h�)�Z�@�r�X�ȁA�$�����I���}���3/2_j�$��6p~u<��x`�F�4��� {��7l�:$��j����V�ZV\]p<�s�ܐ����Z��   h�m;��ʨD5�X�:v	�u�|u�Hk;��q���:s��c;��%�����Q�r�r󗈦G��d�Yw%�mƚ��d{���Ƀv���|`Gm�����{  ����m5;�d�rW�Ⳳe��V�۝��F���p\��p�Z2<�KJ� -��w{������U8+)q�7u�=u�v���/�>�<|���Y32�	����G���$�����G�y����x�[HSʝ��,"��/���9�IR��۳N����-vǠz�s"�̊%�4��<ݳ {� 纝��w�k�V
䌩�p6��{�ޮ�2�`�w�n�f��ZV%r���]M]��u;��� �v��<X�������B9㫰�`�w\I�u�������:N��V0�Ωm.�sp��7�f��� �u�0��|�G�?+_�~���ŏL��RM޳z�$�T�z<��3���~���[l�JMI%�NOG��E���}�I^�Q�$�����/JMI%������Q�ѯ�%2 $��J��ϾI"��Ԓ^�~ϾI+��5$���]�ƿ�QƤr}�I�&�����}�I^�Q�$����䒽1FX�n5���W���tW����v�l�C�ڻ5�A\���zn��;��m| �����}�I^�Q�$�����/JMI$��厘���!����䒽.�RIWy��[l�L'm��gW{�J�+�o��7��`5F��Ԓ_���O�I"���?�Ŏ�o	Z80I�U"��j�huL����c�A],BD���ZtP�i�%�e�U�P�$怗BAf�$"Q�F7L�h��J,�� Lby�d�͙��4��3̱Ic��I!�OL�~�h)HD�*���N$��k�
U�"����K�$d�����H�a�MjSF0AZE�	 F$���
r'�Q�!���F5!H$,$ʧ��P�+�!@sP��X3s��#u�4����q���ˬ�K�CB�*��x�3jA�$��sW-��`M��Bfj2,�8H�bh�]@�	u ���*~����`����ʀ '�!DS������#������^f��r�}�wvn�ot�!�dh�2	G�|���뿉�6���]�m�q�m�W{7/gz�{z��3VLX� ڐ��K޷������?~��$�����$��)5$���W���U8+)ӳ�ݹg]��S��KI��S�]�t�p�n�:[����nŴ����6�{��������޶��L'ԩ/�_�m���Wz�y�����qF\�q��w��}����g�jI.�}�|�^}u������1\�_�(�cR9>�$���5$��o����o���Ԓ_�����9�W2)��dQ,��	�/�������%�;�7m��{��rۏ�ϸ.'`�������零�}�����a�%�E޶��L�8�o+�䂕sw���l͟RI}ݹ��\�ch�ґģID�Kp���c�;=��л�pݮ��d ���uuQ_���_���h-ơ.F~m����ӽm������~���UUK�_�	,�6����p �o����&��h��� ���~�ϫ�II������~���������$�E*JH��_[-�dP�r���>���m���p8��*�RO�v���m���RI|�wǑ�ә��/ؕ|�3~��8�o�ݿ�z�g�L']�߿{>�$��=�S	�n@ԒU�ד�m��%�J�{�?6�������{>�O���^�w�ӽ����m�cf�]�$��l�R�[X l ��   �@�&�J��Nj��z��c�S�6p�ay��Il�ʹ����8��ڰW�.R��7�:ϭ6�^#�w4v��M�[��|` �C��u\I���\�6�o`�h�vx$9g<���8渟O8��;Z���B.�%�Bd�p܋h�Zl��d���{��=��w�>{��J�����_s���>έ�d�k�B���,�r�l�{������y��tS_���o� ?~���[o�����v��̽��m�x��5p�jrܺ�ɛ�������?�S�����m�{���[l���Wv��r��rDI��(�}�Iu���J�z�w�R����M'm�۽]�m�����dXE��DjK�fc�����;&����~���[z�+�sz�6�����E��]m_����o�| {��������/y��g�gm��ד�m��O-�=��U^Z����Ԏ'c*1���ZY�,�n�^�3�������N����yzě�ې�m��n�w����8�6����&��I~�m��4�m��MObwv�h�n9�kr�y����OD !Q =�"*`�k��z�u�s��=�}3v�~����� ��H�U9ǿ����q��m��߯�s��?y��ݽQ����߸s���s���˷�?�y��t3_����xS�@� ;����f���p�-����g{T�+����޶ٗ�ۊ�DV,�n]]d��m����-��T�D�����I%�w����H�JMI%ޘ��	H���V5/cmu�^�hɸ�)'S�����v�Y��q�;�ݛ������99;��Iu���J�Wg�$���3��]��]�m�W�_�W}H�[�BI������������N6��f�w����8�~���W�i��b�1L�#r}�Is�7m���{Ü�"{FE�Q
@!���J�F�B:��&� �I�s<ݛ���^�]�r��^,V�|j4�[!v�'U%K��$"������]�m�����m���y;���_�&����m��>�.!ݲZ ����[o��q�m����R����=��3g���K�����<��F������%�nV�Gzrݹ�k����F�Ժ��9 �ڳr�qk��@]f���5Ym�a3Y�g�m�kߵ�s��?y��ݶ��y��|P�"ET��̶���vn�o�p�鯮WR��.�Y����g�7� ��$XҪ�s���uw���O�3����e�����ȱ �D���g�����W�P˖���Lݶ����r�y�����'�$F �B9����_g9m����7m����k�k3,u�!�5�9�oQ> 1L����m������[l���o�J�R��)UU�n���m�Z�B��D �(K��m������m�����+�����K��o����K�Ԓ^w<J�bJE�W��۲���m<��ʲ���2�"M�9��W��0ֲ�D����f�.e�h�ᐑ�;�H�����K�v�|�^�u�����zD�;����%_�?����PD ې�m����;ߕ*�Il���m�^}N���ޘNW�%K���{�������hp�w���O�3�����w�����T��s�7��N6������[o��d�ȭ�ۈ��$gU$��3/gz�g�i8�o��a޶���J��7���gm��j�_�n�r�(�\��m��0�m��IW��|{�%O��RIy�;>�$�fQ� I$�*��.�����\�Չ@8 ��8�ms�p ^���y-HY٦��sm���1��[#�pkN�p=GN���vn��c�;�i���n��9��m�mմk��4`q�U��X�Z��89{i����eN�IRq}��^���m��۱b�v��MvK:�/:����w&��Ӝ�����ۈ ͭ9s35���k5�ʈ�*?�o��5 )��6+���ֺ�9��K��v�ś���خ�Y�n��̚Ѭ��H�Ѯp��jdC2(�M8O$���'����$���6�o�y�ϕ>(�#<�-����5$���~X��9	���N|�^�u��$�JH�^��;��3g��m�繇{�%K�$o�����������y{���[l���%I/���o>;��͟�F����K�1H�PB�F����2�|���~S����ߟz�~��3���I}%�ߟ�}�IW���4=k�6�ɩ6����m�J��߿3�m����w��~�����������*d@����kvz�R�7#�=u��q��u�Œ��z�أ��w��_��lyE�D�!ܒ_�O��Pyw;4�����U|�X{�ߟ �џZ��n\�L�f]�?_<׹�Pڱ�$�Z_*���Iw�3︸�ώ���5UU|*J���'���n�;�"����=�}��;��p��E����/~|��8W��˖⌱G�������UUW﷿2���??z�p>�K�IUUW���ˀ�kW�B%p�����~�~��5UU%�̽���x�r���w<��r����p����9�{stv��I��pb틩3F\��RkS:�ᗄ5�L0p�G"�~���@���hW�~UI|�)%��2���=���K�2L�k3rN~�ݛ�>T?�����}�x������^Nm$��T*����l����p�B��.�~|���>RIP��T��D�^�_f�{��7�������R�4�l�i/��U^g7��1��Ӏw�giW�RWﹿ>��>��c�ܰ��$|���' ���U^Ͼ���~|���>�����v�eS���x+==����\�ۄ����=���0����wv��'?����|~�?��Zs�h]�����˖⌱G�Àw/���R��Uٻ|�=��pٓmRl?jƯEr+�e�|2�_ �����iRo۳�{󿖀vr�cw0��A��Ҥ��2�pn�8r����.W)$���@m� �o�����=�{��E%��ۊ�rpٓ�U%�e������<���/Wc�$�G">�|�8��(Z��f4`{]=y��V��F���� \ٳVk��2ܚ�%�0�����z� �����U*���U*�RHT~�Ͼ�2����ݲY2��Y�rO<׾�����Ab��FE֧���ٹ'�}�M�9�����(�E�E �@A�UH�%vn�3�\����rG�*������e4���j�;{�׶�W5�0��k3r| �����T�T�I$*Uy�����g� ��1�O�W�$ �5�w��7$���}r�Q���r�p���*J��
�P������k�����dÀ$�~��v����$x�m�$�$°�o|oK.�5&���aYM��.�SV�4f�Vi��Mkr�`�D",a��CB3n�oib�w9�R��g�~4�`˩]08kbȒ�$X$�E�!BH$�SDn��Yi&��;XR\B][�4����^��
�����?�T����i�h�[a���@�#??{�*I����CE�V�6J��S�H@��Y.�.��0�d��m�            ��� +j�,�ب�WYb	yo8�vPy��=�&n�7[A�\_?1��Ig�R&�UEV��v�Gj�;v���(            @       %�    rIl       &�        ���       d[@    ���g���fNU`�Mcg�r�m����|�u+4����U�K�BLP-i˶���h��[�ӷet�6�Lp&봉/�K�.��ǰ� XN��3�Y[;Z�U2�dx6�rը�Ūd3Ν�������
m���}�����\i��)Rx̼�g۸��زv���ƍ��A�1<�L܃o`ÇD�t��^���eH�#�_/������y$�6K!�5�ʶ�uب^��K�%#$��kA��V�s�݂�Q��gQ�<)���[ԉ�Y��q �[�t�M �8�2�0�=��"��� {���ѣ-�9y\�y�om\;���s�dz:ڜ�
���sƭ�>v�5��e�qe��in���7TӤ��F%Zڞ;w!�R�@�� ���!�T'K˔�
��[N1��[���XS<S����N�jX�����T)�]��ZݔWJ9��J�n�j���vz�.s����yU���9���}��vক|��.܆�D2�6��>����|m�c4�pm�-U�3j���W�U��h{���� �y2]����m���ѱ��{b����	�Y6<�@[����9���'�f�ݚ�D�v]�͸�X�F�6�K�v޹���O�>~-����G5Y'=`Ƥ�f��N^!�sPu2��iӤv��v�y��w%W�h��pn0����qm� ��&�����[��6������B�ܭ[(�[R�Q�J�R�.�4�7mѫ�����{����" ��T� EP�b /�> �h���PC�M�(	���y&ffffkZ�e:5eͳ�c�������Pp� H: �  ��nB��ԫ@prc�q��ӍduK������m]۠�c�|�nw,�<b�`7#`x�P^.�,�V�)�W \�m������&�'I\���y#R�\��97<.)�8�
��n���&X��q��A|O@��9��+��k��@����%��f���%���޻���0����d5&�J����ٰms�-�X���5va����?�%͛��fLd�e���7o���??z�pٓ���X~ܚhʿa���& �rC@��vo�T�UIU!��������8���ˣ�d�ő%2�ɠz�M�Ҝ6��o3f��2�p��,Q�[N7drI|$�U���� ��|p�޼��T���8�ye�԰�7$� ��a�6���2�tۻ8s�4�Y��JF�m�JA�1<wCӹ���4��<��yӱ)���&�����豾{c$�	�nC�9Z�M ��h^�gyı,O}��6��bX�'��zk��W5�0��k3iȖ%�b_;��Ӑ��!0V�K����� 8�D��B!��)�%SX� mC�M,B9H`EX��(;�!|���!��GQ9�����6��bX�'��o��Kı<׾빴�@>�MD�<;�'��\2�S.[�Y�ͧ"X�%�����iȖ%�b{�wٴ�K���涜�bX�%��m9ı,Kޞ�]��&��e�Y6��bX ؞���m9ı,O;��kiȖ%�b_;��ӑ,K>���}�y��r%�bX��o�5��a$�C&�2m9ı,O;��kiȖ%�b_;��ӑ,K��}�fӑ,K����iȖ%���;�����Sލ$#�n�=��u���:z��	�(���X�s:����������s�&�sP�[p̷Z��m<�bX�%����m9ı,N���m9ı,O}��6�(�C���2%�bw�K�.��I��Ko���q�[!�ֳ6��bX�'{��6����QD�K��M�"X�%����٭�"X�%�|�{�ND�,K�s�MwWZ-K�q�Hr�JL��L���Ӕ�%�bX�w;��ӑ,j"4C�h�6�B ��A*$T�$T���XdMľ�����Kı>����.��I��K3Fm��m��wy��K��D��"�U��A�ȝ����kiȖ%�b^�fӑ,K��s�ݧ"X�B�V�N��7�N��7�ur�ەn�� T���̔���(�Q >�}��?�X�%������r%�bX��;�kiȖ<oq��������*+J��i�|k�C��Ou&�`.6��{�X��zw'=KV�S5����k3iȖ%�bw��nӑ,K�����ND�,K��{�l���~���%�}��iȖ%�b_�;M}fL��5��ND�,K�{�m9�Ď�j%��sﵭ�"X�%�}��iȖ%�bw��nӑS�"#U5�������L$�2d�k6��bX�'�Ͼֶ��bX�%��m9��a�����߮ӑ,K��~��ND�,K�{ғF��S-�f]kY��ӑ,K>����"g���iȖ%�bg��iȖ%�b{�{ͧ"X��	!xU\�O�"�}���Z�r%��{������ԜAd֕��ߛ�D�,N�=��r%�bX"A�R ?}���m<�bX�'�����m9ı,K�{��r%�bX��K�ܚ ��N
���v��gv�5bf]�<�v���dh�fD2*i�8 �{�"X�%���ݧ"X�%��s�ֶ��bX�%��lG�
B~���%���߮ӑ,K��~�}���KnjL&k3.ӑ,K����[N@����j%�}��iȖ%�b}�w��Kı=�;۴�A�":���'N��_kT��˫�r�5��"X�%�}��iȖ%�bw��nӑ,K����nӑ,K����[ND��7���ۿ{�- �G3_{�7��,lN�=��r%�bX�����r%�bX��;�kiȖ%��|�{�ND�,K����a�Ɂ�2�f��iȖ%�b{�{�m9ı,E���[ND�,K���6��bX�'{���9ı,O�y��2L����kZ��qu`�\ 8G����5Q�h�`  	  ���Y�^�	U�>zr�5���¢	mgX+��!��$�l���y{&�ӻ����v����n3r�#g�ۃ=�W}e7�2c/Mm��O6����&�Hh:�Sq�=�Z�0xщ��<��N��z���C�t7m�M��s��]��,<T�H�uT�ks��w������)�B�[�ޘڃ�ڶz\��n�NSS�#����]]TDR�v�w"� �K�K�&Re&R��ﵭ�"X�%�|�{�ND�,K��{v�%�bX����[ND�,K�wSE�퉨ܲGwr]�JL��N%��m9Kı;���iȖ%�b{�{�m9ı,N���K��K��Z�$��n�K����Re+��s�ݧ"X�%���u��K����j'�Ͼֶ��bX�%�ﾜ�ғ)2�)~ٖ^ۻ�K�˙v��bXb{�{�m9ı,N���Kı/��siȖ%��+vf�R�I��I��4f�챦ܰ�fff���bX�'}��Z�r%�bX������Kı;���iȖ%�e,�ݾR�I��I��{x�'v���s$�ε/���? ��ϳ��g�[sšyMa,��L��ww��?9��Ѝ�e���oq�X�%��ͧ"X�%��罻ND�,K�{��j��bX�'}��Z�r#)2�)~V���av)w-�r��.�X�%��罻NC����G�U�"j%��s����Kı;�w��ӑ,Kľ��ͧ"*ED�K���k�k2`h̦Y�e�r%�bX���}��"X�%��s�ֶ��c�uQ/~���r%�bX�}���9ı,K���k��Y4d�s3[ND�,����w}�m9ı,K߾�6��bX�'{���9İR��]�u��S)2�)~���j�bj7,��r]�bX�%�}�{�ND�,KN�=��r%�bX���bX�'}��Z�.��I��K��{h�-�w.����6�.�;54�!���(���+�A�2ssVZ9挏]p���&��}����{��7���}�ND�,K�w��ӑ,K����[yı,K�{��r%�b2��e�d� �l��ғ)2��w��Ӑ�F"�j%��sﵭ�"X�%�{��fӑ,K��}�f�ғ)2�)fh͵}���a%�|��,K����[ND�,K���6��c� p��B!l@v(�bw��fӑ,K���u��Kı==��W���F]]c�Y�m9ĳ���k߾�6��bX�'�wM�"X�%���u��Kĥ-ɻw�])2�)2��k�n��b�����k3iȖ%�bw��iȖ%�`
{�{�m9ı,N���Kı/��siȖ%�b|����ߍY)��㊱�{�ڲ��F׆B�Z��fI��]��F�S_���3����w=Ge�Y6��X�%��wﵴ�Kı;�w��ӑ,Kľw�͇�?D�K������Kı/N߈k_2adѓ%ֳ[ND�,K��{�m9����b_>���r%�bX�}��6��bX�'����ӑ>�j&�X�}�ɫe���d%ےRe&Rq/�}�m9ı,N���m9ı,Ou�{��"X�%��s�ֶ��bX�����Q;�MG.�	wrr�JL�ą����ͧ"X�%�����r%�bX��;�kiȖ%���a$V��j	�S`�&���ٴ�K�2���[�-8���!�])2���^��m9ı,N���Kı/�����Kı;�wٴ�K�q����������PHrY[]����gɪSi��\6fu����e�J�ꏻ�䱴��ܰ�$�|�ғ)2�)nM۾R�Kı/��siȖ%�bw��`�bX�'����ӑ,K���M^�uu�]f���Kı/��si�|(	D�K﻿�ӑ,K�����r%�bX��;�kiȟ�;��s������W�h���k�w�Kı>���m9ı,Ou�{��"X�%��s�ֶ��bX�%��m9ı,Kޞ�]��&��e�Y6��bX-���u��Kı;�w��ӑ,Kľw�ͧ"X���O��ߍ�"X�%�zv�CZ��&��.�5��Kı;�w��ӑ,Kľw�ͧ"X�%����ND�,K�{��iȖ%�bq�D��iww�owu�z������H  Xƭ.tӦ�:^�a���8 �`wM�l� ��d�l�&����]�͑4��Bv���ۂ�{'j�{CFp훹�}Vz#N�����<4�ݔ�]���խ���b7g� ���]١����:6
��:{/]����d�pv�xάA�Î��]�7f�m���s˵�<u�eۗ���M�D�<�t�����/�/+��\c�����e��:�ղ�Le����9��Wl�2�=�����?�6�u
��{���oq���_����ND�,K���6��bX�'����ӑ,K����[ND�,K�o��1��tJkJ�����7���'{�xm9�	�"dK�}����"X�%���k[ND�,K���6�����?��2%���}��/�њ$�-�fk�"X�%������ӑ,K����[ND�,K���6��bX�'{�xm9ı,O}쳷G5�[sRa333[ND�,�P":��w���ӑ,Kľ��ٴ�Kı;�{�iȖ%��Q;���m9ı,N�æ�ڄ�F]]c�Y�m9ı,K�{��r%�bX����Kı=׽�bX�'}��Z�r%�bX������@S�lWaoE�qՈ��9.���Kj�p�(Wb���x����wn{�;�"7wR�[����_�L��L���ώR�%�b{�{�m9ı,N���	�&�X�%��ͧ"X�%�~��5�5�04fS,�ɴ�Kı=�;۴�:ĈE0(w�b���iek�@��<|D�U�n&D�?s?y�m9ı,K߾�6��bX�'{��6����uQ,Kӷ��̘Y4dɭf]�"X�%��sﵭ�"X�%�|�{�ND��j&�}�w��r%�bX��}��r%�b2���M[/�0��$ww%�)t��L?�*&�k߾�6��bX�'�wM�"X�%���ݧ"X�%��f��)t��L��^ɚ�2剨ܰ�kZ��r%�bX����r%�bX��(��w��i�%�bX�w>�Z�r%�bX������Kı=�=�sYwD`�8{�-z=��v����]v[�8#-n�=	w6\�\PS�zv�`�U��Ȗ%�b{�w�iȖ%�bw��u��"X�%�|�{�@�@��蚉bX�}��6��bX�'{��룚�%�d�3Y��ND�,K��{�m9�H	���b_~���r%�bX�}��6��bX�'��{v��bX�'��zj޳uu�]f���Kı/��siȖ%�bw��iȖ0HD��(LW�!D���Q��)a!��ɇBb�	Ib��U�hK@ؔ�*Hξ(�#7�ؒ/<ү�p]@�)ZB.�*<`��R(5`,�h<"���T��<;8h=H,F@�D�T�� n xHR2%�␄!�Ú�BA]�a\D6A���W�+�� E��*:`�P<�# �H�*�9�I�P�P���sH��k���ć��Aڂ~���=H�� ���
���UOW�'�!���)�U(�@T;�Q9�3Ϯӑ,K�fM�Re&Re/�ז��#wj]�k5���K���}����r%�bX��w��Kı;�w��ӑ,K�H����ͧ"X�%�~��5�5�04fS,ֲ�9ı,O}�{v��bX�'}��Z�r%�bX��{��r%�bX��{۴�Kı<���{��0����3�]�y�j���-�[�=g��pb��z���}��ۻ���/���.MkYv��X�%��sﵭ�"X�%�w�ͧ"X�%��罻�'�"dK������9ı,O����?�6�u
������{��7��?��m9ı,N�=��r%�bX�����9ı,N������j#){f��2剨ܰ���9K�&Re'�g~�ND�,K�s�ݧ"X�%��s�ֶ��bX�%���6��bYI��l�-�KR�n6\���Re'���w���iȖ%�b}���kiȖ%�b_��siȖ%������ZJ[-amW��Q5DuM+����!$�c kХ�ȪHc�m���p���>���ND�,K�;,���YnY2L�f]�"X�%��s�ֶ��bX�!�@5��}�O�,K�����iȖ%�b{�{۴�Kı<�����D��N
��sq�=ˮF�W �˞�jc�L3"V�O������;�k�B7��5��"X�%�w�ͧ"X�%��罻ND�,K�s�ݧ"X�%��7n�K�&Re&R��{�ڃ���fm9ı,N�=��r�Q5��s�]�"X�%��sﵭ�"X�%�w�ͧ"X�%�{��k��d�љL�Z˴�Kı=�=��r%�bX��;�kiȖ $@�MD�}�ٴ�Kı>�;��r%�bX��רW{A-8�wq�JL��L��7��ӑ,KĿ���ӑ,K��}�fӑ,K~ ��w����Kı<��h��,�njf]kY��ӑ,Kľw�ͧ"X�%����ͧ"X�%���ݧ"X�%��s�ֶ��bX�&/�>
� � ��k� m�F��&u��.�6坭� pm pN� �@ /ZX˓S�݀��6��:���)��t��]�^�\R��%�;�r���R���S��w64��;wk��ӑ �u���������t��iJ��nkn��O���l-��g�����D21����d�-�M������[��\��Nl����$���wj�=����{��{�||�9{ul��D8}�=��X�!kے+d���]��Q1�6���ww����?9��㠵&Lֵ���Kı?�����Kı=�=��r%�bX��;�ka�"�MD�,K��}�ND�,Kϳ����4f�&Kr��˴�Kı=�=��r�Q5�����ӑ,Kľ}�ٴ�Kı=�=��r(}�MD�;ߥ�]֫-�&I��˴�Kı<�}����Kı/�����Kı=�=��r%�bX�����9ı,N�æ�Y�uu�\�kiȖ%��5^}�ٴ�Kı=�;��r%�bX�����9ı,O��ֶ��e&Re/+^[w��ݨ9n"���]ı,O<�{v��bX��C������%�by����ӑ,KĿ�ݜ�ғ)2�)nb|v��v;��㍾g,��nJ��l�ì0W[d1Qn�OK�������%�svh�������o��{��"X�%������ӑ,KĿ����yı,O<�{v��bX���c�+�@�e�ܾR�I��E������Ӑ��^B�V,HE � DRAi�!J��"%@ЭU��"Q ��5��A��&�X��w���Kı=�;۴�Kı=׾�[NE�U5��߾)��p�[���Z�siȖ%�b_>���r%�bX�y���9ı,Ou��ӑ,K������ғ)2�)~ɚ�2剨ܰ�-�fӑ,K �Q�O}�؛�H'����� �'<�ۉ�$��K�����Re&Re/�6���԰D&��9ı,N��[ND�,K����￯�O"X�%����ͧ"X�#){�5�JL��L��S�F��r]�S����V���;2�IVݎ��/���t/�s�aRT$S�it��F��S���7���%��{����Kı/{�siȖ%�by�{۴�Kı;���m9ı,N�æ�Y�uu�L�fӑ,KĽ�ͧ"X�%���nӑ,K���u��Kı=���N@,K�����k���h�sW	�36��bX�'�g��ND�,K���ӑ,v� �D8)��dL�=�kiȖ%�b^���ӑ,Kľv{N��\rMe0�̻ND�,���u��Kı=�=�kiȖ%�b^���ӑ,K�����iȖ%�b^��!�t�����Z�kiȖ%�b{�{��ӑ,K�/{�siȖ%�by�{۴�Kı;���m9ı,L���e�F���:!��[�盙zy��]�J	:Â���uMK�q���i�
ָ��X�%�{��6��bX�'�{�ͧ"X�%��w��b�"X�%��6_)t��L��_�f����h�0�[�ͧ"X�%���iȖ%�bw]���r%�bX����5��Kı/{�siȂ��j��X�}�ԗ�5!2[�˙6��bX�'���kiȖ%�b{�{��ӑ,KĽ�ͧ"X�%���iȖ%�bw��v��e�d�333[ND�, �����w߳[ND�,K��~ͧ"X�%���iȖ%�����0�`��������r%�bX�a񯬓2��.fkiȖ%�b^���ӑ,K����y��~�bX�'�g~�ND�,K�3�涜�bX�'�p���+J��Y짋���;�Z ��]Hc	��Ҝ�Wniӯ6͹+WL����Kı<���m9ı,N�=��r%�bX����5�>��j%�b_��ٴ�Kı/�N��5���I��3&ӑ,K��s�ݧ"X�%���s[ND�,K���6��bX�'�{�ͧ �j��X����k�C4f�K�e�r%�bX��>�5��Kı/{�siȖ%�b{���r%�bX��{۴�Kı?w�:�N-�53-ֳ3[ND�,��������ND�,K�w�kiȖ%�bw��nӑ,K�������"X�%�������[MF�#w')t��L��^�朣�,K��s�ݧ"X�%���s[ND�,K���6��bX�'�g�ɪ��Z��e�v�yG�nmdݥ���Z��   h�l��rV�*޼��(���q��(&sێ,[o[[��	��u�w!��X�j��ș$�v�g�r�ۋm��X��K��=��d �+ˬ�{>���������k�ֻ+>�]Sm�<n��ѵ�4�ՔѢr�5��I:�_nw7Z���\]�����d�*N�y�N�d��:�{S�)eS���x����{-��n�5'k�k'8��Gfy��Q�2 ��Y�۵�6�q?D�,Kﳿ]�"X�%���s[ND�,K���6��bX�'�����ғ)2�)n��v�l�p�iȖ%�by�{��ӑ,KĽ�ͧ"X�%���iȖ%�bw��nӐKı==æ�d��.��u���"X�%�{�{�ND�,K�=�fӑ,K��s�ݧ"X�%�/��Re&Re/+^[w�]�K�#.fm9ılO<�}�ND�,K��{v��bX�'�g��m9İ?�D�����ٴ�Kı/~���k2k��3-̛ND�,K��{v��bX�#��s[ND�,K���6��JL��^�sNR�I��I����f� )�B�[�ިⓓj��Gs��58�n.tv����^��-�\�XX���ı,O|�{��r%�bX������Kı<���m9ı,N�=��r%�bX����Zk��-�L�u���ӑ,KĽ�ͧ!�� �=@ۨ��bw9��iȖ%�bw��nӑ,K�������"|�j��X�w;�3T�[��&[�ͧ"X�%����iȖ%�bw��nӑ,~ ��j'}����r%�bX���m9�e&R���=-KA���9K�&QbX��{۴�Kı=�=�kiȖ%�b^���ӑ,K���wٴ�K)2�)n��v��A"䏔�RbX�'�g��m9ı,K����r%�bX�y��6��bX�'{���9�q���~���~�����,��;�O\Vn|�9��y�iش/)�#ł��k�=;��ci�r��˭�"X�%�{�{�ND�,K�=�fӑ,K��s�ݧ"X�%��^�ۭ�"X�%��ú�s������Re&Re/{9�)tKı;���iȖ%�b~׾��iȖ%�b^���ӑ,Kľ�{N�ə��3-̛ND�,K���ӑ,K���}��ӑ,x �ډ��br%���m9ı,N���6�)2�)2�ջbޠ��Rݗw/�r%�bX��ｺ�r%�bX������Kı<���m9ı,N��bX�'�=)֚�&[3S2��2�iȖ%�b^��ͧ"X�%���iȖ%�bw]�u��Kı?k���)t��L��_���S�ܗr���^&��Y��ff�f��:1	�S,��Iy���F��5'��5���{��7���|�}�ND�,K���ӑ,K���{ۭ�"X�%�{�{�ND�,K�f��zZ��q��r�JL��LN��[ND�,K���n���bX�%�}�m9ı,O|�}�N@,K��tf�gl�8�I%�JL��V'�{��m9ı,K����r%�bX���{v��bX�'u�{��"X�%���:k�I�e����˭�"X�|@5_}߳iȖ%�by�w��Kı;���m9İ?'��=`;�33���r%�bX�<;�w2R�)���e�ͧ"X�%�����iȖ%�a�>ϻ����X�%����[ND�,K���6��bX�'���?��ScY�/��\h�א�R� �fH瞹n�P#s/6N��V���u&�.ӑ,K���u��Kı/}��m9ı,K����r%�bX�d�|�ғ)2�)=[�!]���.�kZ�m9ı,K�{{�NC�"�j&�X���m9ı,O{�}v��bX�'u�{��"X�%�������̶f�e����r%�bX������Kı<�;۴�K�,N��[ND�,K����ӑ,K���{�X\�Je��2e���r%�bX�{���r%�bX��}�bX�%ｽͧ"X�%�{�{�ND�,K�3��޻R�!.>R�I��I���7[ND�,K�P������~�bX�%����ND�,K�s��ND�,K���Ä)+("�0���*A��(c���X "�B�b:��B��l��
�Sp� �,�i4uJN�ץ�OO~����߯�               �R��p3��+V���tBA�6�.���.q٧Laz!�Z��ജV ,�5Uj�F9y�+ 1            �       .�    [%�`       	6�  ��    �f�       d[@    Wd��8���;B��)j�v��9�b͒���:m�h2�:b�*��N�0�Ƿ]�d)�x:�&ӱ�m@O�[fH�dcH�N���ʩ��<pYĆ�x�=��q3�m��v9vv�rX��]O�m:��ӖL�usa���+�$�u[&M���]���m ۩AnCKݽ`G����b�m��$g�uc�=��@�u3E�]���s�8��g�������t��m��\��iG5$�+r��)�-@ncZ;s�LnV%�����9�.խ�.��u�;���1�]�d���vSA][����2+=Sc��f]�uʙ�b���c�f� ����c�@�W6��v5�c2����ݣa� n�K,�lb��u�q�M�ѝ�\���܎G�wf��T��+�>4�ˍ����̓�&���R@)�v�eya�֞<�ֳrv �=��4r�8�ִl���<����g���bb]�ЫdN'��ͮ����ֻ�Y[=i.�v�S�4WlU]� 6 9�ѻb�j��UK+�P˖��x��'7a��i���^%g<s�ݳY�c��3ˆ��@[�q�E��"�u6쵣G;��6.�;n�\�Fp�hfm��ʼ�F���8�D<Z�5�{9d���Jys��$�zk.VD�9�2Ӣ�V��v��cw`�i���ѹ�2,��]@�V0n����wf���hE�嵺��-M�m�M �6ٵҹƕȵS�]@Z5*���U/.�$�S2kY�.[u��Et�uJ>�L= A=P������E�(�lS _@=~�Аm�cj�.�n�z�x�[v�� 5�l @ �7:m�$�%�v�og-�u����jjśqô��q�u��m��Rn��p1��.�)�J�&��b۱\X��؅wCiT��d�pk��a9�VǍ��6=*5���L�dr�\�ϣ�gz9.�Q�lvu�:��i�˷=z#P�Lӊ�r9�f�d�,Gc�w����^����K]���ͺsknm�)N�桸솛�����8q�4�m]��T�?D�,K�����r%�bX������Kı<�;۱�Kı;����.��I��Kط��푶�7-�I.fӑ,KĽ�ͧ"X�%���ݧ"X�%��w��iȖ%�b^����r'ê��bzh��Z�2R�S.�.fm9ı,O{�}v��bX�'u�{��"X�%�{�osiȖ%�JOw6r�JL��L��bƶY!,PS$�e�r%�gQ>ϻ����bX�%��_�iȖ%�b^���ӑ,K����nӑ,KĽ;�C3	2��̥��m9ı,K�{{�ND�,K���6��bX�'��{v��bX�'u�{��"X�%��/tj��n��.1�Yc��t���j��.Zݞ��<v�r=M�t����A�Q���ND�,K���6��bX�'��{v��bX�'u�{��"X�%�{�ғ)2�)~ɚ�2Ki�ܰ��Y�ND�,K�s��NCH#`@H��`Y ��(�ԐOUh-�x���D�K���5��Kı/���6��bX�%�}�m9ı,O<ΗE��.I�ɓ5�iȖ%�bw]���r%�bX����6��bX�%�}�m9ı,O=���9ı,N����V�Q�1�fffkiȖ%�b^����r%�bX������Kı<�;۴�Kı;����.��I��Kط��nڍ�q�nK���Kı/{�siȖ%�by�w�iȖ%�bw��nӑ,KĽ�^�R�I��I��؟4�7%�⶛�an��da���u\��V�� ��	��)#sŞ��sa/R����w�{��Y�=�;۴�Kı=�{۴�K�}���������g��̀�Ƀ��<�_>T�M�f�� �͜�Ɇ�v^w�`Dby"Ĝz�U�y�����!��������$�!\%^�ϝ���T�V ����Rh~�į��h��� ��h��+/�@�w�8�ő(Ȳ	ɠwYM ��huVh^�@�ww��o��������C�Ҝ�=��9nk�=c���rm�e��7O%�b�b2�\<�v0�C"������wUf�u�?�� ���h���KY���(�$�@;��Ϫ�&�76p͚p����=�f7���%�%��I���4�)��/��h���{{+vAb�dL�$���<�� �n� {��p?*J��
)FB�]_;��ҝ�v]
�nT�Hhz٠�Y��f��e4��������|=��\+$X�3�]�z��=��x盃,m���n�{p;OC�˯���?v�&BH�� �����@=z��e4�l�>�\x�3qX�H������9��6{6i��6n}����@�Ϯ9�D�dJ2,�rh�)��f�^�� ��4y�O������&�۳���p�z��e4�Em-g�#x�$rM |�� k�x�`kw�\D���w{��~�	 l1�K���[��v�Ԯ�0 l �7���p �@����	N���ţ̻r��
�T�M�7V�x��\��8�U��7g'�PAc�q�c���7gl�q�v��9KB�룷m�GFʲ�Q�h�Zח��5��]�j��y��0��۠S�3&�VN��]Mp�-]�뗬�e�ٮ9�ǘ13�)��Ù����﻽��w�����>��D��N
���9�swRrk#OY��K��*<[��F���p.u�u��I� �ݜ���\ ����Uuz��@�����)E��4�{8��I$����{� ~�d�{9e��&��"JL���@;ܭ��'7V��, ���UJ�J���UUI�~���fl�����|�%M�g �f�V�� �N)�rp_;�?	B�����}��oK�g��9{u�Bp��>���5��)׷jm�ys�����CA�.�NΥ�V�^K����x����ޗx�����ҙsJm-M�ـ��5�"!4�KH.)Q@�u&�����O{����ҚZ"�-g�"b���4��� ~�d�I7��4�{vp�V��,�%�$ڄ�I��f�}�@;�� �r�@�Y���E�2`I&�w��p���߷��s_Ӏ�d�{���������)�d�g,�ьֹ�v2f�֛�j㎻!��Z)�cW6Mvy:�P�����r|_�@;ܬ��f�}�@;/;�I0�$<�!I4�瓚���߷��3o� =���;�ح^-�"�LJ)4�Y�{��E��'��*�l!	RP��!	J�#J�K�c	� ��bT
z,�P��� S"��"�� �1! �!�
RY	D%�	h�v��U���㘤KD�"�'&��u��- �����@:����'�T�L�!���f�^�� ��h�j����X�R7mbR��yn����X��Kk�R����unĖ���������$�O�?_����f��w�Uu���8�����M�q�nG' =���J�l�^��nl�{Mس�[��"d��M��Z׬��Y�z� ���X�̀��E�z� �U�׬���D"�:u|�}��O|פ30�$��$)&�^���g���_��@:��˫hV	F�&�M$�CnZ��܅���ں'&�`�e�e'ZCA��x�H� �L�Ģ�@:���ڴ�욒I.�75����U��m5�F��N�ט���f�� nk�����wīb�BŠm�z�4��@�;V�ֈ��Y����$�M �U��٠{��@:�4s���XȢP�)4ٙ8ҥ웯�����y8}�� m�E5ݲ�ۥ���o_[� -���M��  ����T�3(�r�kgl�wF�X��6Li[��8�w= 0�^S�6�Ź�uӱ����u:6�:μ�n�6
�<x��a��f+g[�d܎S�nq�׶4<u��7�cm�3�$v2GU���/���{�y�q���ќ<�zh�%5V�B�Ok��������="�����3�{)���睌�-*wNp���$]�^�y���^m ~�>�j��� �U��٠vr�!1�Yȴ�Y���@:���ڴ��d�,X�D�$��Y�z���Z׬�>�\xѱ�D�2D%�׬�=�ՠz� �U���㘲C�F�rh�j��f�^�� ��ho����������YN�ms�LnxYݝ�^Ԭ���k�ݘ��X�hdA������!_ _����Y�z���ZZ"�-b?�b��I4�W7��P��S@+�A�$�}f����@:����\�ˉ,a �$Rh^�@�;V�u�4�VhŞ�ݐX�1F��h~�]g��@/��h���f�}��,d��q
,��Z׬��Y�z���Z�f7��R8�iA�H�o�Ts�V�r\���d��=k�gh�6q�U\ۛ:p�<�!I4�Vh^�@�;V�u�4{�,h��"B�"�M ��h�j��f�^���}q�dJ0��@�;V�u�4���y·����5jMVSZ@��P��- (@��
�Mh��&� ��Zj�E֑qRd��H�
�Թ�h�MkFցAm��j�4�Eوrmd���i��S�h5�a�H0YC�~n�h։u����/��H��)8~.�HH��k�H0��.�MhxRE�\�5���I��@E� $�VENASƸ*�T` z�_� �<QD���H"z"'��J��N
���@
��2k?_3rI����r���*ي`dAG�u�4�Vh^�@�e4�ElZ�D�$�hZ���f�z�h^�@���n��^��Œ^n���߯7?t����%���m�ٺX:�qWz@�:�9څ	"������)�z� �U��g��d9?�j`I&���o�?��a��8�׳��d�|��K$'�(�dR׬�uVh^�@�e4��d�$$HRM �r� 9���`CI�Z��Q����f��n,h��"B�"��= ��h�M ��hu+�<����x�
YUyk4�3�V�R�F��̭��6��8%gn�i��BtKD�rh�M ��hu+��f���]�V�S"a$4�Y�Uԯ@:���S@�U������"I$�*�W�z��)��g �X7붱6Ֆ�#r�UM�sf��������@��^�س�[�	\��� �N���I�g@ך}X�����B�
bS���*��U
��.�p�a^^{X�8m 5�     ���Vב��-aR�X3��&&�O;)��7.����+�l�n��ۨ��m��7<�[�nq<��]e�;c	�J�Z�P˹xx��s�ن�����5��ݶN�n5�+�gg��Va=Eۚ�6�v�t����n( ����6�<WLֳ5�l�sVم��b�����BSc[!�AK����M���D�;v�c�X盶t�M�8۪k�Ƅx��:����� s�u����D%���~4���a�L �<�"94
����Y�[e4�l�;��ƍ�"$)��l�@=z��)��f�WR��>��	 ��NM�)��f�WR� ��4�b�J�����b.���� s�u��ށm��>��yI���X��m#�޻�l�d��;{'GS�s����m7`1X�n���p�(�dD�I��Y��f�s&���=�8m�yv֦ڲ�FL�\��'�|�7�B�Z=G�vk��� �~�4�U�b�en�,rb#sI4�S@;�� �Uf�z���g,���D�Y2) �[4�U���hl��v^�p��@C�#�@=�Y��f���hz٠UqW��<��؅��7��;2�Zh��[���!�s����=4K[L�SH���H���@=z������������{��� �ȱ� ��ٓjI%M�{vpٯg ?g�sR���ڛon�հ�"� �n� �r�T�A&�w�s�f�1���(;.2K�p6��7�׳��M�����@��.meė�y0��I��f���hz٠����������LpWa^��:������S8y��SC��T7<Y��u�Վi���	$�:�M �[4�U���hݜ��I���&E!��f�{��@�^���he�w�<�"94�U�����S@;���ˍDĒ�"jMI$���m�ݚp߳'*��-�Ə�&ƫ��&�^�䟽ם5�I�C"q�l��w������zs��8(Ƣ�K��'��"�͋����-�TV�Qóx�za2�x*��Sb.���� 7���6_:�u�n�8n�۶�e�ˌ�� �r� �|� ����㈙�͵��N�˲�����~!�*�X�޶h_���;{+vAc��đ�l��w������z���2Bd2",���w���������0y$	@��RJ� �J�1`@@�HF�!���# ���@�Y�w����� ��6�.t�M���i�� ��]6 m�@ {`7.��;v{N��W�+P���\��5�[�=h�������qN��<Fszc/q�h'T@h�h4�ѶcWv�s�	96�I���z콊#pVCa����v����n�Sv�[�ۖ^_-ٜ�ٛ�	Φ6�y�q��FW�zy�r�1ڤ��Fw_���}�=�²E�s8l�3v�k�G.�9cl�c�pN7��1-t�n�6�q�����������S@;���ˍX�&H���@�^���0����.��
ɽO�W!v(�%�w/�f�Ӏ��8m&�f��@���z�J��4�0�CCj��7�ݜ �k��?<�_ �dÀu�+b�# ��$rM٘�_���;󿖁��hz٠{�*�6����pTQ�j�sx�����m���r�$\���ᩘhz]l
�p+��E}��?_���:�M �[4�U�b�enȑ�d�5�r�]�<���o�j��
�C���k�x��9�Q	%27��2H�dDY2) ����uVh���:�M 콎��Ɉy"Drh��4W�hl��w��Źr!�)�L�	5&���������@=�Y�yuv1�2dj&�D8�����p]g3׷k�ہ��9٭N�m
Lq��b#aZ[)��f�{��@�}V��Ò��1L!�����$/�@���Z[)ͪUTٛ�6�|��ˌ�� �v�7$����"�R0_�P�P�T(QJJ�w~0���9�L�T����0 �$�=_U�u��޶hu,�;{+vD��5?��hl��w���K4W�hwb��Ņd�W��<4csQ��۷3���8�M���S�O6XvMc�m�Ag"��)>�v�x��x��87l�NZ`�L�F��@;�f���H���Z��~4�l�9[�	�LD�$@�&���������@;�f���\q��b#aZ[)��� ;�����W	(��|� ֎��|��qD���fN�O3M��;�hl��u�_�m)�������O/\z,��6��x���������]0ٓ���!�F# ��$rO�-�~����S@;���ı.˂_�LD��I�z��@�e4�l��Y�v,�V�"NLDnE"�:�M �[4��h������$G�L�C@;�� ���S@;*�2�	��"�'&�wR�]s���`kw�T!D�?,�)}�Ha7�lWX�D�dj�Ժ4Z�BHT�BP2M�H?�W�B2Ԁ�� �B1#B�%�%	x��J��ٲ��@��`�H0�c�k|#!@"0`���I�8�B��	 ����(��
B��kJ]cB��D������(�OVh�?Cd"B	!e
��$�!����B'�ֆ�JX�T࿒	a�0 A}D�#. B$]x�,
�H"�����$� B0$@�&@�m\O$�0���_t�Ow�ӿ]���������               �9wM�ݭ�]�v����[��XrW[KZ�IV�4�%�6F�F�m�܍U�I6�^U�P�l      �     �       M�    8^��       m�  �     �       �[h     ���8�M�'V�UP<�Y�vLf�`,	+ۮdX��/1�t�pΎH�$�M+�����S�q��zX2+��*�3gl���wd� �����S�PHF�9�G*�sD����l�M�ΈB��0�-��Wd[=����!<�����,r���2{Nޘ0�$���v�W�L��X�Y�gd������Cԝs���m<n�7e̻�vJ9ɠ��4�M�ms���$���N���ʊ����\v���r �d8��B^�^�%�ݦθp�pN��b^"�9�n��I6eF�-���=�*�r�s{n0t.�69S;�xV�d���1n���p�E��\牵�Ƈ6�[O�bռ[rԳ��6�Y�3u�-W\%<=�����+<�WrکP��!���.�����aتF��
N���P��l�-ۗ�(Z�N.��`��x�ָ�c��h�7>4�!1�e�0X�]�Ŗ��ፇd�x9�v���.�����B���6��/�YmJ��n��ccY��\	fq�ٶZ|���pq��7Ş�AY���l��4vI��u9�����dAS��p���\:��4�]`+j��[Ͷ&�<��]-��@6�5�A%���ۍ��6��-;۰���W� �z8�=�$5�H�Ԭ�Mz�25ţn���1����2�g%+Z�\�-�m�pm�Um��.�4@2[{d�&`,$˦�K5�` �9��[�t��+�ڥZ�`U�m��JMfJ[2�3��J��D��b��]*?� > '��?S����������_�� m�J��:�n�Mk��mt� [@�� � �z�.�f-;Stƨ1��Vra;h�Ddv��"z$�G]�v��P\����}�ӧ'��=w�d�*�pi�^��q�];Z �m�-��^Töf�j#6����F^M'�d�q���vq�k��۩�h�y���u8�r�x����q�9���f���TY�y���w^������7։:D�^\��d��d!���'��t���J�^����9�Ʀ"b	� L�@��Z[)��f�wR��>��?�FF�8��S@;�� �Uf�����%S�1L!�����@=�Y�z��@�e4�B�-b!��"G$�uVh���:�M �[4��m\IG1	"�@�}V���0�;��.��(I-v�MW�Uab�W��=���ny�ς�a�gXY܊��F)�W[�:�sN�y���l��$�٧ =����ǓiRIu�m� b̭�IRj(�8��NJhU
�P�RJ(PXO9w�y�s�sv� ��� &"d�4ܚ�����S@;����p���LA2E�dz���S@;��ةUS��6��^j���F�� �q�nـ����u�k�s��[��{,�pVS��\��V�k:"$��J�<��]�ڎ�Z&ݬɎ�Cn{���I �[4]J�W�hl��ֈU��D11�H�.�z���S@;����ڠ��LU7e������0�!%p�%T>���*����;{+v'"27?��hj��y��8�ݜ��e��~���9e����Y0r- �[4.�z���j�=�1ك&$�q(��l��������s9#���V{���tv���	7�L �"�'&��ԯ@�}V���Z޶h�˃Ʀ"b��/�~��>j�UI6f^��{vh]J��������8�z� =�2pڤ���6���_ �#��
��qR\|I&�۳�y�gu�'�u�rx��PM'�%˫V�ׄ*��"��$rM˩_ �IU{fk�����ٓ�~������Iy���_ۨ/����f���9[�v��'\!`���\���`ˮC�v�%i��?� �� ;[�g�� �+r�an%����@�v��$�~�+���W�hgvX�0��Y0r- �[4.�z���j�ʮ�b��F��@��W�z���=��|��{vp=ը��L���@L�@�}V���Z޶h]g��I9����'���@����l�ۤ�{l���ְ [@	 '@ �  hK�a�&ڭ0 �t�#�f4�+ےu�X�w$��Y_i=!�wT�	�v�����vݮԨ��&�=�c;�?}�n� �[�l�S�����;Y|���k�=2Cn�c�#GW���85��8��a��k#���:����&���۞z\�,C�{]M���:���~�����=���)eU�Mf��1���ɸS�!&vֹ�����������q��#�G��- �[8��2�����|���|��sd�- �[4.�z���k�ҪI6f�Ƕ>Yd��$�' ��@�}V���Z޶h�9������Ԅz���j����ڥI?^i��15�z��mK�QH��j���@��W�z��@��?[65�T��WKa
�&���+�Wa�^�����m�ٶ�8�C���Y0r- �[4.�z���j�ʮw ��$Q���<�����b�D4@�T-M2$d����&������
G$M*H�*!��H	�<:*OK�y��g��| ����I6y�B��L��V"Y/�y�m�z�T�l���h����>�� s�$b�C"q����kw�l�`/�`h�zcň�0�H����@��W�z��@�v��|�aI���\>������۫6�ͻ\W뚖��m7�Z�nx��J1��#�h]J�W�h�ՠ�f���Y̭,����@�}V���Z޶h]J�Ş����K#s�)���Z��}�� 40].�	(�HJD.����:�5�s����.��#Q#�jT�{vp<�o�~��h�ՠ�Q��O蒑F��@��W�z��@�v� �[4
�}�i�����^_%�0�z�u"=r�.�N=�X�r=K��=v�K�q���%�����M� v�B��=!��?=���q�A)�0�-�ڶ�T�䐩)sn�|m�?�p{%��#�#�@;߬�<���jUM�o5���|��<��c �N"G$�<������;��C�3�DD
�Gkw�s�H:L�5`Z��G�z��@�v� �[4.�z�?x�i �	8+���M�ZK��<\7=��Mr퓃���;@�sŞ-�]-Յ�a��Zs�hz٠yu+�=_U���c$ȏ�,�9��ֽ˩^�����ڴ��1��F��4���R���Zs�hz٠y[����LA1�FG�z��@�v� �[4.�z�}q����8��j���@��W�z��@����>���n�FےI�`.ܲn�um+�� �m���   hUjN�r�zvUv3�ِ�4uG8�<ltzs�.{Eɱ���� ��=�F��۶���j�ٺ��"�An����s��m�,S%���݋�N{��4��p]�8��'P���PR�{ksv�vQS��u�`v�˷On����
J��f�!؆����y�ӗ��$'
>����t�F�b��>�֕�Dn�y��x�ݗ�L�{ ����a�������R���Zs�hh�ZZ�A9�E$�<���u�p�np����BID��RV~if' �Ԅz~w��;��@;��˭zb�ev	�('?���z���[�g��]s� �ݖ2L���"Ƀ�h�k�<�נz��@�;V�}r+BmƢ�g�n�����\s��� 6���=K]:ŉA�`�4�PiǠyu�@�}V��v���z��pɍLD�&k5�'�u�zDr ��1�DI�J�h����P��
":���-��6y�ϒ�&�c�$2�L!�qh_��@�z�˭zW�hZ ��##d�-���.��_U�{��@�D*��"%�9����<�נ~����ٚ���_ ��e����f���vҖU8*]ڬz��Ԝ���lk�#Fݬ6w�4S1��u��t�q]��S���������/�`<�`�jt� �"�s����v����.�|�~�ͤ�6Y�e�(ʐ#Qw8��Հl�u�����5J�J�fBD�ˢ~Mf8�*XL9��BЄv�@��	"0"�k�2^�l�P�N!T��~0mc������$"�B��JH����x"��AE<S�.���8�p`� ���*�*+�8	D�	�"���B���k�p��p�˙)�..�n(6��<�נu}V��v�������51LfǠu}V��v����.�����DF�c�:��|��ۮ��ooi�ɞG,�2����juKh�
Lq�A)�0�-��Z+��]k�:��@��OLx�C$qh�W�yu�@�����ZZ!V����4�'#�@��^���Z�ڴW��=^�:��R �Swu�s�s�oSs�t�u�� �"�Y�P�X�D�@G����u���g��q�M�A9�ԋ@�;V������]=���b���0��*�9g��g[(M�	��nZ�<����ll���nۍY�E�L-���/uzW�hyڴ�U!�F����/u{��3�"�w��;���@�z�ˮ\2cS1�`�zW�h�h�W�yzנ}Ϯ8�C ���G��;V���z��zW�h�T�ǋ��!Z+��^��_U�}�j�O�#�h1JRYĄ!n��;x��������U�4�Nk���N�@!��� 8�`�$�}h�pڣ�:Θ�kv�2��dw�.c˷K�g� �Sq�^b�H��;�Vg�)�>���.���spwmiό�Ё�K�ێ�ul+���\��퓀`�t{��z#�&�c��z7k��2�j�s�6.�7k�k.M�/K&h�����Nj�|�0�Z���w����<����N
�\���jΖ*n���H߯����ˤܽ���:y���P�r7'#�����@����;V���z��c����"cJG�u}V����@�z���^��Y���M�A9�ԋ@��ՠr�^���@��� �=�c$ȏ�,�9���z�������Z�*��?�JE�z�������Z+��o����ߴt*�:,0��e�������4�fԹ�e����s�;WX�%�Wu�s�s�{i��:_:�B������=]�� ��/�0�Š}�m�U�Hv���y�r���e�e�5UU6fja��'���2G�W���^�����>�hh�Z�� ����q�~�Q���Հ?��8�����]`�C��� ��)���Z�v����/uz�̳pm���Q��r�g8�V�}��uk��!�t+��X(�7�����b���16$��R-�;V�������^�*]a�y����l�E�L�@�z����˯�_��Z^c�UI���͂%KnG���:y�X:�8BP���""6!%
�j�Z+��V��&51LfG����y�5��M8�{/��U=�fށ���d$2�L"X��@��M���
���_U��U���)�N
����m[�a�PV6��<.� :LGWMq�q��A�<X�� C@�z��e�e����dӀf�Ƕ�v�[���r�?����UR����|}g�@�z�ׂ9��$�&4�z:�8޶`/�`w�`�jm�s`��jE�_t����z_��[��P�0A�!dXD"�Q��$@�$DBU��� r֝�v�Ee�r�ɻ0�ΰ;ΰu�p�l�7]���Z0S��l���z�N�Dg�:�E�a3Ep�,���uBC,bMu��
,�z^�����/�S@�z��r����&0qɠu}V��t����z������$QC�D�G��t��[�h޶h��@��?�,FF	!������e�j�����7F=�˶�2Ә��M �����hs�ޯ�����?�ϒ 6�4XC����z�V��n�[� -���t� �Q  z��uȰ[Y�ķ����['�:_"-Βzobm�'t8�q��e�g{rr�4d��{,ݗ�fa���,����K�ݰڅ��v��nYȎ.�q�5����t�r�rt8^��[�=>*ݸ��ݚPD����Ȭi�W�܃�Dd�Og���]��V���ۻ�����ͅ�Iy���_����[>{9��b�-�S�ݛ���5ɛ81�=)�VD��N�����@��U����u��g��������5"�>��h�f�}�f�k���2L��Eɂ�h���}�f�k���Z�
�Xa?�JEN�u����>��h����n\ 51L`�@��Z���ޔ���o����q���z{,����^�2sI��M�Krm&v֒n�p���+;v,3�*���Fӗ ���g� ｓ�UR���|wSZ��V�b�R\|��g�BX�D*��""�w�=��@��U�u�kSA4�$Ԇ�w���3/��m$���y��n�Ӏ~�#��$b I&�k���Z�)�wY�{{9�9����)��>�@��4��4_U�z�?���M�l�/�60�]��mC�]3�<��\�p�vvm�'hr�E[։����`����9k脖�w�������F��$�4�� �~�}Ͽ-��hV�2cS2B�]]��9�w;�Ҏ�	B�u�"��P(��k�n��������H��/�0�b�- �u���> w=������|wSZ�%Zi�A���-}V�}�f�k���4��tm�F6�cIbѵ	�G\�X�Cn����q��i.�7i������aHLdI�1'Z��4_U�wY�Z��Ո�<�����$��������9�w;�5J���I���)�}�f�k������M��- �:匓"!�D�$��u�pϝ��9��$���B�)��;
�
4C�W�'M ���G�a?�ԉ��Z��4_U��@��Z.�^TG�Rˌ-j�������GZ-��\8흜Nr;OEQ�]�K�q�����o�\� ;y� �s��%�~^�S�2E1)�Kqh{��-}V�}z���h�YVl�x�A���-�M ���������:�
���ȓNbMHh��h��@=��8�R{��8���ӵ�JZ���h��@;�f�oJh׬М<__��)DRDX1H@Ѩ��D,+m�?��O�t��l��@�UN eD�%E���6��$.�Yc�Q�|<U�MZDc�|����>:�$��<$X�$dI�����U��!�֤�F!#��xAC���I4��d�(O����  ��          l�\�m��&%y���m@�v�Y\W:Jqs[����P*f�I�#�8
�*���^��ӵ�D�            �       [%    8_��       'M�         m�      �      �I����--�IZ��m���vv��HV��ŕ7k�6zT�j�lT�sN=dخ�0H�mòr]m��ng��ݗ��A2q�kf�Pq��۩�㢪��U��ٱ�B�[�\pr�`i;V���.�`��،�eň�2u�mj�G[�	�m'K�v��S���`7j���UN�"GFȈ�c���n�Z㜭��ڶ�;&@y���xN9�����OnzTpɷ3�;��]q�OgaقƢ�{mv�g�Yt��9��s�F��usqϝ�JuUvٽ����nZ냮0��k�$*m�T�[#�[s۶�Tݐ�W����=���cv�x�n�L���k��~��s��;���ĶE͖^���n�R�yD�)���T�[�E�$�]��Yd�d'SȪ�����e�P����5oA�e��Y�y�^Kvszx&�u_=]�<M���N�ۀ��=6���;O��X� �/d�hpojTk��WF՛i�y��0�<BY��`�8&vwD[y�*����\�99�24�v���v(
�;"�n:sv��t�Lkl���ZP�;a6�V�@�9����vd��G��[kv�v)$z�yAƝ��Cv7��֍v�t�ô��`x������7d+X��s�툵Pg��:tt8���W6PXT�j�pE�y��c�I���;&ɺ��9ݭ9lc�wk$h��e�I9Mn 	ugeS��i(�嚜�*Լ�f��	")�F8���m�WI�5��	��5.��O���G����� ]���P8 "�P6'����w{���ws���l���v{)�m�WUU\ �� �    ���+�];*�t�#z"��p���v{)��rբ������6"�;+v9�X.q�$��A�I�X�Dx#��tё�l]��-6�cdw*2�q��a{/6հ'=m6=����lkv��m����nJ;��kd�>ج��;�vtA����h�1Y4<�KJA \��}�ޟ����$��.�4��"���nA�՞6@��m��U��,�n�dr	��O�_�>�Mޔ��Y�Z�� �:匓	��YRMޔ��Y�Z�� �u��
�XdG�d���4��h��@;�f�oJhG\�cjb& ���&�k���h���}z����$QA)�Kqh{��-�M ������>���7�"�7����N|�N-��mgĴ� �+��ټ`n��&k�5�<X�ƈ8���)�^�@��Z��4�B�jh2$Ә��� <��\BJdn�� {y� �[9�=����bRշI' ݼ׀�� o�����R�u;.ɛ�	Q���U$��͜w&� ｓ���$�fk�嚶Y""R����)�wY�Z�� ������C�~��d�g,.ݭ�VlWe������N ��ô�0Ms��1&�ѽ:���4��4_U�wY�[Қ�.ژ��	�rh��@=�� o����y�BJdߩ�����(�.eM�� k^ �[0�@�bA`Ċ, 1h) 1���!GBQ�Uc��s���9YqJTܦ�294zS@>�@��Z�u�Z!Q��dI�1&�4��4_U�wY�[Қu�^��R7N
�rj޺ů7I��lv3�'G�H�!f�*Q'�'���J`I&�k�������(��[��R�:����0��H���7�$~�g�@=o�Z�� �:匓"?�"Y���)�wY�Z�� ��� �Z,2b22D�N�u������sr>̈́��A�� ,	 @���JZ���7$��፩�����G&�k��������n�Ӏ��p����ͽ�]����D8��#�8���9��س��'����p78��Kiv+�RYۋ�L~m���Mޔ����-}V�m�E�?�,QcD��)�{��-}V�}�@�D*=�4�$Ԇ�}�@��Z���ޔ�=z&<O*3#Ɣ�rM��h��4zS@��^��Y��a �1��)�_u��)�U�@��ZwK I*�Z���0���e|�	zk �m��� $�z�7$����ۚ����+���Ϫ���u7`����ę8��n��6}�gV�8ǒM��քB�vIlq��"��NE�C�zNJLI.�mr�<�ٵN����-J�Z��Nw+4t*c�0Pt��֭۵���nZSl��9[�Bl<V_�5lR��xn��8\��VH�y�����g[���3��`��g�U\U��l٢c��FI�̐�dB�|��~4����f_��UU��f� f�]�1L�cI8h޶h��@=�@��4�m�SLiL���@��Z�u��)�z٠}_\d��0�2qh��h���}�f��UU=ٚ��Sѫ�iƭ��\�}l�kw�7\� 7y� sR�w�"����YK�w.뫃E��K(b��}���'<K�+�8�r��d۠F੻<��׀7\� 7y� �[0�'��)�ܚ��ٟ��?�P��Q*T 7y� ����n�b�g;	���'�R- ���ޔ��Rl����7o5����%�"((�Y���)�z٠Z�� ��� �Te�LF)�,i' ���j�[�5��͜3�ט�ٗ �l����7Pv��z�;zⶍ!ْ�;��t�jļ:i5u�ڴu��I�_U��Y�[Қ������I�?�2qh��h���}�f�k�늋�1b� ���+�f {[�)I�T�D*"a%M�U��Y�u��D�sjC@=�� �s� ��x}l�5��ʌő�`7&�k�٘�����Y���l�>�2�M�m	��Q��r�g;���>��:��Z��7�$���a�u�t�a�#��K���E"�{��-�M ��ɵJ�Xn�k���l�DEK"�@��4���_U��@-a��d�I�@���@n�� v���`��(*n%Z.YwUU$������l���7'�S��"�E
>��_��Z�;�$j���,QŠ7��ι� �s��J'~R�t�
YUyk(k���%��o���Rԩ�9�U������X���ɬ���Y��>���-v� �u�WɊ���4�$�@���@��� �u��h��+?�F)���@s�� ;y� ���ι��V���A�c�'�z��4�j�>���*�@;=r�I��dQ,�RM�78�F�o��KV v�U{�s����� m����5I]o�K�hI��mp ��� )D�8 ^��2�KQ&0�u�ۘ�6��y�ڨ6��]�/I�nԑ<�x��9���:H{u�mi�탷[���
qV����׍��B���\�e��KK�3�I��Ӄk��ف6;/������k�n���f�@m�����Ӝ9��+�y͸������������������V�LJ]��cv�ړ�����]6�J<14�)Yf�z3��s���YՒ,i7ߟ�
����Y�_;V������A0���qhwW��@�v�������#��?� �G�w���ڴ��
���/�= ,QcD��hW�hwW��@��LTx�I�1'Z��Z]��{��/��@Y���DǑ45���ܙ?���r���י�E4غ�}���6��7k��Q��ȉ�?�qx��P�{���|@5w��b����k?�H���o��BR��(���"��:[u�9�wϪ�&��l�EmF9' �_��@�^�@��� �u�|.a�18�j����mRO��v��; ~�Y����m��[��a#Q	Ǡc�����{6t}�8_�e���?׷��U^Z�/gϧf���t�
.,�f�bMaj�upZ�v,3���oW%�Ǡ{��/�����@���ۊ�ł��6A�ɠ_YM��^�Wuz�u���b��#ls��0Os��s�7b!\z���M$ ICЖ(Ł @��o�(:ҡ�n]��Y�|/�1B��R1R�i�F�ڤ��[q����`��B!"�H�!A�mM�5M�
�Ev������-�B<�@! �̈́9���ͨJB���)� 0L EBh=xc�*�(@�h�(1`F�e4<�� y M.��W�#�?
�D?1��: ������lt�1�t�
h!M/��H�	ȏ��kFyJiq��}M��z��	��F2�j)�f�J"��p=|G��~D=S �����P���*���Њ,g�w��ץ4^���"&��$�@��ހ}�f�ץ4�uzŞ�w$��c�'�N7�wY�u�M��^���o@�x��$�pDƐ)3(��;V8��Sێյ���V+cIg��n�V^ne��I�2L&C"�dB�hzS@�w[���]�%��͜ �	�f�D��X�'��^���o@>�@�Қ�ۃ���F��@�v���@�Қ˺��v��d��Hހ}�f�ץ4����? ��F���V��t#�� @�}�[�w�K�Mo))�cd�^��>^���kz����f^���l��ډ�%��Fծ�;=r9�4�����2cq���a��nx���(ŊH|�_�@�v���f�ץ4��ƇF��F)�9��M�`�w�s�f �[��Z�ܓ#1�0��8ހ^�4�)�U�^�k�� �z匓"!�D�&�����*��@��ހ^�4���,2f$X�N�h�[��f�}e4����.��I$m��Ee2�{c`�ų�B0 �� N�J$ ���-�k�j(	�6�&�ˉ��AC6���z,�==��Inw���g����ѐz5��+¼tM�k��� �+m�Msaa�qtpmuM/�ɤ���#U�nt]3�b��W^8^{A�]V���9M�+\�;�4#;
\�����t���kz�pδ���-��i0���{i7,�6���#���#,���ь���D5��cj �H�D���?~�7�����a�%Iu���_ ך�Yr��2#�= ��h�S@�v��r�7ڞ�_#CRڻ!v�}��_;V�k�� ��hW���@�1(�4�j�-v������hu�J%���P1��k�� ��h�S@�v��إ�0SI�XE��N: ��9qp��t�vK� {u[��39�,�nn�7T�,mzp�;��f ���������������$ȈdQ,��&�}e5�?����\%�"!A��<��n� u�|b�3	�,i'�ڴ�̻᪩�s6p۳N��b��œ	Ȓ�h]���@��M�ڴ]q�8̃�S �I��f�����h]����c�[$ʇ�9�z1qv5�P�6e�6���H;xo 7i�&���4v:N]e*�m�l��|�Z+jz{��>���Q�
b�Hh�S@�mO@/u���hu�J%���S���5�����Q	(��v��h�<2��F' ��8ހ^�4�L8~����I<��w�/jخL�fEȚrh[)�_;V��ڞ�^�4{OVЛq��Kb���ۡ�"68�6�q\�Όv��u܏�AU���ɘL�cp�/��@�mO@/u���hgu�[��a#YR>�˾j�M��l��f�?^c��㸜FF�S �I��f�����h]���= ,�cdRM�e4�j�:�[������T8@��D�T ��s�ܓ�5�x/�����/��@��o@/u���h�b�(�jF�m�J���廮1k�Ƒ`�t<�⃸��#�L��b)��J`4��:�[��o �v��78��'M]�Ur8ހ^�4���/��@��o@=��c$ȈdQ,��&������|5&�ov�����Oř"���p5$��n��{�| �{' ��M��cksL"�#JE�um�`�w�y�f �������d�lu�7nY7iz붝3��� 6�     h%J����%�	%׷4�Ngs���(1P��������ZǮ܂dz޺�^�9�:8�j�f�!mհ���Ll�lvj6�ª��̉�ݹNgqn�6�����G��ml�����g��=��s��a��1�K<�+v�˷Nۮ.����7M�y��j�O61@q��U�����B9㫰�n:�u�u��[y���e�,��C��JL�l����r�k:�/Pހ~��h[)�_t����ށz�ǦLY��6����h�)�uv���f��|�
��
b�Hh�w4������>�S@�cN`�b%� �"�|����۾ }���<ݳ {��V�M]�S��'��@��M������_�߿�����\�$J��Y�}p3���݇3��Z1�q�8���K�g���k"�D�&����h�w4��������ɘL�cp�=��7�E0S�EsS��ַ$��M�e4��፭�Y0�,�93@�M�`�w�y�f ��,���e�.�Pj\��$�$��6p۳�_u��9[S�/\TX�ɋ#X�ےp�L8���ٽ]���Y�\\�ؒ���k�mA�ܻ�]����T-ñ��x��1�掞� �b� SjC�?u����= ��4���>�!b�K�4��:n� ���0�l�5J�髻�������� {��7l�����������f��]��,�&D3"�dM94���/�g �^e��R�M�g 7�xY�ɘL�cp�/��h]���Y�}l��U��+&D�q(�A�do.����������%;fm&���oZq�T����Y��aYrf���ހ_u���h�w4]q�8̃�S �d�h�w�sv��<X5M�}
!%2}g��F���&�~�������@/�����Tx�A�n����(J_SŀsT����g�JdYYCB��� H���FTa�h�J8�b�# �H$��ֳ��7$���,���F)�#����@/��[)�^�M�fY��J`��E��Y��%ӹn=�[��sn�8�SG6��\�Xb��I���O�o@/����h�S@��o@>ιf92&�(�Dӓ@��M�Jh]�����T�o��`�R5�s&��7U�[���0.�U8��Dq�ww��͛�| �n��ɇj��I=��j�e�.�Pi�.���'�I7v��۽��������krO�����U�E_��EZ
(���(���(����@�������
� �@X*T��H*Q��E��V
�AR�E�� �D*Ab*`�E���X*T��"�H*P��
�A`�E
���E
�A *���� **���E*� �EB"�H*@ * �@��E��H��R
������@"�E *
�B
�B�"�����D �@
���@X*P`*`*Qb*�� *H
�@��E"�F���E��@`�@H��Q��@R�
�"*��`*V�"*B�
� * �F�
���A`*E
�U
���A��D��B�"
�H
� *�����F���"�@��E��2""�U��QU��QU��QEVtQU����QEW�E_�EU�QU��QEW��E_�QU��(���b��L���^Z6�e� � ���fO� ��~  � �@     U�4( � �� =�       IH
TT�T�T!��P$T�U*"�*���� ( �ER*$ 0   �    ��f zQ��V��帳�����������a�P˻5���|�׶�]r��|   ��W��{��� >�������<��a�01hW� �޽EMu�q��6�Ws-� � �� h  ��0 <z'����p�qk�ړ^0�i}�pR�r�[4��ʤ���_<
)�����8��3��/y�uU��
0���{�|5���˪������(�ON[�^׋����Q�wi^� @ �*��)��_}�������P� 4��R���Ҩ� ;3���� ��JS�(Δ���
;�  .3JR�A�(�;��v:R���4��R�3JR� Ҕ�6R��6R�R�iJiJ  p
   � �0(�JS)J)�� S�:;n��*g Q��.�i�}�}���ίv��>pʙo,��ws�n^M)�������T���{m��Vv]y<�O_ �K'�Ó]��>���y]x��
     �0�Uϩ1��i���NMN�N�|p ｦ���m�{ʧv������Vp���ˋR�5� Ӗ�׼Y�|xP���S˾�)��{qp���|�z4s�d��y:���=xN�>�� =!&�JT� ���jf�R��  Ǫ�DҏQ�2 '�U$zJR�  T�Д{T�SH  ԕ5@�0�)�'������/������f}>Ͼ���g��_�Y�PUt�
����_��*�� ��@TU:=@����)\lѭf������p�Y�[�h�,�B%�o�8�B��5��<���7��G!HL������c���􂏛���Iz@�.$)��F"FBS4y���C��u/5��|C��ϵ4zW���>���]ᴉЍjE�d @,D�B�n6�-֎8�B�"@�@h䍐�֎�%�0�H������$#�U.`�2�, ��0s&$�%�`�X�5����2�,.�3�B�虻�+��j427.9���[�ljBv�e�;L	@ H�,��]e0�
�9��#�����_O�����c�C��y�x]��� ٢7!\B�]q�۽����5��R�g�,Z��H���Xkr1�6YK�	R8D�C%!���)�o��n����8���OYfka�l���������PѮ>e7�8Y'ƾ�N7���ўy�r15Ϗ|<��y��3z�8]��'<��B�x0dB��!�P���`B����;�ձ��	����TME�M�}3<�6��D�4��B	�.n�J�*&)�:���w^2��i4�A�2F60��4�r�Ԥ���,����$K���Ēg\+��0cI"HD����w�\M@�`B�=�X�$ E�!r��m�����q�%I �b2$']O��IJ�2GO��
�*F2bB�ؤ��$����m0�	`�ĀY0=��D0�6�	���]j�L��H%$�vl���T\�Tc�t �/�q�0<�J\%)q�R$�A��`�(��s{.���0p�	MM��S�@�&%8�!��N��ym�6B�xbe������$�*h7�;e	 ��F�1�!aE���3Gj�`�X�%-�5k�BD(I��JBȐ�) ��ĹD4RF����	,��4G@Y�Đ��R@
�41tH�h�,�$l�ġ
�<�0+��A��"B,g��l�ن�xy����)�����9��o��Q!BT����s!\��Ɣ��F@p�p(�eˬ�1*�\I"D��1��˳A����0ڦ!�xp͞�o�ߜ��)�{0�m�*�#	�.kr�s��.��k�¤���[󎂛j���1�(�*��4�b7�aM�˅�cW	Lh�YJa�0ر��i�	�cE#��)X7>TSھ0��&]�ﯚ>�����q��"T$!Cg�q��3F�xq���)5�����fh���A���h=��o\s�/����_����!bR V�`h���;�a���:���s�to��3A�͗d$!LD��#���t��7ŗ����I�����
�<Ԝ�:������&��/$9Cƍ	�A���!ZD�8�6��o!%q4�aW�Ai����8��s!F�p+����P�
�M�\.h���i���H��Je0�>�B�^{��n�(M�ɞ�|y�i�S!>r�vp8z�@,���I$$ ���b�r{��w-����4a��&��>�>����6'�� Q����P+����+���X��]������aL)�d$� ���B/#� �0ӆ�xh�,hH9�6pׁ�2$$�35��8�a�����e1ӳ���$���x¤+�'����0!�C�j�(B:���{)�0,��$u%�1�L4�$Jc��b�d� ��@�C�"�J䆦�B��gU}Σ��(O����_.��2B�*��Ԥ� R����$76O�\A	��������B%��b580�ĉ���h��!L4S�tB᫚$bW4\�z�a�4i�SL#	��jɤ���ũ�+5�}ߔ�]�2jo�_}o��G����U|UЖ<Me����Pnz��zg��9��jo9�r%6�L�6D�&���(�aL���;��E�ī���1�ks)�f�7�6�Ja��B�q����sn�'�k��Tx-�] H�B�����š�'��I���#�hă���F�IC�1�bx��f���P�w�9����.s�>{�)-1>�ĉ6B-B��WmqM}�Yޖ�N�[S�~�\9BQc�\L@�)
d�h���ϳ��4�5�"���Ͼ�kG�6�o�}���|�0g��zs��x|i Oa�#�f�K
f�T\�RC&*��T/��u"Ջ�v��0�%0����}�xK��6�<I"CъB$BG \� �\��4�\3�i=���2�5^g������=4L4�O	$aSĢR�,��(JQ�Nx��5�3^$.�Ä��>)��>cR,1`!L�`T�4��"�$$�9��tqPӼxlq �0�G�D�:����C0Ѵ��qѰbB�� 	�&�E�Ȑ�#VA����A���#F�ٳA�&��<!��,a$���	'�E*��)$$*|����P"i## ����7�ѣ�U�6�(���B@!$�+ �5�@�&!�T�B�WA�D��������^.��P!M}H�~������\�g�8
JG QĊd�G	1��Xf����L��ĪJ\�!`�$I#!�p�CS �C7v�@���"A��.�_<��͘x�H;|�6aC<=#�)�hD��n[�p㰌�C&�|�9�/�0�.٪n�%�DbA�\
��b<|!pѻ����э\�ą04�*��P�R������+��o�����N	� �l=`�xl>���LO(p�f75���O'��y�������1�!}4��h�/��7�>7 �=�"z�1l"����3k���G	W�RD�\*��АZ��,gjo�"V�ߥi3L��
�B��槾��,by/����K�rpɻ�u�Z�E�� `��C�sz�#6��v`E���I�d�\��fd�L�l���8��R�6���5$�f���7S�)�炨�Ņ$dH�p�]��(B��:-�:ɸ{���N�3����M�0� Cp�,caF4|u7�=��&�zz=#)$  D�!$D&.�)��уWS|�V�f���J���ٵ�ͿI�U*)w}M�A$��ā@��FB��o����]s�Ìn;���e��p�~tz1J��T��A�Ȅ�q�ӳ��,��f��pѰ���ˆ�M��14�H�y����!�?����%a58$dJ�e���K�:4��3<x�C!14¸B&��:�Hx�JC;
f��4�4��F�:)���#L4�Za���Vsg��~y�g���^x1��8�sng��e��X'��C��6D<|M	y�9�����ZF`p9���h�e9!b����T��L#C5�����7�Z�gT��]:؀��8��je�I%�` �̶K�����m�m�.�4u�kjIp d29fu�pj��h	 �m�                          �                                                 6�                     ��                     �               >�          	    �                                                   p                ��� l  	4P                                                          �        ���                                           @[l0��m$� n�  $:��kX@�`� �`$N��%��n�L�G m  H5�A�m�  kX �M�M��	5�@ R���n]n���Ő�s���'�LŻj���6%$6�bl�⮷$8�ɶ�3[L�pS���M@m&���UUT���k(n�K,�T�����v�BNm&�m���B��D�[O; ���$�m�����I�T�:�������m��f�ٶ  ��v���%v�:��):S ?;o��l�Ͱ  	y��΍jۜ �KkEl8      Kh
Q u�v  -��[Kh5�k�T�U�,�ljeUv�H1  bCm��[M�����8]6m�m:@$-��i  ����� 6�.E�W��K.F
�W�����m۵�8.���� �l�鴀 �z�-5u/;Z*˽���(01m�H���𷭷��SB�W��S;M�TFB���`,��;�Ӓ^R���Xưm�mծ��Ӓ�h ��6�l��8Jv8ۈ���U��ۀ 6�6��E� %��Ʒ��N�9#ml�i6UZ�Wi�Am͹\k%��yyXN��M�V5�*�U,���j�ug.ˀ   l�3��㩠��lٮYM�Y]�8���Y�N�)�u��lۀ��cr /P
�ꗖU��UT�.l�m@q��oi�l�J�m��$��6ȭ�gJ�ʁǂU���J�[+�~g�}� ��Tb�n;c���UJ&*�Wo�*�Y�mJ�<����-�[4���Km��) ��U[��[R���s[@-[Z֑�()h �dh�����V���)P��
%Xㄆ��6�����+��ۖ��Z��)yj�FFX)-U��9�^P��k[�$�36ֶܡ�m��2�*�[J��	6�]av�m� [�ʻ�q 9%Y"ۃ�F�ʭT����T@� 7X+j��d��*
���V�2K*�N�U��n�2No��|m �*�T Ȗ�!������askml �IW%�6[vRBZcmf`����}N�e�Zl�[Vԙ�h����P%Z�Hv��[sI�6�X^��0�޶Ϙ�h��I��-�! I,��	8Im��`��}��Ŷ�@�WUl��7!5U�*�ʵUKf�2�[*ܓ��j�����p5U�*�4�6]�J�T���� ��K�ß �]h�c�!�pOoN��k�v�J;j9�՝:\���Ju��cb�X�[� �K,�+�L�4���Y@ m���t� ��n�T�I�l3�n� �q����]���
�L�c�Ԭ��@[E�6�`��`���kn ���i7$Jsjڀ2,PS���n�k$z�Aöض��(l	����m��v�JgCZm�%�]�5���`$9 ^�a��[�Y[��l� A6��j�i����Vՠ(i;vm�lm��8$thūd6٥N��m�v2l�!m�[pm�  L�X`�  l	e�CjZ�Y�nZ�e���VT���6�  �t��e�   5ї���/*ղ3�E  �`R����  ����ut]J�'J+մ�Pm��$� ,�"(�f�l�n�n���ݶ6�r��$ 6�w6��06�bD�[��ۥd�6C>���m]����i���}z}g�'�ݰH6���x۴��P\;�]mjݠc�%�Km��鰶��mf����)J)U	Rٕ�gF�԰T���v�[v�y@iyUj���|�\��5U^�y���8q�1�����G`�t����R�UN|�pv�UG �������iA"cY����1nGM��B���K�z�n5s͐نÉ���>Z-�v�=UPx�&X��z���8���,
VY�({=l��v�@�l�:�Ź�ʕ���V�v�I�&�L�hmŬ�'4�<�*���ښ�m�e���hYHjɮ��[-�Sݵ�r��zZ�uV%ۛ�m���{9<� �sZtPZ5�C�n�ےm��kh�y�x6�` ������w��Y� �����^�����BN� �f���`9�����"��J��vǬ��nY���A���p5�Wn�d}]RʱH��VI��/Z��hH �-U+��j��W�X[$�$��ې��lMac��˶��7�J����j�yvntHmT��R�;K�lQm�m�����X��]��yU�N���A���8/i��M�mm�,��N�v��������]�L ����n�[kC]��Q;nܕVՄ�C��[TT.��a4 ��MUT�mv�6ڝ�f���$m��E�Tn��5+*���/[f�v� s��t���J���Q�m�6��!��U�R�ʰ
��Ϋ���@� m�[vٶ�����npn�� 	��bKk���m���p9�i3�  %����/E�A#�w���m"teK쭌��@q�ېj��U��Z�j��&A�i�X������� �Ҩp�F�7W=@��a��#�8U��5uUH����l �e���-��P���kR��� ��K�9�Uڱ([�5f� 6�ٶͫd�	 [%	-+ci/6om%�HH-6$������ �I�ɵ��;UK��Ү�j�Fط[�$H-ѫ  l����c�(Ff�y�:�'e��h[dN�@����j�fQ���j����r��� p�$�ʤ)vjvV���e^�tr���P7f�7b��\�W6������R��UJ��[@  � hH�۶�IBKz�! p �ۃknζ� � �  �7m��u5��> �i�6��im[E�6큶� � �	��H [@8;m� %�$ڳmځbF�i��z��� �e��l��"\��  ~�-�( m� ;m1��(��-?��ͷ�L��E붒L �>-����[yoPm�$m�l 4l�[@ 8 -,:	٨�Z���ri0����)@������(l6� ,���n9���m,��z�m���b��km�@ 6�m� �ly�l7Z��錐�  ��h�ia��Ͷ[B�#��A�m%��U�
EX���,��eI$i8խ��M��N -���y^Um�P��KUUm�h�j�:�*\�@��Ͱq�$:�z�F�ۇ;;G��ڎQ�ól�7Q�c�b�Q;�6硷h$&ږYV��j��L �V]����v����v�I4q��V߀�u�sZ�l�YE�����u�m*�T�P�4k�@;m�N   �Ӭ��͔]Ɨ�w*�2�\�q�kD��[���m&�Jݭ�� 6�8 +���� 6V�յS$UR��l��WJ�Ad�;�� ��M@+0];f�m��(u� d�i�	6�m��J�4�H��[z:�g�� ֤�֎�d���   ,;n�� 6�������g��m�7S��Z�����Nf����5vζ���$p    $  	 6� �Z  6� Zl�]�[%]6    �`e�\5�� ���ݍ� ��Atԋ{{P�F� кl/[m�v�m  �`����p�m�А 5�H�}��Em��8l�  �I�kk��-�kZֳ_�*���
�o����*�?���(l��F�����DV����Tң��@
��|	�v���"EI��� �h��O�@�U|sѠ���U�� DZ����1V,$�XEa��"z�p~�	���)򁀆���])�\�T~7A�0�v"PD>@A>!A�@���j�`#�搞 ��E>Y"�� @�"0H�2�1 @��F(A"�`�X`B0"H� Dc�QO��P �B��HAB$FH�`$ăU�P,h�#�, �}�DXA�I�B)!�d"��1 ��Ry�>�� �ĄH
� ����P��H� F"1�$) �j��A�E��� �CJ)�R��XU� �U�I#b����ਛ 
����S� �����z���x���Q�W�_ T>V�> PDӤ��*�*`*jG�E]��(*�Q��TR {w{��{��*��m��d)T)f۬�(ְ    	     $        l       m� �h            m H     m�     �`  �     ĲT札��ޘZ�'C,V�a5�F�^��4eT`w<[:�W�5�1���g��f�rnG�T�q�CSUT����s�B�*K6�d[�Z��)��#N�L��4�f��뜯f��tu&nq��p�l)�*{��f3�V)uUv��[s��}�.݅0`;:�f�lOn�1�b�`�k%�v݌8�<B��h{n�=c;�1���M�#�Rʄ������K vv@qqBfx�+ѱ��1+�����a�b���v��kn���Zv�]�rN�����Z�.�B�#ۖ�j�z�,�p5b�����xb3����\�:Ca��vy�/�;N�(N
��&�c(v� u]-��c!T�&�=��5��C�G,MwV���>9Ό����0%�[M��H��^��������7"C�v�u��n6���z�����s8�ے�v�)��ZWE�m:�+��U��K�;��\�U���	v��롧g�]vú÷:�a,1�r���mm�&J�NO66�n�gz��=1��c�N-#�l���"^�sHt�#%;sc7\[���vC���t�۔v���XE�&�1�E����Ӯ�����dӳ�bɀ@u����!��A�C�h�[n��h+���8#`�Z��r&��UY�ZAl�q;�-b�ֲD�,�w5�5�n��Pr�؍���+\�U+)��Z�wBdX9��8ཱུ��r
�N�O]�Cm箤0\Haڜ�g��rF�k�9ڍ��$���e��fqi�9ꠁ�[;:W��.��A���t�ė�����5m�	��0$�k�wL�8��n��!�3U�n����|�{����C߅_�����A:�U��Q���)sZֵ�I�kZ֤���6���m��  m[NvNWf�bu��҅�������B�����%ی��wZ�-���v���W��7r]�; ��sn&�V:L3qv�(��&wMr�[u�z�RM��dF��4a�+i:�:A�Nl������M�vqX�#�7��$����4�Cӌ5���v:����=��w�{��#*ga3��=�c9�{&W���d˗�S���r��o�a���k��C����|`��0:䉁�)B�%)R�K�$�@���wJh��@�[^�sލ�,���D��	�@��M��0=rD���� �Ԓ(��*�14�����+k�--��;�S@�Q���ƌm�$z�h��h�)�r��δ��iBD����:��)��x�p֎�8p;�y��� �<�a�)���FLCN9$�--�`wvA��$L�L`oR�IJ�AB$��+��au��B����w���--��<��<ɐ��Q`u�d�32��otݵ`fd���cx0��?'#�-�@������"`uJP�IJT�n��M�����4Vנ�f�{�U�8�⟌��"D���#���6�g���[q��yٹ�4X�PQ��!s93@�Қ+k��@��s@;��نW#ic�)"`K�BGL	ݐ`z*����N4cmI#�*�נZ[���?~mBI������ɰ���f)����s5USa��V�V�^fM���^��c��1I�0d��^�\�0%쉁!#�D,��,�%�icq�s�r�I��+pں�����Sq7/;b���1[��"`K�BGL	ݐ`�:��ǒB4���z^��Kw4�)�uv�����H���%$��e�;���I7�;��7��`_��C_�d"Nc&h�S@��6La��� ���Ԓ(��"�E�Ń����D����wJh�"u52E�E188��a[ ��u��@��m6�s�_I4��*X���>j�n6D�Ki��|��-��/t���ڴ<�긋��rH��#���0:)-�/dL�R�)S��X���Jh]�@��^��,���yAX�2c1
C@褶��0$$t���8��NAJ�US3Q3T�fM��	F��x�ύ��h޻�mdrI H���	 �awM� ]6 w6�^@6�:c�%�GMָCI��������S]�-��e�R�� Z����f^0�ep�H�;�����l㣖�G��|:�wNfru�[���$��ݲk�ɚ^-���α;�s�\Iv8��*��6n#�:��i^�g/B�݁�n"M�庒<T��A�$\V�U�8����w��+A�H�7�W[<�Ӑ��"�d{uYW�N�x�[����k�J9룒��'\v���o�����{�4�ՠ�f�{�W�7T�&�X���3gu��v�Kw4��m�eq4��8�tR[ �&0$$t������E��cm9"��@��s@�ҚWj�����.8FLDNI$�$$t���E%�	�cJ]/E�U�[<�ؔ�N�ۣ<4����6���NV�#����;:�Ұ3��,��; ϳ+b"#�7M�Z�<��&
d�2b���ڷ�f�%Z�P�RBIB �5B����(�D+�ˬ��w-X��h��0xI�����Z}�h��h�S@��ZeǕcV4H�`�E$�--��/t���ڴ�l�/�z!��JCRc&h�A��Ill������\�ku	u��g��Z�i����
d	=��J��<�<���l�g<;`褶�&0$$t����T��ȡQ,m�$Z�h��h�)�uv� �?z�"�d�D�cBGL��2�����껸���,�=�ucw"�,!�wt���ڴ�l�-,���<��I��ɈRVנ[f�Բ�wJh��R���"Q5��RѺ���ϵ�(�d�ȧ)N�Y�p�L�3S�T;8I���6�z�h��h�)�P��5����J�/h�T�Ҥ�&�r��wd䉀zI��z!��ғIɠwt��U���٠r�٠��ن+�51���a�!����ۻVr^d�|�\/ߟ>�hםF�E�"ƛ�G�yrD��D���\�0;k���2���ٷ[>�g���-Ƀ|�=�f�^�j8�%8��+]x5ͧ\hJ��m?+��0;�:`K�&�H�)K��D89�X2D��;��h[^�ⶽ�V��yB�&% #�NS\�0=rD��D����Nܦ�J*�73J��M��(���ݛ6^���rՆ�����́�T�d�'$JBb���@�կ@���h[^���^�fg�߿q��$�L�l� 8	  �  7m� m� 8��b��n�a��	�7;{d�;<�A�u��]�]�8���n���1�M�6��.�y�=o����=���sV�.����6�]�;6����%��F���rhJ��n$8�;��d�:
��m]��V��42[9����"��Yʳ�Z����]�� ���h�zʗf��gs����������s	u�Xذ�>v�7	�:;2,i��v��
2�qr�5�	��!�)1�8�����k�<]k�:�k���نW����2�Ǚ�~I(l������f����V�����ȱ���.��]Ș�0%� �}�,Xb2ʧ.��l5(P�i�́�͵`c�ɰ<]k�=����D88��'��tt��$L_H�Ș��w/1PBD��ny��p*��#W\��`{v�,��m��P�i��]q��a��	rD����\�����qGKMJ�U*nf�S�����i(�T�&Ί�Lގ�䉁�>U�2�H��I�ի^��u��*���ֽ�{�WRғ��@���h䉁���� �)$QQe�F�ŎI�Vנx�נujנ{�w4{,�R'ڎc"��C��[[�Ge�lu�<[��s���k6�^}��Sv��N
Ba��G�x�נujנ{�w4
��@3���*�Ȍ���zV�&����V<̛���{����Zo�pp!�$N=��s@����6�=[����"hD$F0#A�VYX��X��-�A)Z����>t�SH}��6��!'��H�!��,�*��&\�yc���a
�ѣ#�Ĳ��@�h@�d��HL��B�"b�D���Y�����@aX�%˂r1�����Xȕd"Q!U�ԍ@�<�1��{d�B���E�@�ƌ!�
¬aѫ�!4j\`ef`bF��F��`�ģ
 Č"c��ֈInS.�R\�IxJ�u�㰸�Sp���L�(U�S�H�cc@� �c�cvK�n�����U 4֮h�0�1&c0�4F��)�*B�$h�j�@�.�"ck8�s!B3.eX��(G��c&\¤�)���S0�"���d�7�<Uv�hAS��b����<�Tb*DES��D!GR�����6�/�6>���Jd�c�	��*���ֽ�V��빠^0븱��L�nc�G�z�D��D����.H�C%�L�a.���k���N��^�C��V��Μ�7Omg�9���Jj�<T���D����.H�U}UU����`_�b�Ĕ�4��$��=Vנx�נujנۍ��!��ʺY�L	rD����\����ց�yr��G�4ܒ=�ֽ߲��nI���rS��"���8�ꪯMSɀW}�,T���%x���WH�.H��,�p�YhZ�..V�`nu<B�ڥ�Z�����㥮�c�s�e��r�3j�ݝCM��{��y�6s'a(��{�`{�>�ĦLC&!9�Vנx�D��D����8����J�����Yy�������GL	rG�\���ĩ"Q�/đ�Z���:`K�&����X��e�av����fZ�6I$�wvx^��V�����v��(�rI&H � H ��%��  N+��ʑ�l��]�����C\�q���0�[q'6�D�r����˽��Y[��E]���:�\��N�vƪ��OH���]�t��3m{tnu�=D�����Ɨ��䅺�a�2�vv�CRǵ�	��W���h�G��;v��-���JG�u�Tw79y-֮j��]:̶�\޹[�Wjq����5�m��ss��L��٘�R$��G�iLNG2�Ww�@�^�@�U�@�m��<�.V�#���f��l�s�(�ُ^�X��VVנ���*��b#x��@�U���#��"`w)-����JT� C8������k�;��@�U�@���\ĦLC'Ṛy�6�̭��1�ݫ�̵`b���+%������χZ��b�r0�%i��[s��sK�H4���:c�m��;(��K`u˓$t��$L	[��S��T�M�:�`u�̫�K吔|�!]���V��f��g1��ID6gL,C>�s �pi'&��}��U���ՠr�٠n6�+Q�<�uSJ�T(I'���`fN�:��U���wx��V�r�uLt�r�j����g1�^_����W@�߿Z�1�d�g~�Z�!"0�z�כ���v/�Z�k����s��L��H�U[B\S䏌�*U1T�u4�_��Vٙj�Ǚ��0���h�?�7�L�$`��@��j�zd���6�����ǙV}+&�ĦLF9�73@����j�s����@%V#H�@��
р0 �Ѐ��, ��	F�%�ߪ������妦QT���N�T�yBP��)ݿy����>��V�����6�D�)��U:��Zc�v^<ʰ7����5�����Z.�SR'�RF�Q����d�6m�;r�gn0T�6G���#j
�m���;�2	GI9<�����k�;����_/��~�f5�Ʀ7#��c�ɿ/Dɻ>�5���`}���В�S'}+��SN���T�5US`{ޯ^<ʳ[�ݵ`k�ٰ�w�<d�R�2�A�'^�X���y�6;��,�N�3�J�U�i�U���j�ճ���7v��:��U���ǂ�#	X�E:��s�9^z����<��F���.$YM�߽����Â���\^�́����׏2�8�wvՁ�0�n,L$�6�(�z�S~��W�v���V<̛����N�eS��%��4X��Ձ��j�(�������6���`w��I�M*��-���؇���`k�ٰ32��؈�;^~�X��f�F(�s�L�*����/!{����ޫ3�j�_vs2ۮ@p� v��m�,� M��x�J�4��n���o'c؜��䵎�@tOE�M�ͺ��ɺ���S%WU��'\�u����v��!�f�ݎ7.�t��6����n^�l])�mv�9�zv͡�u�9턩.[��XJ�u�P,b}�O[�݇�ftA�h�s��]�ѫ��'M�����������E�wHr�=��/W��߽��.���%�G$\%=�+v���x^���/� Q��lq�����[���d������!��4o�	���nI�_��S�*���߶u�)�X��?{�`�vG�MJ�əTX߯�k}"Ea�2~���7$�}�M�����"!z!@(D(D2g�����J�U�i�U��o�X�2l�IzHI(��{kŁ��ޫ�J���K��5c�m���?��.~��ޛ���`u�̫�^!"S�o�V�G�hNB�Q34�:��3;XX�Q��v��m�fM����.�K�rItOg���뇃\�m��ͥd��@ꚅi�1�Y����|럈j���~`ǯv���gs��m������/
_U6���m��t垆��n����۶߾����|
`�`�苮j��W�v�o��_�m��:�w�"L�o����|�b�1���<I/���$���s�b!D)���[N�m���s����VN�.MD�ə�kYwm���T$E`����߼s����^�m��38����P�D	
�~��[m��k��ɠ�T�3�]js���}u����P�A��B������>��m��2��o��-����ci�-�u�i�%f6�ye�Y2G*t]�P��NV������������:���$Ӛ��m�{���o'2��y�xj���Q��m��ש�m��[��I�TȚ�3K�m��˒�D$��B�����_�q��|����fg9����F�&dsN3RI}����%ΩbԐ�Gj)��/9�~���9m�����������?P�#�6�����~ֻ�v�oww��m��˒�{;��9Ē:�h�IQ��NE�$����o�/B�_���6���~9���㬧m��c���0n�.�u�-b]�ςܝguN��7\��95!��»<�{��n������FF�9�H�w$�����ԒVݧ�$�:�&����3�J��+��2b�I&��m��f^樉�x�֕m��wx���y9�7������ǉ�&��S̃�9��Ǯ��m�����=�3/gv=I%��oǞ$���c˓�1�4U��%�J����������M����~�嶻BB	IbR"���-B)V��$�0��C� ����K���N
bS&#����7�2��m������|�x�֕m���;��������B��C�۞�`�Wg�/�ts�\g��p۝vk)��2�������o{y(�����TL�'NiOͶ���|�m��*�m�ٜ^^Q�BQ��o�������}w����h:�����XU�P��I%T߳���l��j��o��߯9�O� ֵo�%��?Y$�Hpi'	�$������$[w&���:�<I.UJMI$�ۂ�*�do�.�is����B�D(P�}�|��m�k|�����XU��!(�(H��U{=�q���d�s&LS1�ɩ$�N��W�E�0@�����׶����Ü��3-U�ۨ�L�@ZI��� |za���P'�y�x��V��l� !����OI�"@�!�=>X#0$^�<aL4P�A+����3��
c�.�,�r�<Jh	#tj�R)�H�%�O��V�R���0�$3o)*r��I_�}GA����yI]�)��|\S�7t覀׋���p�����K��4I�f9��Y p�kA0�iD�>A��#;�R��h�>��hHF�x{��\Iu6Ra���D6�i�~�{�}ݏ���[mM��T��&띄�    	     $        l         ��         �   H8     m�    �     �    m��m�-ӗm���f�����>{�~d�vMre�̽�F`x	6:�僭�*Z��^�sMQaQ�[!n-t�-[5˷`�t�[K& .:nz�(IqtuUUJlO`�Pw)��;OnR���J�]�G���C�S�����j�6�ڻ\,&�����ģa�,F0��� k]�`t\�������8W��9�ms�.78��K.��8ǚ�n1L��8_Tz�bɷ ���vEz0�R��_*�w��݉s�����e�������ݝM���/�v���O��Z�1q�#���v�ni����<ܖ��oWPͣ�t�n�+;-�'��0�7l/� m��5P��[-���J(�:�y+�ϒH�kuKU�����H�ŏ��&�mg)=u�Y���I��@v�c��1��86j2@�۝��:,=rf��D���:��K��콈�K�m%�97&�N� f���!]�v�\��k�r�pГA��I㞜Pu�c	�n�:��q�S��#��j�V����3��P���<�-]u>.�0@.��%���	Ӷ���T�|��\� 㪏���Cě��=����]���9s��Vd��+a�:�+jɳ(q�׍u��b�z�xV�5.�5�y�ݻ�f�� Z���r*�VR�� 5�rj�-�k��5=��v�+O�d��ں���Z��;�^�����u�s�a�Pj1�R�9��͍��ywkoJ�u��dꥐ��M�v���
��R�:�����u!�D���b9��B,Z��������h��ٶV;]�T��V�-���6��m�̑2@[e��y�U�j\�n����y~��� ��@�(TS��A�D=V<�}}�{���;�߷Oַ��p� $ � �l m����K�M�e:5h�ZT˓&����ϡ�^����n��XWY�`'�8���K=��ܚ�;k=������������8��]ۜY��a��q8�3�9z��r�:9����r�u�T�!n�c\�q�'����~���u�G�����u� �d�u^��a�i�%�)��k3����>�{��F
�Clh��f�v����N��wǳ��:�m�Z�FWOl�r���w{�w�K��F��������_�| >�38���32�j��\�m�Vk�m�rJ�JiU�tMm����.s��$�U3�����~��>q��$�&�m�+���%0S&#����$[w&���:�<Z�(���+I��{��.q��DfZ��TL�*�4��z�B�����ovJ�m��}���6�"���m���R�m ���	Ӫ�q��$�&�m�(�����H��&�����<I/y�-Q�4�j��|��aN|��n;d�v0�i��l���)鹹s���{��؄�֬��&l� w�y�x�E�rjI*���Ē���RI.�౉U��5#��$[w&��% ȉ#��4�	���`&�)b��9�8+��)�f�с�0����N0��J��J���EtĐH�j�]�7h��T�P�T?<�-�w���[o~ɯ�7m�>���=	/BIUS��M)MII�
�j�iU�����y��̒��oa(S3����l��Um���u�<r�*�&d���q��"��zM�����s��fe��ިJ&v�6y����rJ�SJ��4���$���3�H��MI%_u~x�W믹� ��P�R���#V�Y��+�����F'�.PCc=���ځq�e��ww��ۛM�*LSP�i}�m��j���O{��6�^:¼�B^Q
�M�g���6ߤF��NB�Q34���V�o'���5%		US��m����8�gs-U����-`H��2&�~x�UU)6�o�}�r��(�(�? ��`"1 *F*)����H �  ` �H�,����l����w�s���ӗ�(�%�D�抶��IG�I$�D$D+����.q��~�j���O{��6�6B�(	����4�m�yH��
�.h˭f�r�g���[m�z�^��{����m����.q��VV�9�)7:��^�ֶm���n;|=^sgS�z��Y]�1�����θ�i�������󍷏e;m��fqlBP�G{M����m��ůS��U&L�SU<�m��*�%�e���8�fnګm���������ܩ�~��r�WWh��_�����l�e���I%3;9�<�m�뭧m���q���!��9�\�oa%��V��Qm��;��q��q�S��(Q��W���{��s���	���5�D�Ңf���y=�O8�~��	G�Ϟ��I/����y�I.�a�$��چ�q�8K�\�P�q�chKu�ݓ#��#�{����t�N-n�s#[f��Ȕ�~ }~��v�o>���m�2�Ԓ�L��s6y��>ˊ&����$�Iȵ$���3�>�����v��{9�<�m�㬧z�%2�W�Ć,��$x�Ƥs<�$��톤����<I*�-I%}���Ē��)MII�
�jjj�m�DG�BU^��O8�~�:�;m���8��ޤ�L��(��o�������O\et�����_c�Ԣٛ����y�t[m�O{��6ؒ���_��D�p8�H �	 �cv�   őI�].t��Ms��n��wj���ێs����.��wOG,[W�[֗[[8mv��S��m�:v=��c�һ���^����e�����b�ܕn���j�U���n�T��<��ch;C�V2,g���8���m�X�H�P��'F���P��gM˲�c�5y�5��u�A	���Χ�(#�jkMz�˔�q�<ܜ��/LGQ���յ�9���m���\�m��]�o������/�J���?�~,O~n&������Vw2��(^JDB�:�}6�μXw]����qba&F����h.뛒{��_M��S��AX
D��j���j���߭X_)Y��
jJUJ��k7'@?Q`!�G;����'��훒}��lܝE�b@E)�n�lV'�.[�*�m���,wGL�0=}�06��0	��e����ul޹�]a](]7Z]urg:�%���$�f����u�����s��F�%*�NiMS�_��Z�8�ܛ�Xj^$" �@����Ձ��^�R����$�TҰ8�ܛK�Q�
&IY����fZ�;��W�$���� I
�����O��U&L�SU7$�����'=�훟�(B+V**��߭X���`Y�
�4��R)�E54X�rՁ��Z�8�ܛy""�R(�b�������^��?�@恊�9��`w���BK�BDDH������I>?~��;���{��q�4�jd0Y �?���vD�˨y4�u=W��:v�ŏ�N7q�5�I���6����^��[)�y�w?�?	bAR�! !��j���+ޗ5HSSL�TK������o�T�E�R �@"���DDU�~�`{߿Z�8�ܛ �=�SL�ȢI���4;��m�76
��(� � *�A@)�@? @E�"! �!!(I
M���l�x����e>ɣZ�5��˭����� ��B*1T"u�����`c��M��c�,w�j��b˚M8�E �&��������Q	y(D%	R(�T")R(@>�����Z�33-X��4�r�M�lr]�.ܯ\�tc�;�6�X�c�˘.˸��2̙� '�"� #
@�9vs.kV�fd�j��o�ο;ܵ`ffZ�8�ܛ ��xU)�T��MM9���{����"? A1""0D�:�����Ձ���6َ���D/З�P�	
B(EX$������n��.h����V�߿Z�8�ܛ��XX�rՁ�#��i�UP�f�K�V�H���� "���ٹ'߿]~��s�~ٹ?��$$��@�O�"$!"߿_���W���
ji���uR��/ ��tt��GL_tL�,?�}�2�n���[s�"�ܥ03\�Z��S<��W�Q7����{w{���?�N�sD�揀��X���>�'W��}!�����#^���N���T���W�""l��l��u����-^���	L��/\�H�$�TҰ:�~�&�y����:`�.eiȒ��6��z~��|��@�߷4��V�Nf̀b�zU)�T��N�,�����I0=}�0$���*��C�p�Q��L艪���
��$�����$m�e  �` ��l��[���Ê�Z,�S��;Cb�jݨ�B[��Y.D}�� ���>F�!�a�PK��ƍ��<Ţ�ln�A
��pc;s=��9��<�sZ�4�%H��*c�c�X��M����.8��#��Z-��6�v�s�(:ͱk��b�Y�k��{ll.^&(\H\a�4�%�ǉd,���]\���4��l�����P�#a�S�1��L,��o���|q�����ng�w�nh.��nJhw]����qba$1�24�8�ܛ�
��芣��ʿ{߭X����I~_�(UF-R�~�5HSUMʪ%�M����_��̵`ffZ�>}�M�|�O��ԺtۚT�a�^ I����|�{޵`|�ܛЗ��BHI"�~���X��l��&��JuD��Ұ2H遷�IY�GL�|KX0n��.2���N �bַ�ܶx�)�ɔ��%7N�����B�����\��H�*GUSK�k��M�����9��V��hvU�Zr$�1�9�oƾ��x>(@2�q�f,�(U�i�_�@�]N~�,{}j����7�	z��"����y���UJ��3R����Z�33-Y�IB��^f́����>}��̪W5%��\��r��U ��{�+����XX~��n�X�w54�*��f�˚VϽɰ?%�B"""�
������X�e�>��}$�hHB:u��q�*��r��9�z�q��gKX��5�%�ԍv�c=Q.�l�a`s����2ג��D��	%�=�M�j��˟&�Ӧ�����̵~��DBDɻ�Z�1}���=�%4����Z�&�H8�`w����{�e�P��8P&fI��	���0��|
�5⡨@�B�xI~q�"F"��=P�@���&�4F�J2B(XBm_�u��\4RVI����(J�d�ki"�$��f�4���$	����㈆�D%��#B"
 �A�����|W�> ��>��������^!�	��xkٹ'���f��YsI�H�*G3SJ��(P�g3f���,w2Շ�D��{�`W�O4�IBbdr=�rS@���=�w4Wuz�n�)�)N"�c�{���6�ɐ�q�\����Vڣ����o����
��T���Lԩ��;�����Z�>}�O�Q��v�}�W������䒬�X]��V�e07�t���*��9��W���2k���,��L�CŔ�����07�d�07�t���35HN��&��56	z�No�<X�zՁ�s-XJQԒDg�/�\$Q�o|0u։IB$���@��b��X!K��b����۰pA����7$�=/��:R�2�4����s-X���|����=뒚z3��M��q52cpF�I�x���=FʛW`�s��gNp%�{<�{��U�M�>K��2�Q554�7޵`m�D�ޕ�`{�t��*5�u,�����VϽɿBK�
&L�*�`w��4z�� ��̭9P���������̵g�B�H�H���zՁW�= �0���I�`�x�yٖ���j����6IG��BS���_$���LR2LM9��n���rl����9��V ��a�@�U�{����[߬�,0�?�~��	 �at� �`p�<�mzv��+�Ge̙��N&Q�ܺ�ƺ��Lm��Kʺ.K��z�%p{Bu�k!۷Q�qD�gNS�y��"j�.tX�.�r����:�p<=���
u�+Z�]ڍӎ�u�XS���Ic�z5������!��2�V�.z�/2���������Me����wu���!jƄ���������/[9��q�!��ޙfd�)Azg�{��wn���v�?8d���35���k��M��qV;�k�	(�����V��� �iL�E:��>�*��D(l�7mX��VϽɽQ�d<�=�s��ɠ%Mw|遽#���&��� �]"�u4�S�&��+(���{�`u��lz䦁�u��;-ˮ,_��~#q�`q��6�(�j�8ٛj�����;��	H�Cj8�b�O�v���ϓ��|{;�7^-���\t��m�u�5ŵrHŘ�O՟����􎿟U}������r9�B"78hw]����R+6	$ ��B0�HVHA E$IB�$�U�=̵`s��v��X_�!B^�_ʣ_��L����1U'34���֬v{����5V�ٛj���q6K�T'3P�iXqo�[{�@f�W���(��nh��<�� 
8��Š}�U���{�{ߺ����V;=�`s?����g#	u��h�_<m���c���P97M�d�L�S�ʜ�n�Tch��,�:`{�K�zç��ƀ^��_5k��I��n���q�wa`s��W�ًum�6R���]�YL�~�����}�_���s@���쵕�"J��h~���~��`l��07�t��.��;�-r9�̈�ǎ��s@��fu��3�=���z䦀{��*�iB@��#^���&K+��cp]��\8�g�n[P#�1�y`�Nco&'&&����V;=�`}���K�>��V1�Ć�����G3@�U�{nJh��V{�j��l�b��2�u.���'��}��@�빠w[��y]�@�|��h���N]0�4XjI'���`fnڰ9���.hIY �����:���v�㑼$$��w���J>��|����;�� �w��1���]���λ
��c��n]^sgUy��<�^}��Sn�f�q{NYLE%�6J�0;�:�_z�Oߝ0�/���"J��hے�wrՁ��Z�;�V��!��MT�uJ�/�,T�`O���t��� ��*S@������#$ƛ���+~��`l����Y�GL���P�t��i2�����a`owU��;����w4��kPO$�I2I$�$��H �	 t� � B�u���.>!h6Á3�8���6_�ގr]�h�^L�λ����t�fH��G�#�N݌��h�b�]L۩���h^�˷g�-	�\v��S<1��ݧ>���猄���4���i2��4�86 �j嵴���an��v���]�q��u!./N�:Sd�bz�-ϻ��e&r0�^�ڐ�q�chO]�M�Fd�<�[\�س㡺�NZݸ�R��MH4����>4{���n���=�O���u�%��,p�=�:`{�A��VA�n�.�pq��L�;���<�)�{nJh�]��ܺ�X�1��bn9�C�6��;��K��-X~P�I�n�X}��|ӑ%	�m��hے��[�������YMަ�J%Eƺu�:�QÞҊn�w#[�6\����	�P^�'��C�b�#���x�{�w4�2Ձ��a�a��ZX�=�
��Ia�s4nI�}�~!b� �D��K�,���`w:���-_�1U�$�6�"9����{nJY�Dzg7}j����X]R��f���K0V�`l��`ott���ߗ����/��P��E�������GLt�0'J�0	�\.����nu�7����a]n.��.����<;�kNwf"�߽���c�|���Y5]�����d�d�0$��M�D�#���`s�X^�ٹ���:߷4��h\��ӑ%	�m�j�;���>�rՓ
�$��\��ۚ�ύ �ak��#��O4$t��L�������R��cM��:۹�}���~<��O��빠\��mƠӉ���:�s�ַ<"3��sX��u�	0����#���AI�	2Cs#Nf��YM�U���{��8�7vՁ��+u˪�Yif
���$t��J��;S�b���%L�CSE��ͺ`t���2��vQt����rD�uJ���)�{�+���`w1VIqBP(P�8�B��_���;�4�R:��&GUSJ���XX^Q��珀��������u58�P�b������td^�r���۫E�Vq��>KV���ɜ��#diȒ��6��4m�M�z:`wH����E��3+_Úr��ﻖ�T6fnڰ>�֖يS@�ث�)H�1��h��h�+57��ZX�m������UBs4���a脓��zX�U����w4�w43�yjj@I�r8Xf*���IB�sx�f��ead�_C4���lڱOtc¢D*' �q�#T�RIFA��a(V4�4�6�*�J�* _7��T�s V�ά�     �         �   m         �          p   	�     �     V�         s[`�[tH��ӵ�Ú���3�Jyե��r�L�1p��t��nn�<!���V
 %N��x��a�H�A��j��\xvT��s!Ut��)r�UU穭i�._l%��<۞�8D���l�Ě4�ܕ�!�lF�-PWn^�i�p3XN�,\���ik/\�B�[v��9O`���F)ÛC�w8v-���6�uU㍡��`v�C�5-��6A�����;-��w/nys��w]@f�;s�{��ܧQ��8�R@�:;��Z����r������Ţc�-r�9�S}����nއu������W�:	'L,��Y� �c\��p/d[�(�f&52��L9�GTĳke�\N�F��ś:^�8yg<�v��Q˓۷m�v�s=���7n÷m��ѳ���˹S�+�����q��uu瓵wd�s�ôϵ�Ͷ�;j���^�j�Ht[�;����3�r/Z*M����5�9�S����Eۂ�ե��[]N9m��5]���Eu��m�W[��Y&觍��J���V�vFG'2l���nÚ#m��	S:m��m�ޅ���e8��fR���
�R��t��I�^ݻ<���QF;IV�׊s�]�agt�WIAE�j��1v�h���ݡ�e���P.���vV����$�e�c=�9����-`V��8۞9�`p��-�<����� V9X\u��ƙOj�8���\�+Z�ee`�7\���4�ъm��.�Չmb�Ь��inr�ʖ�]D�$�$��]$��ȶy�S���Qq;�R��Fz��&�����|�TU�(����!�8 �����g���� �m �	 �cm��`  <FrHvN��t�vmga�Sڛ&��nĵ�˕�:�,��m�\Qd����j֥ɞ-����m�{wWQ�s n�G/�:l�Lu�ݲ��m� n��.{,q)�W'�,�f3�����7c\��ۉ�hÂ��N����gs8�/[�ݞջt�Ft�	i���M���;:t}�Kj�����K��=�!�lg^L�G2��Yhͤ��d�#�3o=F7\Dg�;����쎘�:`{fA��a-�n�.�tqȘH5��w[��y��=����Z���=�z�q.��.�M+��-��a-�����GL�t�%�Sn�L��j��zC��,�k�t���%��,H���aE��K�GL�0=�K`l�����]��LYJ�&�-�1v��]���[].!A������hYL�o�E������cM��~�s@�@�ܔ�=�w4
�\2c�����h��뺘*2$�$"B$�"J)E
Bc0aD���VH`�bŋ �H	bŀ�1!  F$X�E""���p�H$F#dU�"&<�}����0;�t���U�����	H6��=�%4z��>į�}��u|�{��qE�N�n��#���&A�ml��u^,�%˪V{�j��̭��;�ZX[w4�qS�Č�cQLCajC�����Z-�,��Ȏ�3:*]�:�)�<�:�e�LҰ;��vs+I��7x��"X�%�����"X�%�O�vM&j�rRd̓UN�p��L��]ݾͧ!� #�2%�����iȖ%�bw���6��bX�'��{v��bX���Dn�L�T�J���&Bd'�w�6��bX�'��xm9��P<�Q�(B E!
h� OA�yQ;���r%�bX����m9ı,O��۝�sRkF�h�sFӑ,K? �ȝ����ӑ,K����~�ND�,K��}�ND�,[��ND�,K���&I����f�˚6��bX�'��{v��bX�'���6��bX�'�w�6��bX�'��xm9ı)�(��[�N��N]9U"�'�/o"�Ⱦ^�yT㳩�ԃi嚼��%mnf3Z�3W��Kı;���M�"X�%�����"X�%��{��,K����nӑ,K����i,:k.�������Kı>����?)��,N����ӑ,K����~�ND�,K��}�ND,Kľ���%;��k2k&5�iȖ%�b}���ӑ,K����nӑ,K����fӑ,K�����ӑ,K��{�f�Y�f��u��ND�,����nӑ,K����fӑ,K�����ӑ,K�v���Mw���r%�HL���6M&j�sLd̓UN�p��V%��{�ͧ"X�%�����"X�%��{�ND�,K�뽻ND��7���{�{���`
��uხױ���q�(K��F�6}
&��,5�����|��%U*�p9�3E����L��[����Kı>�{�iȖ%�b{�w�iȖ%�b}��iȖ%�b}�Y��WTT7H�4�L��L����p� �,K�뽻ND�,K��}�ND�,K߻�ND�,K�>���Tڙ�2���	��	�����"X�%��{�ͧ"X�%�����"X�%��{�ND�,K��G{e��r�iә�w�&BbI��v���Kı=����Kı>�{�iȖ%�b{��۴�Kı=}5�K�ˬ�.�35v��bX�'�w�6��bX�'��xm9ı,O~�{v��bX�'��{v��bX�$��w~}������ H@8h ;m�@6ؖP ���o�:�9�gK�����v#!��ݦKWi\r�F$:��t���qb�e��-t
]\t�NOcN���K�YR�<�8�T�<<m6Ɍ�ݪ�0tj�7l����.%��8�j�ۆ�����a���B`���֮Iu�[mq�z�U9�n���:� =Q�e��˪tT\9�����z� ��(��[2�3Y�5r�яX2�)� ����������q��r�Nvd�s��4=�g�t��w�w�{��7������m9ı,O~�{v��bX�'���6�șı>���6��bX�+���4��j
�e�L���	��	����ݧ"X�%��{�ͧ"X�%�����"X�%��{�m9ı,F�wd�L�T�3$�S�\!2!2���m9ı,O~�xm9Ƌ��wj�B]��w�B]���̷+.K�M�$�O~�xm9ı,O���iȖ%�b}��۴�K���"w��~�ND�,K�v���-ֵ֤-u�-�ND�,K����r%�bX�}���9ı,O����9ı,O{���r%�bX�t읹̶Ս	=[sѡ: Wu�mv� ���pg��,.�خP^�;��s�I�r�������bX�����9ı,O����9ı,O~�xm9ı,O��y��K��{��������\�+=ߛ�o%��u�ݧ!�>�P���Ȗ&��8m9ı,O��xm9ı,O��{v��bX�'Ϧ�Ia�Yu�e�&f�ӑ,K�����"X�%�����"X�%����nӑ,K����fӑ,Kľ��eô�a�̚ɖf�m9ı,O��xm9ı,O���6��bX�'��{v��bX�'��xm9ı,N���h��4�3Yuu�6��bX�'�w}�ND�,K�뽻ND�,K���6��bX�'�w�6��bX�'�O����WmY'drv�y:=o6�n}�}�7ǳ��u�ڨ�v�l�r����m1��Z��w�x�,K�����ND�,K߻�ND�,K��ND�,K߻�ͧ"�	��	���i�ҙ(C�ni�.	bX�'�w�6�����,N���ND�,K���ӑ,K����n��!2!vz��rꂪ��KsJ��Kı>����Kı=����r%��|�GA�,`���R�/��,���c	�"%�V���(Ak��PȎW��᨞��߷iȖ%�by�{�iȖ%�bw!��Q!*����RLҸ\!2<%$,���ӑ,K����~�ND�,K�{�ND�,�2'{���ӑ,K��j�%�6�uH���i\.�	���뽻ND�,K�{�ND�,K��ND�,K�~��"X�%�����v?	��%�O&���_&�ӑ��p�q�5�M�BdЖ,�7*s[��;���e.f�ӑ,K�����ӑ,K�����ӑ,K��߻�a�	�L�HL���y�.�	��	�o��<M)S�ɬ�fkFӑ,K�����Ӑ��"dK���ӑ,K����~�ND�,K�{�ND�,K��y�!d�3L̺��ND�,K�~��"X�%��u�ݧ"X�%��w�ӑ,K�����ӑ,KħO����Ԛ�YffI��iȖ%�b{�w�iȖ%�by����Kı>����K���,���w�iȖ%�bS��w�K��3U�5nj�9ı,O=��6��bX�'�w�6��bX�'���ND�,K�뽻ND�,K��{��!jH�5��nɒ۲�ր-��[a�na���u�ݗ�v �+Edu�.f��"X�%�����"X�%��w�ӑ,K����a�Q'�$��L���q\.�	���a��tkZ˓4Y��iȖ%�by����?r&D�>���M�"X�%�����iȖ%�b{�{�iȖ%�bx|k�l���3H�S4�L��L����pr%�bX�{��6��bX�'���6��bX�'���ND�,K���j�ɩ��UMQp�Bd&Bd/����Ȗ%�b{�{�iȖ%�by����Kı=����r%�bX����ŭM)SS%I,���p��L��]���"X�%����xm<�bX�'�~���Kı<���m9ı,OO�쟍�0�g�[@ �@ .� Z������N�{f6��9ɨ۳�.�ϐ���ι�V�N�vd�r��պ�����t�ݠ�����mw3�C�)�t��u��f��[�-ZWk%�`ͩ���6K�i�ιt]�v^u��<���2���m�.=clb���(z+�a�j)v	nHp�$���������ir͕֘ޞ�:�ey�����a۞k�BΚ�g8	��ϳjmP��j��Mߞ����oq�{�{�iȖ%�b{�wٴ�Kı<���m9ı,O}�xm9ı,SZ�d�L�T�3!3J�p��L�����i�~�DȖ'�w�ӑ,K���߸m9ı,O=��6��b2!>��٩SUJf�j�h�\!2�by����r%�bX�{���r%�bX�{�xm9ı,O}�}�ND�	��=�t�uD��R樸\!2��'���6��bX�'���ND�,K�~�fӑ,K��߷ٴ�Kı;��{�jL5�eɚnf��"X�%��w�ӑ,K��߷ٴ�Kı<���m9ı,O=�xm9Ǎ�7�����e�%׆83d��5�/`N�֌�ny�{]�w+��5���ws�[�T�&�Nf���p�Bd&Bd.�/fӑ,K��߷ٴ�Kı<����Kı<����r%�bX�Jֆh2jd��ST\.�	������r:�� ��T۸��bg�w�ӑ,K�����ӑ,K��߷ٴ�TlKľw.�4au�5�.�jm9ı,O=�xm9ı,O>��6��bX�'���ͧ"X�%��̽.L��L����	�����Z�ND�,��"{����r%�bX�}���ND�,KϾ�fӑ,K�����ӑ,KħN�'d�4fj��Y34m9ı,O}�}�ND�,KϾ�fӑ,K�����ӑ,FBd/�7��p��L��]�ӎi�tU$\\][�7:��EM��nZ-�;v��3�:���zI�3�{��N��n���.6O�r%�bX�}��6��bX�'���6��bX�'�}�ͧ"X�%��o�j�	��	��+�4S�	R���ӑ,K�����ӑ,K���ٴ�Kı=���m9ı,O>�}�ND,K��Oe�I�0ֵ��i��6��bX�'�}�ͧ"X�%��o�iȖ4]� ���)�D�oYsX@鸐���GI#!b��!���(d`���M�xbABIAG<�a�r�i�RHT2MSRZ$H4A��BV��K�sZ��XF!�Z1�t��֓��W2S2\�spt1"�(U��� D���M��DP���b���!�H� A0]�Md�i\�`|��R"i���"{� >0F
����>}Sbʏ���t�'�3��ɴ�Kı<����r%�bX���ۗZ���73V�6��bX�'���ͧ"X�%���o�iȖ%�by�{�iȖ%�b�̽.L��L��uV�3A�S%V�jm9ı,O>�}�ND�,K�{�ND�,KϾ�fӑ,K�w�z\.�	��	��n��2f�E]�����sc�d!t��%G]��s��m�1D�̉���M.��=ߛ�oq��O=�xm9ı,O>�}�ND�,K�~�fӑ,K����iȖ%�H[�nP�m *	����p�Bd&Bq<���m9�$r&D�>���6��bX�'���ND�,K�{�ND�!2Z�dЙ�3LNe���&%�b{����r%�bX�}�xm9��,O=�xm9ı,O>�}�ND�!2]��4Lҙ(�L�p�Bq,KϾ��"X�%����"X�%���o�iȖ%�� ��4UM��7�.L��L��V�.h�T�Y���ND�,K�{�ND�,KϾ�fӑ,K��߷ٴ�Kı<����r%�bX�:k��35�S�v^��u��c�(qa|�gLFz�[H�9M�6Y�\k�����7|�~oq�X�'�}�ͧ"X�%��o�iȖ%�by����Kı<����Kı<=5ӷ5����73V�6��bX�'���ͧ"X�%���w�ӑ,K�����ӑ,K���ٴ�K�L��uV�3A�S4�UUQp�Bd%���w�ӑ,K�����ӑ,|)!I����p��L��Y�~.L��L��Y��f�[u,���R�\!X�by�{�iȖ%�by����r%�bX����6��bX�'�}�NE2!2�[�&H
�dn�i\.X�%���o�iȖ%�a���y�m<�bX�'���ND�,K�{�ND�,K� �@�!��{�����~?_��D���   $m��`   yIMםI����Ν�mmӷ���G���]�n�nn�z槄�ݎI:.�*n�K�_Y'�/m���b0�^ulKȞ�\s�8�q�����pK�9P�dtْ]p��Nݞ\v�	�$ۧ��l�v�8ᱴݶ�1��f���%ӡ+i��s�����浜ׅ��cl�8��������g��0���#����]�;u�Y�m�����;�Ǐ-=���&s_�����;��t�19�T\,!2!2�ޗ�&%�by����Kı<�����3șı=�w�m9ı,J}�OzF��S%���.L��L��f�m9ı,O=�xm9ı,O>�}�ND�,K�~�fӑ�,K�k뙚tꔌ�U34�L��L��{�ND�,KϾ�fӑ,K��߷ٴ�Kı<����r%�bX�ã�T�*��ʚ�SJ�p��L��_fo�iȖ%�by����r%�bX�}��6��bX�'�}�ND�,K��];sY�l�ә�˚��r%�bX�}��6��bX�'�}�ͧ"X�%���w�ӑ,K���ٴ�Kı���C蟰�X���u/q�f��e-�JtS+�p9�n�zFr��ٓ�qzYΰ��֮�6��bX�'�}�ͧ"X�%���w�ӑ,K���ٰ�	Cșı=�w�m9ı,ON���G驖�K*d�4\.�	�����\��H�OG�q5������r%�bX����6��bX�'�}�ͧ"2!2qe�C�A27U4�V%�by����r%�bX�}��6��`	bX�}��6��bX�'�}�N�	��	�[�hLҙ�2fBj��Ȗ%�by����r%�bX�}��6��bX�'�}�ND�,KϾ�fӄ&Bd&Bk�#vF��S%�u4\.D�,KϾ��"X�%��
{����yı,O{���ND�,KϾ�.L��L��h3X�S�\ӗT&j�W<��'.�:�����R.a��]K��1,Fr�+\�WJ��������o}�xm9ı,O>�}�ND�,KϾ�f��3șı=�p�r%�bX�d>��I��5�]7Y�iȖ%�by����r�dL�b{����r%�bX����m9ı,O>��6��bX�'���v�Rٙ�35�5���Kı<���m9ı,O>��6��c�4�MD��w�ӑ,K����e��	��	��.�ֆh'T�MS�6��bX�'�}�ND�,KϾ��"X�%���o�iȖ%�by���\!2!2�6ܴ=��mԲ�JuFӑ,K����iȖ%�by����r%�bX�}��6��bX�'�}�+��!2!{(��>sM���t�2]c��JnǊ��In�5���țc&t�I�3���)9r�H
�dn�i}�&Bd&B�߷�6��bX�'�}�ͧ"X�%���w�ӑ,K����iȖ%�bU�vM	�S4��XMQp�Bd&Bd/��}�ND�,KϾ��"X�%���w�ӑ,K���ٴ�Kı*�ݑ�j���̺�.L��L���fӑ,K����iȖ%�b{����r%�bX�}��6��bX�&�����ӧI���M;��!3�P�D�����Kı>���6��bX�'�}�ͧ"X������"sș���m9ı,N��_���M]fM�j�9ı,O}���r%�bX�}��6��bX�'��}�ND�L��_ef���!2!}���N�э	�^�^#�^�u����V�S�Φ©-�k�f���3`�ed[��{��7����o�iȖ%�by�wٴ�Kı>�~�l?<��,K���ND�)	��,U����S�Tꋅ�!8�'���6��bX�'���ͧ"X�%��w�ND�,K���ͧ"AmP��4hz���	��b�
>��ĐI�{��p� B�������Kı=���m9ı,O~>ݔ4m �"�t�nL��L��sy��Kı<����r%�bX�{�xm9ı,O�߻�ND�,K�>�4�J�2�f�L��L����pr%�bX�{�xm9ı,O�߻�ND�,K�~�6��bX�$2�P�!P�!mE���i�V0��#ӽ��[sZִ$ m m�H���m�N#��.^�9����b��ͥ̒�ɯ'P�^�c�s�p�yx�rb�n+�5�v��Y�{5�睃	�s,J���1ki��1�nuۅ�O[ey۵ʹt�3�A��e6���t���=vût�g�|3�3��Bې�5�';����P�n��Lg6���	�L�!.0Қn�ۯ_�����(b(F�%/��^�M�������7>ļq���N�j7jt�6]l)6�{���oq��O=��6��bX�'���ͧ"X�%��w�ӑ,K��o�iȖ%�d-YXh�j����LҸ\!2!8�g�w6��bX�'���ND�,K���ͧ"X�%��w�ӑ?T�	��L���h��'.�nL�ı=���m9ı,O;��6��c��DȞ����ND�,K��fӑ,S!2�jٚ�*��f��Ҹ\!1,��Ȟ��?M�"X�%������Kı>�~�m9ı,O=��6��	���i�UJ�:uN��9ı,O=�ݻND�,K����ӑ,K��߻�iȖ%�by߷ٷ�7���{���}����L����c=�9#���i��Bt���r���d�s��Tt$�9��K�ʙT�L��L�����r%�bX�{�xm9ı,O;��6��bX�'���ݧ"X�%����r�H)��9����!2!}��NC@���|4�'"X����m9ı,O~�{v��bX�'���ͧL��L�֬�4&iL��3!3J�r%�bX�w��m9ı,O=�{v��bX�'���ͧ"X�%��w�ӄ&Bd&B}��T�SD�@�]M"X�%����iȖ%�b}����r%�bX�{�xm9ı,O;��6��	��r�����*�dL�U;��,K��=����Kı<����r%�bX�w��m9ı,O=�ݻ{�{��7�����~��R���6��#;qk�M�%]��RLs�6`�e�H���&�&�4M۠���M��	��	���oӑ,K��o�iȖ%�by���r%�bX�g�w6��bX�'�ƺ�f��ʪ&\�:�W�&Bd&B�r�m9ı,O=�ݻND�,K����ӑ,K��߻�iȟ�*dK!jX���UT�ES�.L��LO~�]�"X�%��{�siȖ>�Th@� @:4n&�}���iȖ%�b{��iȖ)���nZ6h�r�s!5N�p�ı,O�߻�ND�,K�~��"X�%��~�fӑ,K���}۴�K!2!w[�kf�)��9�����bX�{�xm9ı,O;��6��bX�'���ݧ"X�%��{�siȔ��L���O}#uNi�.��M�IC�v��7[sP[�e��=�z��*Y77-v��V��u��̚ne�3GȖ%�b{���6��bX�'���ݧ"X�%��{�siȖ%�by����Kı)�a;ܚ���2P6UQp�Bd&Bd/�Y��p^B9"X�ϻ�6��bX�'�w��"X�%��~�fӑ,K����JN��ԕAIL�U;��!2!d�6nD�,K�~��"X�%��~�fӑ,K���}۴�Kı=�v��J&�m�Rr��p��L��_w7���Kı<����r%�bX�{��v��bX��O���ͧ"X�%��~���Vl��D��������ow��}�ND�,K������yı,N����ND�,K�~��"X�%��������L�a.�w&u�:�Ѷ��5�'X7`LR��=	�BX�<ܩ�o\'a�j�˫�]jm9ı,O=�ݻND�,K����ӑ,K��߻�iȖ%�d/�/K��!2!|�m�F�.]]e�&kWiȖ%�b}����r%�bX�{�xm9ı,O;��6��bY	���f���!2!w[�{.���3%��k6��bX�'���ND�,K���ͧ"X�%����iȖ%�b}����r%�bX���rvL��M̲f�6��bX�'��}�ND�,K�u�nӑ,K��=����Kı<���m9ı,J{�N�&���Y�R[3Z�ND�,K�u�ݧ"X�%��{�siȖ%�b{����r%�bX�w��m9ı,M�GdӵD��M�:`b�)6HJ�a�ى*S���a W�s�.(;�"��4�U�ۊ�}%`IX���RnT�b�7�h���uh���\#%0�	

� �"�ГrV��9
:���`jB�D�D����@ ��ؐ`A���[D�^sd�f��� `�@������@TW@h�7*�¬�M�ؑ��͉�f#��9.`B�.�͊�jc��$i����1$�Z���O�G�S�Z	��ZA�]     h    �   �   m�        m	          8   ��     6�     ��         �Z
�e�bB��Gc�	zu��:9���/U��\�4�qN���N��ѥKX���7lgm"�V]9N�6�"]5�+�α:]�\����M剎�z��۱�]FN�`:�������I���`�\Wj@�e��W�my�ج�gm��c��R�M�z��k�nϞ}��[z�\a��q&(��X����r�7l�vv��y�۴tNUٹ�wb�HQYb;#- �Mqe&]�Nv��`�����؛<�#&lvU�:z�;-�Nzݶ�ݍ�h��2�9�ݷ�;Q�A%.ͱ��݇����[*��Z�gv��IX�R�ٜ5C�e�eN��R������&#Y�Ump=�sLi80���ًK�;0���ra9.Sq�vv�ç�s���Gl�(��v��J�b��v�.]c������hzi�ö�e�<�pI��'l@��,�gkZ�(林�]J).+j�8c5k�����9-��-�'S��#���p�h�nm���6J%��]<Ge1�z�T���m�O��d�[T�N�d�����q����FG�/mY���8C��^ܧ
�>�n��_g�YJ��v��8��ֺeM�9�PK�F�tU�m���*��i҂�R ��a�j1vs��W@ :�/OO �s��&������9�GV4X�qʜm�z�HTc"љ��Nћ�܁�H�$p�8-Tsj1��1Prx6���j��i��Lv��j�x� *�jg��-��ܚ��q���q�Z}�7:\���mճl䲁��ԃt�;\ݛ7j^*��A�)�u�����{������|C�OC�=6�"��w������{�?�?^`$a�m ��� ���	<'GdLѹ�b��mc�;I����w\�;:㗢:.:��y�]]N�Ƹ�b�\k��lm��Ɓ���iuq�wZv�lunӦՀ�ܑ�A=�1=\�k�ѓ=2Y�r����j��ĝ��׈�N���I����zz��1�X6��jG`k�����n����MvL�ﻻ���w��3�>��!"฽]��G&N ^ݣ�WV��sێ�m�V��띻/L��s,έ�L~����oq���}}�siȖ%�b{����r%�bX�w��m9ı,O=�{v��bX�'�-y��M�T�9uSp�Bd&Bd.���m9ı,O;��6��bX�'�뽻ND�,K����ӑ,K���[��U�TI3T樸\!2!2��}�ND�,K�u�ݧ"X�%��{�siȖ%�b{����r%�bX�GUkC���J�4U:��p��L��_{���9ı,O�߻�ND�,K�~�fӑ,K��o�iȖ%�bx�m�C�u.]:�,&i�.�	������ӑ,K��߷ٴ�Kı<����r%�bX�{���9ı,O�w{����ߧ�e��b�j#�/�<6��[s�rs����<� ��&-U�P�Y�)��9��B���L��Y�~.LK��o�iȖ%�by�۰����&D�,N����ND�,K���I����)2fBj���!2!}�{6���:����H�M��Ȗ'��;v��bX�'���ͧ"X�#!w�z\.�	��	���u)Ԫ���fkSiȖ%�by�۴�Kı>�~�m9ı,O}�}�ND�,S!}�z\.�	��r�����U��ֳWiȖ%�b}����r%�bX����6��bX�'��}�ND�,�"�"{��~�ND�,K����a4SmJ���M��	��	��ܽ."X�%��~�fӑ,K���w�iȖ%�b}����r%�bX��~��1���]x�1͙�G���ְ8qv��"�󋎻Jc7�S]:�t�M��{b�m9ı,O;��6��bX�'�뽻ND�,K����ӑ,K�����p��L��YU�vFU*���:�iȖ%�b{�۴�Kı>Ͼ�m9ı,O}��6��bX�'���6��bX�'����K�]e˫��I����Kı>Ͼ�m9ı,O}��6��c�C �ApȚ�����6��bX�'�����Kı=��w%��ѓV2]]kY��K�� �2'����iȖ%�b{���M�"X�%�����iȖ%��&D��ٴ�K�L�֬��	�D�P�Z�T\.�	�by��iȖ%�by����r%�bX�g�w6��bX�'�k�ݧ"X�{�������B��q���������zhݴ�۴���8��� ��-Wkv��'��&$9���"�-�~z��Z��h��X��H1�Z_{�~��M�d������g��ܫ�	�Ǔ�=�}V�岚}�3�^�~ZV��s��7$$�cpNE�w�S@�U�z�W��pA�u���wrN>�%ϲ]]�������6����� �'5���iʉH�CqO�d���zݑ�`#���W"��x��]{N���:He+'b�ѻ1%yx�����{"`z.��ݙz���tLJ�1�6(��@�vA��2���{"`ձe	V$�^`�ݙj��{#�=�)��0��x��ٓjC@�R[odL��`n����\J�D�3�E�x���ޔ�=��Zz�Z�r�i�$�L�I&@p  � ]6 �� �j�����o�m�K@����I��7ǣ���U�qm;q�c]R�:�[VVt��}���z6�:�lS
e�s���r���b6��{7&[�f
q>��s#�3����<���ƶ�������;7BU��cn��r]�Ӧ�:^qV9fkvt�)6%�:�>�{��}����6�>Y,�%��u��ío<;��/�g\�Am#Q\mZ�2��$	�xLMH�����ﯪ�;�j�<^��2�[�	F��^f����K`z�D������CfGT�C��ӥI�j�i���v�dL��`n����NĮ�ᘐ�ĕլ�`z�D�����l?]���@����K��2,7��ސ`n����R[ײ&��v��ݨ�.�vz��wgn�g���PSs0/��n�θ���\曎Ml��
rV���j�l�%�={"`l��V��S�U2*Nf���ߧ1�%��B�(! �`A��lWga��1g�B0�b2P�RIb���j�T�0!��4b G1 BRF)A	 A!`�#��8�b�&�Db�"F,�8�Y���s��<��;������@���\�"B#�H�?�&��;��������� �U�P$"m☚��������@���@�{k�<ˎѹ �S��y���]-�����dL�0>���>�C�	9�YW�F ��N�N��i��d�"3�ԑ4r���=��.iUΗ
Ĳ��K`{fA��#���l�ѵ�Q���X9���h����7����]����e#.�Ie��`oH遺�[.�_}U���T��� �QQw��}�ܓ�-X5��5I̕e�3J�b!��~��~��GLI0
�Q"#ġ2cQŠw>�@��w4-�����@�aj�8��5 �9���v�r=p;�뛫khV����G<�L�r��8�Y�e�%����0=$t��]�bQ	q�d��ݚrE9�N�*iX��W�R�	L����9���d��pܐJ)�M@Rf�ﯾv{=�f�wvՁ��ڰ;)9�S&
�@�}V���h[w4=6 �u�}����x}�)o�5�Yy���`{dt����ut�s�
�ru8��,j)�l�Ƥ1Om�s\����rXy!le܅�ftY'��u���	f2,hn(�x�}��ﯪ�;�S@����R�2�#>���,���l��0=�:`zH�V)b�xbEeZY�l��0=�:`zH遺�[ڸ.�K#0�>K/0`{dt����ں[�t����e�����b#��ym��<��Zs�=빠o��jE�I�I$�$�m �	 �cv��  �bI#&�m��p�z+@;����;Lb�;˗����k=f�=T¹��-r��Gq�)����
qr�S����{�Vb�`-�ܨ�ݮ��r]����A����ꋍ�듀:�I�hG��5�خ�;s,e6��Ё�����ݗ=������F�9͙�+	3��g�G{���	F4$rt1��N9���6�j'��έʧ�כ�anpa2���6)�QB,j�=���w>�@�޻�����{���QL�(A�����ގ��:`{WKʫ�W�]]���Ie����������hϬz{��+$L��7s4�0=���;�LLoGL�ږPn	�~M�M��<��Zs�=�z�h�v[�IH�Cj'Q��lۭ�Lcq��!�$�/���$����tn$�5�4dĜ�h���=빠v���]-��\J%��e�%���nI�=�f�. �,D������ZY �RԶ��"-%~u�}_mU}Uۢ��˥�$]10<]�W	�x�"9���4=}V�k���w4ܹ�R9�E��U�`������t����t����{���QL�(A��_X��J>�^��������v�(��Q��I�0�\���4Z���#l�nۀ�te����3v�H���:8�X��1x韆�d���.����<#�	D�QI�Қ����̞�M�ϻX^�	Cf5լ�MRu%C�nf��>��2{�6R����B"Wc�)�x�9@aM�aN(@#�M��!�^f����d�l%#�&c	))3@e�XC���9��f�0��)� �D��'_\����q��@|��" .&
:�Y潛�s�u��{L-�5�4dĜ�h�����0=; ������P.�K#0�>K33���d���.����*�iBA550��D3;�&N�*�Q�a78�}��v.�k�OL�qmDM�S$4/Jhz����=�zS@=˝E#��P��c������t����t�����R�wR ���-}c�<����}V�篪�.{ѵ�X��"� 
H�od���=���߾���Wș&{��R9%ME$4+��3ޗ��|���{Қ��u�H�B�mͮ�nװ���o�|���n�N�,e����fs���]��:��~m������bE�����l��W�J�*X�75T���S�D(I���i`}��-�_U�{΂�[�2B#�q�����t��t��_T�I0��7��I����_U�[�a�y�Jh�s��s��S�����H�`{{ ��R[}^����d��J�T	X��o��v� H@8h ;m�@6ؖP ���o�s���V��s�c�r	eVƮ�,lA� ��S��u6^Ø{����a�n��y��u�2F�{\����i�KjCg���`��#�1�ѱ���O�u�l�qː�.&�,\6ħCu2��gqv5r��mG��i�V�Z;F ���x�,k;-Ӱ.��5:�a��_��������E�l~9K��ɝrb�Ѷ�nZݥ��Ű�@��������r�5�p��5�#���ߞoGLE%�=���.{ѵ�X��"�!�������<�ՠy����4�:'��9&%�v�/S�Ilj�l�40=�w4V{��dd��I��篪�:H����A�褶[\�ʻ���Ife�:H����A�褶���@��*�iBD�j)�LS���g���h9�v�{�U"��s�e��e�2B#�8��zS@�V�篪�D(��ے���[�UT��u&MTܓ�g�]�RH�HF*���V���ꈩ>��;�.K�w-^�X�\�/�Q�H�LnE�{����40=�0=��ﶔ��R��f �f���(��wy%��smX��z���@��F�*�G�E�C#4oGLE%�=���:H��7N�e����u��z������zΚ�s��60�v�Ū��]�� &�������$h�_}�z�z~t��]Z�EJ�RT9�檝�ϧ��RM���%��smX��w���wM��5U@�I���`f�ܖ>�Z���Iv>�QO&��v{�������u5$�2�sRXjJ$��o����9�����n�$�>k��U"�/>2�Y��Ilj�l�40=��,�[�zə�tK�r�R��ԡֺ8�&���vs֮l���]�J����9�5��yߖ���f���[a���2:�Z�ST��f���̹/TD(M�w6Ձ��i`s��=�X��X�Ps�f��w4I�`{WK`t����]���-bʴ�iI��e4=}V���և�dH$Y��I$�A$�A,B@D@������9g�ȸG�#'��M�hz������z�h[)�{�MN&�$J&�p\�\�xs��ݱ<��Q^܉�|s��%�.;e�$�S$B� dcnH��V�oGLI�`{WK`o(���xeU���V���t����t�I5��;*�G�`��b��yl���]-��F����Һ+X�U�*2�fj�l�40=�0�I$�۷����:�s��UJZ�D�;��&�����0=���=}%k��8� $m��` l ��;U�z��N�z�dH�j��n��nܙg�]Mv�K8��2-���sv�k�ys�<�zn֠�Ϋ8v�\j$��f�p�n�����òr�kvȝ�A�ڻ�>a�Vs�g;�[��̱w8���rnw9�ڃMԽ���m�mN�h�����U�Ir5um7lp�Ͻ���rX(c,^֮�ٶ��#�C]����b�݆+�sr��@�2����,K�oOΘ� ������I���F�:�sQ4��f�岚�����I���遷[R�F*��eX����t�Iގ��!��(� ,�F6�@�ҵ�{z:`zvA��]-��J�#3̳�Yk1[���Ӳj�l�+Zea���q50�"�������T8��uf��e̖�3lu��E٧���%E�`��b��yzS@���hzV��g���z����_�q��5��'<�~��EX@���ϳ��-����Ӳ�iK�)I^f"�	e�:vElwGL��������`lS�\��k��1���5�y�w4+�9�Z^���΍�u8�	FҎ9���Z�����ށ�u��<��S��ْ&����I��k�vpt�9�s]��/��n�I:99s�n95�rdd�6Ӓ-�}V�ץk@��v}�����r�}�Hے-yu� �y�ܻ��=˥�7�@X�#����RF�;���}V���� D�$�0#"�";	����UM��K`MR$���K����F&���s4+�9�Z^���~��_�� ��Ӎ�Q�8�܋@����D����%��r���*�NoVU�ш݆�-��6�6N�\��\�d�tp̞�^�:c%M�r�!�tI�����[ں[V�%x���pq9��5�y�]�����_U�u�Z�;���'T�`�m)#���Oq��{��I7�����6Ձ�=ʋ�y22bi���>�@��컒s�~ٹ�,�"�U|�)6s]�,Xl�t�UT
����vNȭ�����[ܺ[D��CB6��x[�%�;u�U�����Rq6�)p�t�r�qls:lZ�lV��tt��]-��]/��'韕�5e�/�P#"LM9���Z����Jց�u��nujF�&�xe%�lr�l��[����t���:��XԎ%�'�ץk@��V2{��b"�Y���ܩ���u8A���Hց�u��<���<��h��˹'�=���	 q��Hb�>���͆&�Pь� �	$cI0��`�0v���Cc���؇8�2���X���mh�+��
��j�da!Ȕ��	!*�qX��HD�  �4��a+9
��C(J�	0�$c$���8` B�P�F��2H���2放"�c��k�k:�    ��A�           �`        ��         	    �[@     m�    �     H     ڦ�����8U�v��N������re���B��f�3�FS�vF��J���b�v0k����hv@49�7d�&��gW
�G6%�\���3��ճ9�\"�`�'&�]ZMX-���.����g���V��u>���Y]��ԗ��<npkUjPF'�ɬ��s�s+��@b�;\�ꗶ^����  �K`
,�d�]���Z[38于.hՋp���9ݳ��d\Z�l�G�"��2uX�.ڣM͝�����i�j���;�1��-�,WElD�۝���g�p�7e[���7a�d�	�e���2�OH�{- vZSO��7]��-X��I��=�h�P*+��v-:��-\5�歭�)�Y6tnc	���[����ʞ���,����9vu�u��"�v�*f�^��n|��ڴu�q����ry�mɶ�ZMis�$��-��h��ֺ@���`�\T�cZwG[q@>{T�y��/ld���犹["v8�ZĻ]jv�����Lm��PrjKkbrQ���OO:!.+�nݧi�nzۓ��;�ά�%A�<'�mӓ<��G�n[�<� ��,�uv�ou���.sf����`��pc��E*�R;��$�����ݬ��*�[�X*�ŉ z�Wk&�c�'!@�6��'FR�x�G�t�muFwd�:Z��r���x�ݶS7\��.��(k���t�gʏn]��sV�+���gP^+H�g-5�:4�-�K�F�8�*� �6����b�@@5J��R�O@9֯]�,�fʃj�%�m��䆟SM�:�����(�����	a�Sh �D��E ����{����Y� �8	  � ln�  �`WW	�k�/]�n7c�΃�u��Lh�m@��]և��=FOE�e۩� �;�{w5�=/X����H�vŽx�5vNzۯl�w1��p웯���O�g�������@X�ݧ���u�70�K2�v[�f�v���'�����f�מv͚4�mS�n}z}����������#�0n�+e�#�ict�'c�e�t7K��$3�9w��lX'��wϒ��ǉ��EJ8�|W~Z����Jց�w4Y�T\#��!%k3-��]-�Ӳ+`{z:`z.���q]��L��rE�u�Z�=�0=K`{WK`oR�h����*ʵ���=�0=K`{WK`t�Z�<Y�+�b��y_U�y���+Z����:�T�Q�Ƅ�fwY�ܼݸ}���Rx�2��q�k�z.��F/L�s%-Kk���o����l	;&[����t�VҗBRƤ�D�AH�zX�~����w4,��ϧ���	�Wr�ZoeԢ��4�32�����lj�l	;&[�Ώ'S�`�m)#��^�@���;���v�'�sx�k�6F����F6�M�_U�u�Z�<���yz��-�$�N!��%S�3n��<��0my��
^9ۉz��e�s;����q!�?F6�@�ҵ�y�]� ������@���L��
LF'����� ��j�l��[���Wf�Y�K���b���~����N!���3�!�AH�0P�V�D�Y��z�k컒w�w4۝Z�����D9&�篥�:vEloGL\�[J]+QI"�<��hzV�=빠x�W�y��.2��8��jd���#S8���쩈8�p�<x�l�ԍ�9�ЭbQ�"5?F�=빠x�W�y���+Z��7��9�Q���)��ں[�dV���t���s���"1����z���J����� ��"�yb��ϱ	,̶E�&����tL;�_}U�&1�+Q���~]�<��d�>ɭAI���7�y�]����~~�;��:���~�캗ɨ�"Q5J&ON�����m0�<0�nq���*�m���bzeRR(�FFc���x����<��ZWս�z�h�9U$sj@��b`{WK`t]`{z:`z�D���X��"II��@����y�]�>�K�����-�X�"���Y�0=�0=s�`{WK`t]��9�x�q���$s4��j�l��LoGL��Wuk30p�H� �� lK(l� 	:��%/#����ԓr��k��շF����W�pX.��:^1ȳč�5�f�^�N�+{��� ��ݾ6ل�Tm�0s�Ş1���J�죶��Lh콣`�@���NH��
�tzw�ג�j�L��"�ޞ�&�>�@��d;pK��f�7f.�@L��]	q��q����yƧe&�k�����1��e��|�F]��z�Z+!Z�[�l�Z��L���b��RH����h_Y��w-~��a��ٰՆΧL�UY�!%����$���t����}V���+$Ȥ�d�Hށ�v���0=���6)`z*�w2�U�1��K)���ں[b�&����sx���목��]�)78�����0=�0=}"`{������]vGa'����s�w���i�7Z�p\i�<�7*s[���qR@�3-��H��#���L�����2�y-�T��P��;�fZ�Jr.�����:�y07�K`l�%�	��S�#�#iI��Z�}}V�g����v�ݵ`|�WrF��I�1L���L���)Ill��}"`�q]��L��rE�{qڴ�">�� Ǜ�`}����e7�4�*H�..�8n�P	g+��3.��p����`��<���1o,��F�ܷ����#�_H����6R���R��Q�S#1���.�����ێՠy��ʪ�9���LI���]-����ͯ����}�U�RZ�u�x�נv{��������@�R�ll��{"`n����;����	j~X�Z�۹�}_}���~Z�U��UD�N!��F�	�H��_��ٷ��#qs�v�x�7M3��M�fToI�JH�h�������S�z�DG}��V�b͑��RuL����&��l��[�#�^��=�+��I��cNH�n>�@���ײ&��lN���Q�����SN�RQ����V>�́�Ϫп�3�ϞIV��<�+#x)��̠K)�ײ&��l��[�#������������da.�e^ítx��g�6y�9�ٳv�+�/l�#Ji�\[yT8�PjĜ~���@���=�s@��@��X۸�H�l��h�]-����dL����bWWu�f,W�]%�����ײ&��n>�@/����c�`��RG3@��ut��]-����]]��&)��)�ﯪ�=����#�^Ș�U]�%	bUk33008h8��$m�e  �l �����9D���ڻYG&W᷅�w^�p�/Rcv��nz\��lf��3Kudt2[>�ٴ����g��a�[	9dj�ݦ݄�qp!���y�غ�p��&<ݥv���#������n�·s�.0�ƺ���,�
�Z�OSC�Y@}n��E`Y͛����^g��ۧUP:�AM�nn�[��[��#HN�uy��ཱ��n�q�>��^LOn��]��b3�ק#Q��~�9��>m��:`u쉁��[ӫ,.�F*�Te�b�Ylގ�{"`z.���S�w��g�hnәC�JI)6敁�߿&��l��[������Y&E�P&$��<���=����빠r�נ{�X۬�����@�K��;z:`u쉁�[*��>ࡌ�{Z�l�^瑉\�.��i�d���b�y�i��#j&�҆:��/���2��w&�z�u-�`�����M�$�4^��f����f$z�D�����?�]�u*~Eы&)1	�)�����n>�@�z�h���y��aO$���I#�=��[���^Ș��0=��]*��'�XH�8������^��^����h���j8��DE����r�I����6^�Fl���2���y�H��L��LI9�/mz��z�U�w�w4ەWȈ��	�'�:&�]-�����dL�N�i�x�N6/đ��}V������ lG�zK��X�`�!�҆h%�x	�:�B&�(O�Bb �0�@�HF��$Hb� ��A��d�D��X� F$HA ���%><׌J(V��]j�M�R	,����^L3 � @� �ʆ�� ;�L�"�#���xi�%� F@"�!	BBLM�:	HLU�Ѳ�`D�M��A`�X�H@H$B1��LX�
F1X�H�h�pt����1v�+B�'�;,LLWX"qae��"A��6ƅ�nᄉ��QpP�`ς#���&߀W�A�z!�U=6������{޽���/D�,��$RF���ގ�{"`z.���K���6¸�Q�$�4W��<���:������i���l�$\=F�u���S����CA+�]��/;����	����b�c�<���&�z��ZJ]-�����tL�Zt�ڬ�21�$Z\}V�����9[^��}V��c���q�P!������t��&��l����T�i�2bI��9[^��}V���rwFW� �
hA� �*s����}��q���	@����W�h�9�����V^fM��D,�5�rD���$n����v���Ӭ���ʦ����nI�Gg]RQ�]����Ǣ��3T��w-Xy�:����`j�D�,�D�~1��������+���Z}��;$��1ffe0:䉁�[�)-����ŝ�c�<���&�$z��Z\v��빠r�� �3Ӭ#I�!Z��`t�%�;z:`u��t���������_��ۀ8�[@ �@ .�  �`p�h�sp�/`]ћD��L�;sJc�C�oS�o\Sp�v���;�6��;����x���p\�:���a��58ȑٯgd��Y��v;
���-�CC�.w��l ��K��@p5;:j��؏�|�K�A�l��k��ݓ�vݦ�^�˴č�k�v�Ai��{��n(�CB6��y-=�����;�]sRy\2�Sld���zY��uI{;7a"���oۚ+k�<�����Gf��v�+A�9�:��JM����&��l���oGLe�F$�LMI4+�qڴ���[l�=ˏ*Ɲ`�n�e�$�%�;z:`I�E��^�m!e�ґA��7�����m���Z��Z��4�q#$ML����g{l���M�����p�ɒ{ge�pO�\��(�`ԓ#�
1d�g�}��@�'���9��
8�;�j����d�NjL֋.f��ַ$����q�@�TL_������;�:`I��Zt���&cNH�qڴ���~��}��@��~Zu��7r'�@�,�&oGLI1��[JR[ܪ�7��ɉ'3@-�hW�h�h�]�ˏ����Q%QH>+u������>גznyȧ��k����]�/L�v��2,$�1E$�<���-�j�;޻�m�@�.<�u��ɂ�e�$�%�;z:`I�E��^�M�q�E���'�����m�߼��UW�}T�Ų���[ �� ��b�$� �٠y_U�[�1�l%
���X5�l���C�L�Y���E��R���0	$�m��w���e!�	��ٵ�>8����y���)���(*�u8��+^gH=Wm9Z��`IJK`v�t�$����=����LO"�$YZ{�s~��}��M�����hs�
��
@c&$�� �٠x�W�[�ՠw�w4ۇW$Ȱ�j��@�^�`f)�v~�Z�Ű���Q�	$�D(��r�v�-R�Թ�	�3@઩�$�%�;z:`I�\��D1��s	u�.��a�N<�a{$v8����;=[b��%���Шaӹ����2��0	:c�:&��[ ��l�b��I3@-�4��q�Z{�s@�gqX�)0rbrI&��^�n>�@�_U��� �x�[�U%C�]UT�jP��U����lN���Ή����JVU��0�d�h��޳@�^�@�U�y�������d�I2I#�[@ @6�ݶ    x�Lݱ�moMu���}�9�=�c��\a]×of��E�,�Fۆ�n4�λO���-�\ח=���Ж§��&�lv�)y빶r#b�m0��6��.�J�U (n�kvfCt
�i9ó��i.\u�&3e{in�����p��6롳���١��p]5a3G�Ν����:C�HZ� �����#�y��{FgW���8ݹ֊�e�����P;��1(����x�W�[���;��h��I�a �	�)&��^�%.���]-�I�R�.�R�,M�_�#�-��h��޳@�^�@���h.1�F��E��������- ����<W��-��h��fu��
1dR- ���<W��-��h��;,�R'ڎ~p��C�[�2�Ǝ��|�>n�Χ��=���ϳjn���s�ےI<�����Jh��޳@3�ܮV��?&5$�@���}7���)��{�o�$�޳@�^�@���18(�Ŏ`��]-�I���0$��0=�`<���(��u4�<�!&�sj��}~z��s@�_U�\:�&$&��:��8�6�J7Vo ��k�z��%Cj8ƜML��,l�f��ö���K��h��ɤ�;�T�9��Î[��ĜB�I�n[��wt��[l�<Vנv{Ѵ��P���b�4��0	$��H�T��ޤ��+��� �٠x��O3�|��"����|(�w�h���{Қ��o$y�ےI4<̛1fZ�;���D&�wj�3�ܾφ�FɈi�$z�e4��m����z%[��	���.��nu<i�=c�V��\{<m����u�ݛ��25�̘�`��!�wt��[l�<Vנ[�S@�PV$�R1
C@-�h+k�-�)�wt��{p��<&(���ȘT�0;� �$�R�.�W8���G�[�S@��M �ٹ7��T�|Aц	�BU��"��D0���������"�#X�"�Q�v���srN{��e> �"N~x�4��m����r�h��Q)�n)��	� �u��6:�{;k�F�s�s��'mq�I�����1H�((Ŏ8h���mz�e4��<�.Tdo"q�rI&�Ǚ�zٺ���32���ʽP�/����I䌘���G�}�}>4��m����n:���0q'TXl(y�zX��Xy�6�DC�6��>�Zi�C�
$��TXfeX�B��v~VΔ�}],(HU���"��� �����*�� ����"���"��
 ����� ��
�"����@��D�"Ȋ�`���"�b* ��"(`��P"��A��AB��"��"Ȉ�"��",�"�F�(�B�",P�"�#�� EW�� EW��_� ��Ux*�� ����"��� ����*�� ��� ��� ����(+$�k&e@� x�{0
 ��d��-��h
*� U%E(P`U-5E  ��@@ 
%�  x�B�      �����@��UPR�@*QUPU)T�@R��JR�P �% K   j �   P Yi �=�S��g���P]}�!��ę_t�Q�)��{�|  �Y]n>�Yw� gT���(���0�n�:� �� �P��L��X���y<�uYj@ > @ *�D�� ;ԫx�9�v�-����@����)�}]+�smwt^�l� ��ۜ�n��{sx ;�wv����G����}V����ƻ���w]�㻶�w���;���O!ш|1�K���@ P �L� =S�1:�N-ciO ��\m���7�u�vܴU��Pp}�}<���'�Ӑ�o��ށ�`� �`�g��s���_f���rk�94v܀� �* �     �  �#�q�#�I)����o!Et�6PR�bh��JR�0iJwH w)ALm!JS4JX�)@���JP�B�Δ�,f�R�3J)Ll�(S)JS�@:R���)JbiE)c4���R� s��� 
 �(�� zR���R���hiLF��1�}���2z�q��;��� _"�  v8�� ��/���G�ӓG� ���P��'ӫ�n�r}��y ��l��   �� �*�`  <z�T�5(�0 '�U$zQ* @S�	S{T�*   �OT�0F!��_����g�_�9��?�1�;;������"���3��QEW"���EU�QEW��QX* *�����?���SU��[��Q+0gT�D(a��#�,
���T\����400�H��Z�S���})'hyٵ��Z*�TKՅ	�F����p4S��@�#pS&��
S�\��f�ܡ�!mق�<M��~\d�!��/�B�,i
bE1 F��`��IB6F$�i���kP����Ș ��۔3	
c9	�cytF���	~�3���y5��tկ6�M�e�V\p魝C/�h8bЁ\���s9w�}�p�	�cX�`r0���\Cf��m"�`��q3W��)��6o*$� ����	H�aw���yFl�`2�Ç�>a��鐙��D�Erh!�@���F���)R���)Zć횳سe
|��s�o�o�,��Θ�cX@z1,i�*���]r�D*�N���#aD�2���}yWo7c:��7��	 |nHՍYL�8��
�8��,��j"U��u
����9_�	 ! D�$
ģ8a��`����M�~�S�ve�6��3�a�q�`��Ό��a�%0�L��9\C:6.?��#N�,, �� �ā
`����1�ҩ��v::�`@$b�F���^��Aԉ
0!���5#	�6XdF1 ������ܛ4"�A;F�K4!�:>:�\2.s~H()��	��y1�6od�ypf&�7�!}!���2B� a�n!HHd��0��v	�2�B�$b` �0��0k
�$(Ġ`X�d	K�{:8�(����y44�'�zB�2aɆ%XN9�1�.�dʐ���G� y	/`�#�@J`�
`9!����&������4���	�ϖp�+!j<�BFR��g�o��R�W�(�3�^j�O��ye�����C����+��K
�3ơ�x�T�/*�LRu�A��>��N��rky� ��-��F HH0@�)ȵp*H�!O���>� p�Hr���: H��[���)8�n�)@�ܢՆ�� �G��BI��"��K1Y$J��+	�$���V4�§�x�/z��Oe�(E�ȿ�p��:M�)��a~H�#H��E�a�!\9�I"�i��`�K�[�(J||�Hf�d[�0рѦ�t��I�D�fB3>
�g40�^���NH�R���FW&e��z�+(PS�C�a>r��DF{pq^���V�j����mJAt��䌸.WS~��� gpִd$�# �,�m�F(D�B�6f3Ť�i
��V�%G�x��j�Z$xa	�N�X�6��X�� ����1��2��7L<4ohl����a"r#D�pj��i��!��>X�B�;>�A�y�$t�iyx��gA��ɨ48d�݄J`2h6�(��E�dd
fD+�b��
}��%�t#��4�$LK��S ��X��0�L����V�HI0Jk��
T�HF������B�"��B��B��S1��+����D$(B�����`�G�HaJ��ra�ZV��R�WV��ԅ�$�7�4�up`�Ɣ�
�,$��ǂ �4bÃ(lR,a.2����D�+�M����>�@�d^���5qq�a�q�9.2i!F]��y��D�N���7�t�G.d<`�A+-g�mF�5�
R�o��4dyjj��m!5p����)�<��r|��*�F�>�$HG!�k#�8R#ơ��j���W�&D�=g��p`C�� ��̗�.�u�iC7��x�M��z�Vh�������(^
1�S��8ky�@�����FV� J��2UZ�8jm]�OBBBr�uH��
�4���4��>�z�&���4o�p`0B@�¬�-���ޢO�%x�)���md1��&K�[�D����*�	� �2�Bq{p�	ÄB�p_ؙ�4`�σd,���ݛ/,a��,bG0��J�Ҥ��K��!,*�%�-�s3�$P���%��&s#1N¥I�VL���U3A�bM�[ˬ��i1�`�p@�f�%�{Íl��@$�H�BB0��lF� P�	E A���������N�.衏�1$
��FF�V4,�1��y�T�X6���Xc,K D��3�!� �`B"Tb-g 2	�$P�&���\�S�32�cqlH#!I0 :H�$B0pw1��.�#CM�����SLB�����bD�{4��E9����h鳧��˭������:p0�#�ɍl���q�4�a�
�2�d�S4�u��RWA�� ��`W |�!F��g3�c{���n'7	��� �D�l�0|d��sSZ��Kw�.	�����~N��b�.�ӿ��Ld�X����! F.�
c3F�����H��Aq��~սk��ib�Q���Q"���܇+�q*/"�e%p����;8L�S�HI~�"�=�x^���U��Ț���ki��&��2�{ۊ�yjp�����o�g�!4�Ue�D��u(|��7B���)aL$K��\�\gMC�N$���G�R԰N=)U�-�b�dCɐx=��ۗ�7
U*=iŊ��W��T,Ì�0@n7��}f��	11ۣ��X�¥2긄4�BH0BgWG���vcf��@��y�Kf�"m搔d0p)�� �2��	a�Hi5&I`�Ó&���<\d�ώ�®�M6|q��
`ˡ�}�Ò8�s�N�<O��LdѰ>,N���| Qp�!
`�R%$$h`2ü71�w$u�eO�L9HXS���,$$�� �ɧ-6l�nkf!��]���0ZF������pÙ;%LEB���-\�{���uQ.�JS�[ZS�]k���XV2�.sư,Hi!�36��^��E��
�Qyϖ���ЍcW��IC��>!��]9�~xqHP��[��qaLM>xp>��NϏ��lk�ɭ������WM;��F3�Tx\H�,"����HJ4�B|hm�D�$rѽL`��|LbIB�b�)��"š��),		"�,d!Z�h�BA��! `�,����0hs��
rc&@�F�F��0�!\9cR���
0V)�I�Ö5��d�GsaL��̄
`�BV� �|�eXR.]������A�`2�n����OR�;qa&H�6i����$��F��H&&T�@�@"`�-I_��0|��y���c�ϕ_U��V�w��#D�nڜ^Q������jc��CC�<��T0F˘�1>���荆3�I��%Æ ���Sc`�GL!�|+�wrz�����-�&�7eTE��>q0z�M�FM^�YD�U��#�� B�$�HD�b�d����?����   [@                          l��}��                                 mp�` �llإ����ඍ��	k� �E	���@,1l�R�{$���Mi��`��`m���CSamI��J�Zj��;tPn�	��ٶ��rԙkEm+��[��6���m��#m���l       � $ GQm$�[Gr� ���kv{e�Y�Z�+	��۲�*5J��٩UP�<�3jr�EUR���.��� h6�Vն� m����- �� �[p   n�I��`���   ,�ڶ�1�����UR�@��*      t�m��6ۃZ� � �  ]7f�m�`�   J�֗e��URZRZ�8$�K�3k��-�l��                             8Ҷl��          �| Ā �"�           ��                                               |                                                                         �                           �0�`km� -�                                                      �>    �&ڦ�k� �J�b@۶���n���mK@��S`��f�:���	 ��U��gRK%��&���{�
������1��d����U���H 8��`��6�$�m�n'B� �-[o[��Y&��8  ��	6퀶��8t^�h h 6ͱmIH�ؠ��n�6������N�$�5Vڤ�X|r�X�VVU�T��XW�@pi��4��vyV��/l5!�"���Ye�  8��*W�:����6n���6����I6��%��ݶpv� � 8�m��>o�6�5rޠ[�AI`*Vڭ��X6�- �f�m��n��� ���6�Ya� k�     < 	�Ē'Y�ݶͶ��4+O<u�ܻ���@�sk�ښ��%2 �N� �Ԡ   G-��[�M��{Zml��J��(HR�Y��m6�\-���u�l�6�   ���
�T���J�C��&G�Z�7ST�>�8���`�-o]��FY-K̓��j���[�z]9��Z��Z�+*�ƒ��\/N.��ix�����N�^SI��VӠCm���$&�d��6��v�,'Ei�i7 �f� � �`N��	 -�����cm�m�N�cY ylc����U;e��v-f�$���m[ ր���V�^�[u�[Am�Zm�m��
�p�-���V�i��-��ă��t�cm&k��n N�$�M�a 9�#VKE��m @�u�.ۢ	��H���-����1J���	5R�7��UU�l�<�lk�f� �E H�vImC�(Yq��Jd�iT���:[�*�d9��Wg���P�����@*˶Ā��RҰg ]V�U\^�����Iz�� ����7PRʠܲ;m�����t��m��� $[�p!x����(ԣؤ�&���A ִ�R�������]�m����&P�vj��
�i��\հ�r@��Uj�X׶����ŶӸ��b:����F^���!gn+�6ؕv�y�XK�6m� h1��\*����Y$�ڨ	P㝥�#;
����gM�H[$�U@Z;1�쒂��>bI�J-��)/im��:��H lv۱�m,a��)$��:\� z{(&�����Mh-�g���e��Њ���&� �͐��zEV�F�j�B/UTB�T�U�e���E��C���+�*��ڲ�	ͽ,��j�[c(�z��eK��r�XZ���Ӷꃚ��]�#"�T��<�X�{kq@UB�It{m��is ��m *5 T�UJ��%ZR��z]� 
v��$�B,H8 lm�`���19�U���UP��m�Κ�u�Ҥ� ��6�m��%�ٺ=5��qĂ@mkK,���^U�V�O*�@v�!5U*ͪՄ)g=%@.ʽ��F�VU�+[�����;3��r�1�[U�qt�Rn��^�
Vf�U�Z�v�(�=s��Ɣɵ���;9ݎ\f�9��Y�;
��^�[+��C��b�8KkH������&7[<�l�  m�p5lڮ �ʙ�hi\C����� ������LaT8Uh�հ��� m�R�h�M&q��L0E���m�Ͷ 5��  �6�sͻ` �e �I8$�iܽ.p5�X)jW�jt��� �6åsI��MU@m�*ҨUR���m#m�m����u�mm��}h8N�p�`Im�`��m���� -�s��h-���L�S��H�@ -���vH�K,�mcS�m�A���ZI�6��zU��Wc3@U+���P`�)P Lv6�YU��6� $ [��m%�B��jڪ���e���.vnu�\��Ҡ%�^*�N�l���$ӊ�Ν;e����+to^�'��$�d&	4�H�C
��Y|�/+X;vz�B��p�����6�b8�),gw@ş]v��P�1�v�"x��";=�I�����=W �5u�=+řgj����>���0mf�Y4hUy�"�m�*��UGYYV�������cu��s���jd$�$�n�e��o�]R�j2�m*쬑rF����<��.��B��0$�i4��,u�h-�  �b۶��m�����Yn�#u����p �a���hD�^5������ uu�o�|  8�� M��k��z{e�v�n���  ��k@]���  H �,0 �d��6۴[J٥�`8ڻcj�Ŵ��l8 &��շk����6�m�e�i��"i�� 6�� 8֭��m�	��[%���|�[m����P$� m��     m��fطY.mt�) 4��)��^j��tOl�   m�fy�ع,�쁍yU�
��n��� ��m�8�KCm�9k�t�� �V��x8Wm01����,]���3rKiz�h���[�v�k�[@����U)]3�C��k]- �P
cPpn��gPp -��E��/����g�F �n:�Uq�w٪��]�.ܙ�#^�����c�i^j��jUyeu�v�iH%�[p �yN]��m����ҭUR��i]�'d�lcb�q�p�㎧R C����U]Nt��Ur�(��qoW�֖Ԇ���}9ώ�ǠE d�5m��I���>~o�O��=��V���{e v�V­ U:*�j�v6m�Q�ԛV�L���NK�JK:� � m�UiYZڒd,�U�I&ҧ�m�]:�I� �}d$/'m��6�I.�5��+���[mѬ-�iM��h��V�i$��:u���%�&Cn�������HlUAK�U�k���m-�@��##m�9���k��m�+UUUR�
��m�8�vZ-m� �&��K#l�n���   ٶ���k *�-� *�Z�y3l��06�A��l�m�� 8�Z��hR��9����k�m� $h    嵶� s"M���`�`$�e�4�\=U*�s�*��U\���yj���n�mu+$�)m�ꮀUW��;r5BVv���\�]b���A˙�[td�(��f�I�b���� �v�]�Mmxmk]�q���`�rD�ݰ 86��d��4�ۖ��;V�H�dm̕���m��    � :��j� �P Zv�mom����m.����:��S��[Tdg�Uѩ�@l�@*�*�Ym�MZ������Zʚ���v�T�TcUW)*���&*�+�yZ���cQ�t���� �m�iq�L�I��,�KnI��a!#���;m�m�    ^�    ��	$v��mp� m�Em�vvn��	e�������]�Wj���<�յ\�[V�I�����{����O� @b������~A��誟�|�a_�L(���8;D"�}�Et��O�D��E�.� �]�	1,�0�HBJ(� �_�v�H �x'�hT`����~>!j�P�E��	�""XS����W �Dbdj,1C��mZ�>A>DS�T8F ,U6�h:"�C�%H ���|�Qh ,T�����(:@:� �F �$ HD��`H��	�a� �A�dHHQ(a��BV�$BG�
a^T"�#H$I"@��C@&z����A�,��)�Ȅ��E������ ȂW�Ƞ;T(uDt�� ,AO�w� 2 �t�Qjt"��*&A�D�=Q�C������pD�/ʈQ:�� b)� '9E8 �uU���W"�^ �DJ P ���B)�1EW�=D_��$C�ӻ�������{��w����    Z�      W$�i�̂84�rC��Z���zuM���� ��]���S�;h���>˶�.!�[�����U�tUJ��L�YF���Al�]�     �  �m��`        m�  6�  $           �     צ�      �   *�t�u#��q�Z\���O:�JA�y�m�S�[�(:L��;gc]t��a9e�-��n�A%��B9.5��-�]��p�g�M�E�ȷ� pnuKRY�q�l�m(�ŷ��l�l��e��ٻE�)[0]u܏9�.�$	p�ٞ�e�Ը�&zֹ ��" �B��um�v�:kn��M��9������a����u���{
��wjF��3B������kYD��kI��v�p`�Sq����6�{5� i�*�j^Z��O�[Jt�Y]k����G��F]��׷�PG4��jB���΍�p�5��<F®6�Ź��,��������� �Hwr]�t�Ǚ�ض�m��]�u7Jۤ]Ƭΐ�c`D��E�P���,�a���zj1����z��{n�4Ph:�
0+��;��nEunl�8����7;�v�=�ǀ��T�������]8��C��A��z���{ã���je�ie�vM�m;m�]ŷv�f�q�p�V������&��e4J硈�����:�jRRyFc�rN`�I��	�s�kZy�C���MJ69�m�X�<�� 6���Z���q���䵊�񦸧����E���q��nϭ�%Ձks��:���Q�.BeNjݺ�)r�TN5�;�U]@U����{<pV���k��tҩ\v��uw*:�S���%*����,�v���`+gTF���ג�	݉%�CucE�]�i�:ۻB�&3�����p�)�4�UW~Ax�� �W����������w{߮}�m %5�'֧��OH�ڜl�.[U� 6ٶ�	 8m�6�ފ��^�ؗPr�Op�Ŏ�W�q���7и�Ś�.3b�FO�U���˰d^��F����$���n�n}:T�T�q�G�Q��(��mK�%��jGA�`�ލ�3�.��uv�6�#d�rƢ[=s�H\��$�yj� ���{��{��;�޾~|����� >a=��E�&vys�;ݍ��>˞D��� �"���R�76T����@�Қ�|������F�L�/��h���{�4z�����q6��(�5�h���m��-뛚��h�_)����M��)�[�74m��-�M�bXq^8�I�I޹��[n�oJh�M�lM��F����N�[�ٰs��wd.g���n�Tt�=�XĔncȲ4ӐɌJd��w4zS@��h��� �ם�a#��1�c5$�y��a��(x�G�ZX��Ձ��j�;�O0rL��D�&��4m��-뛚u�������:�� Ȇ�i�@��j�;��Vd�������`�7e��rN)�3@�s@��Z��h����4��x��JF�o�����(x1ep,=���TL�)�78kl���	DA�G3@��4l��o\��-�s@�r��LMbm8h�M޹��[n�oJh�Ê�A����ss@���7�$�'��)���(�(��P���.j�JF�R�؇���`n�i`fYM޹�����8��6�nf�oJh�M޹��[n��>�ŗu`e�@��[�:�Z� Z@�����|�>Wgp�^m�
��aʭ�H~ﾟ�ss@���ޔ���:�� Ȇ���o\��-�s@��4l��v_-m�i�rj�ҥ`ffZ�3;XY����7sss@�Y|��n!�j��-�M�j�-롡�w4V��L�D�&ӆ�k�h���-�s@��4z��J�`�m�m��%u�-��<v�ׇK'9h���,ɒ�c�7kO�a$��@����m���)�Z�ZǑA�9�Ĥ�w4zS@�ڴz�h~��"�(�x�	��-�M�j�-론[n�w��cm�x���-v�޺��h����U�ui
djbm�8�z�h۹�[Қ�ՠU���D��I#RA����cO<����M��Am h �    �ږ�v۵v�!۱�6N��4]�UnNd��k��d�)A�Ѷ瞽����ҪD�wG:v�Y��w2��e��.���N�5��㋶絺Ē���k�p-A����k������6B<.��#`�a1�:۷��O�y�sI</��}��ww,I�K�10R�W�q�i��/m��y�����t�nD�h{�m�0�<��G7mH�����-�M�j�-론~��\M���5�h���k�h���-�s@�o��������Z�Z�t4m��-�M�|�V9��I��9�o]�w4zS@�ڴ�k{�"�r1�H��h���k�h���9u��	��B =v�]�����]�����Ƣ�8�b������ԧ�ț��8�M�x'3@��4����凒�����:���m9x���-v��g��/0�3�%(�UX2�
@���S{/��(��Tv��h[���L)�����-론^�s@��4�ՠ��[O���j@�/[��[Қ�j�-론~��\M�1%�Nf�oJh���o]���^�if�D�D��(�y0Y�G\�ҵ�c��ۓt�c��9���z8��#y�J`�I)��p�/YM޺�w4zS@�|�V9��I��I޺�w4zS@�e7��<�=�|��ȠƜ�LbR�����ޔ��%�Q�BUO6��7�� \��U�H�I�����e4l��{���z�� �V+D�m9x�!�^����w4��}\��;B(�}�q���ѰF�8��C�:쐝�<A�-��A�����\*e�;ܰ�33-X�V�#�7v��ϼ��7�R �q� h۹�_l��m��/u��?V_.&��dmA�G3@��M�)�^론[n�י�*��M�PL���a({�zX��grՇ!qB�̫���'%�*�1�I<~I!�[�C@���oJh���}��s�N$�,I<��j��s^�v��q��<�ۍ�+�n]$�l�+��(1�!����[�s@��4zS@����g����E$Q���nf�oJh��@����o]� �R-i4�6��5!�Z��޺��h����U�ui
dq�̱�;Q�sx��3����DB{�����˕$� ����T��h���k�h���?fy�g��?��6��_������:���M�ܢ:���R\� 6� �  �Ҁ6�,��I���^ΓX2��;�9� �
�۴�͖�h��g*v�D@��;Sr�M8������>�f��1�e��ARã�q��̙u�ك�ee����&�m^rv.��r#�\�9f.;[�=��v�vݐ��U��<�=P�W\�a�؊:�j�%{��$���9�j%^��ۚe��k�y�4�sZ/�#��-֡�n)�^�V�JY-��}���ՠ[�C@�����<)&&�IOӆ�k�o�y�f$n��X�����ݞ�BƦ���x��E�[�C@���ޔ�-v��Z���1�"ɌJ@��������X�ZX����兀.gg*�a$��Lo�h���k�h���-�s@��[k+DCq)mamdw[��<8��9��nb�;6��U�68P$i�7��r�ՠ^론ffZ؈��kK�6[)��s0����
�/$��%�DA��J��e4]�@=������q� h۹�~�S@�ڴ�댾\M����5�h���-v�����m��+|xRLMA"xcn�ՠwu��?[w4��h��/l��S�]��zh�3ٗ�4���&vv��W�&ܶ��A�m�3^����A����A@_wR�/�x�7cy����<���,�Ĥ��s@�l����������y��A��_�5��7��%P���@n��WyZY�����aV!0'�b����A�Ԧ�@��Vd�1\S$H�	
�"TeX"@ F1䤆.�G�X&�en	�0�\	� �|}Me�T��XdRT�\$ P�
�%�2�$*����(BD�E(IU�A���!.p�L!�F`0�a�&KA�i5����`�ă���J9��6�X�J!C�+����pB�����3�!������`���$%0�� �LaqZ���*Ba0˜��)p	���3$
��
0#���BĂ,@�P � ĕ�K
�n�K�\���Ar�o�!q��R�΀8�"��PL �A>~M�Ex���� ^����Wb�*
�X����oړRNs�ѩ$����m�7�6�rs���n���M��έ!FH�m�8���
�z�}��{΀���=���PJ�yö­��t��wB�r�us��{�Ş���&+u�r��,�L�{�J���‽�������w}A�{�3�>�ۘHڃ@������}V���C@��w4��§15��"J�7���A@^�R�/�i�{ε�U�c0�x��E�wu�Л�;�RM���ԙ"�#�@�_��~�7��DRE����~�����{~��6;�@fl���r"���?־�T�!�u���N�t�7��'b��4r�Vn��|�Ȏ*��ɜ�������g����a��0�����G�������C@�����
�z�}���6]��L9q����
�z�}��yV�{���6��!��j@�?{Қ3+�Oq�D�3x���ff�T���L�`s2��=	Dy.���}�����M�3����$m�$�H��^���;�պ�s=z���a�� m � ��e�3աika�c���=�����Mў�g�ظ9�z*ۑ��^��kZ^��N��8���+��n`�L�ʲ�QF;dW�v�0��N켪^{`[>a����Wm����;j�a)򕪗���������d�:x��8�U�j'==�����ļ��)Uk��ol�! .�k�xGD;��<�-��8�-g����Nbq�D���8~-������S@�l���:�V9��IUE���,/��;�^,������)�g�ߗۏ$x�Ȳc�4�+K�����7�ei`ff�X�g;�6�4)�{���{l��;��h}������|6��o&Z&��9���y(_�B^��t:{�����M ��J`ْ	8܉4�V�ź"�N����]l��t\����{hG^՗���=�$�)�L�'J�ә�L������a`s2��^(QHwg|�ǽ$̊j�MTӗT;����d%L*@��(@�!(���3��vw���{��P? �(E@) @�g�?���"�ˡ�����߫�`s��vjIG�DB!�$�ww�wkŁܜ���.3�ٖ�35'��G��*��=����XX�kQ	?�oK�;-Z�R"��1ST���a`~��п��ߎ���W���g���)��l���,Q<�t,�v�n���;��ˈ跶ݮ��H}��~����_9�y�h���X�?�O�o?�����,�w�g��n��fG#c�8�kK�Cg�9���Ͱ�9����S!���������9�-�]?y�$V"6*W�81�7T�W�VB�R�W���U�sk��������Jk&[IR���Ӱ�
Dz�!*��~�X�W��ϲ����(��%��; ��?~�̵5C&�i˪��a`l%�$��������h��h��4��x��JF�]�=�����×�,n\	]�90�;Jv���~�З�P�v�\q9����i�4|���jI�c���w���~���" ��;�^,��$<據��PI3E��c����($T9�߿jM��~,�+���BK�!$���O�h_��R"��1ST������af��^�I	L�=^,��ǖ�UJ������	�Q�		%=�����`s��v	B�
!%>���`������Ix���}��ي<��;����XX}������N��K@�[8�Du�m��D�r;���9O���'�]k��k��w{��5�*l*�a5G�w'�vw�a`}�k����C���`k͔צ[IR���Ӱ3���
;ܭ,�֖>���	zJd1z=�&dSTL��.]PX�^,�+=�z"��O��n����)219����i�-��B{ݽ,�;����,,6Q�I)��x�7���&jT���f��Nc�6!G��HP%��|����ϲ��%/�ٜ��[@4"�Z��������ދ��!� �`    e��<�xA,Nћ�.�wa�lc��.�npWGVL8��A����M�n9��':e���cNFօ��`:� �M�sƹf�R;q��f�M��q�;=�^&�+�� ��i�d��۷��w��><��s�{v;7�GV�Վ����nf*��5,�T�`�{��{��,*p� �J�lF[�ۋs��v�q�[y��M��T���LL�c9%? A`ַ�h\jiH���MS�?{��,��arN���y�X!�BDH���BK�������jUT�����A5A`}�k��H�HH�'�����O���r��<�
(D����.�=�IM�T̩rH�Q`{=^,}9���%�A�W�{������X~l�&e�f�2�XMQa�#�
Or��`{w��v���K�%>�~�4�Xg��H��#i����/uа5DG{�� ��i`s��vϟe���QD9_i�s��`W� l۞<]WC�y{C�u�oa�߾�{<���w5�����V�}���ϧ1�%�Q�}a`w�OG��4ʩ&�r��`g�X_ Ȱ|��!,��3�~�uپ��>����D/$��D	B�7���&ZtT[�,��������a$�	"" �D)�ͯ������KB�1���f$3���O"��E`B�BQ>��3kŁ�eaa��G�$XEHD�@`��u��ԓ��_�%S�jf�j�PL�`}�kb/�� H������������a`u���J�2� �l���;�]��+��ڶ;�Rkg1��.nq�\�?�E�`�7��y��M�LbR����~�ڴ�XlB�0�r�����3-�49�2�j��Nc��(�I/�DEQ�ޯŁ���h�)�g�bE\�ϾY�m6Оn���s�'�s=��ءzhP���~��ߖ�{��X�1�6�M74Xo�J'3y���z�X�s���B�n�Ł�I��j\����Kr��`g�XX�^����?���x�>��������p<�D��e�mg�3ec���@�����#��*WX�����wU�����|8neX��΀�������s@��XeX�#��E�^�M�G�(�36�X�zՁϧ1ޤ�A�N��_ۏ$x�r9��@���h�mY�G�!D�r}�`{v�X�'ܥ5Nj�J�$���D)�{�+�>�N��ԙT4��P���KlJ�����~��N�Sߥ��&hs*e��+�Nc�6�A�$�/n���fmx�3��V�^L���l�`����v�Qt����<vxci�ӯE��0��il1�[<�~�	E�s�C{�,�r6�hN/@����h�Қ��?A�"$VD"D>Ĝ�?~v���I.bj��T�˚,��a{���bF*� @
�LI���X������a{	(�DD	((X��"\bs�'��L\$c�&������4޻V�{�4}�M��0�dm��M)3C�30��0B!H0 "�"Or��`{v�X}���aDG�P�(EB+)"?w��I?{�м��HT�(*j����a`~P�<�Q��H�P�}��~�߭X�s�k4�By�vk�`�x0�G`D�����0ˆ\2�t�f�	�1p��2,��0K����`�cP�@̈IŹs�Fq���I0)�v��e�F��B��C"�6��hT��٦HYy�J0�H�2��QW� |=�����a��8�q A�	 �Y��c\!�0XgA"$��,��k�8��j��@��H.~��������e�0�f���!���	��#q�$<�(A�ĂF��� &����hr�dCAB�(��T��r®ȉ�L�@!�L`B$$�6�X���O}��?�   ���      
I��gE�ۛuL��C.�Ʉ�d�nPVp�lA�<�q*.�v\OK-�r��V�W4�b�U���Biv�ְq�`�V�    �l  ��[@       ��     H     p      ��    �,m�     |    �_hv2b��2�Yĺ]������u�9F�9vaˣk�5l�5�hI��L<0��]Z��u�v�У�� %GZvU`ڪ��RWS�W
�p�u�����U�M%@j��=�8{P���1�l�����9��Vz1U[�����i�m6h��&���mK��}:m�Ʀ6��v���h��m���͌��p�6�n�h^ʝ�,��gv�ݘ���6��ⰵ��f��ƶ{v6mCtiwf�*��j���RO����-����v'S�s��=�Wj��Pe��u���6���6���bn���&��7*�I�:,�%�v�.�G�����\�hۍ��@Qf�Әѱج�:�g��nPjy����y�	���W�ęvɵ�S��`��E���Ґp5l�b�X�#c'F�ݘ���Kգ[5\ӳ�:�Ea�ks��6��[���Tp��-����uɺ��H��^i��_l��a�����i5��4����:�K�[:���ۄ6mg��uET��Mmq�(��ݹ��jg��;n���[�2�4h�4��Gi]��1��~�>e=����T������9�nA]�&��J�Sv�z]����v������fj�ttf(�Fq��\�n�;s%^���
�S��ۚFx�6����n����CZ�s^�i4V�X1�H\`m΍�����SvƦ#n��m��4���rq�v�w!p�U*9�֬��,ﲧ���!����e3`]�L֢fL���L�"�G�'4����B�8r�<L�u��"����DT:k��s�nj�I�<WH IѷLf�xYˀs�>�k� �`8@ � ��y"�K��a�8�ݥ.u�+�)���ñ8�7�q���za|��ja�68fv��]�u�f!�m��-؈�;q�US�%.�C�!b�R�����j���E�v2�7!�c�V�0�hknh�r��Pmi|1�vWj|�u�kSȫ����ە����z��Vn�ݔ���x��L�q����nz��2�������s��?;��fZku�x��_�>̵`s��z���̭,=�+�b��LBR����FfB�S'r}�`{v�X}���;��d���"��73@��h�SO���K�ύ���� �L2ѥ��(���a�BOs/K����ϳ-XjP���v}��0L��#i��zS@�
7��\���3��,gp%
��U(%^��۳Q\��ro=�夹�>E5��]mc�M����w��=�G]N`)n�������Z��4�w4k�0�TL��T7-�+>��w0�
�r�cJB%y���g���'�!56�t��iU�p씥$40�P.��%fP3�"������`}��V}ܵ{�	(�7'e�y����U,EM�kŁ�fZ�R^�3��Z�=�^,a�Y蚙���TK�,6y	(�g��=�^,�k��(!(�n�ŀ-�{�ST܃��&���_m��/t��{�4�][h(�!������@��;�]d�p t�b�g%����#�E�p�{������r����r\̱��-L����=�^,�3٩'~�t ��_�` s2{�?�P�!~�Kj��u$̺sE���a{���!!(P���o�X�W�3���{��X&c�c��ӆ�o]��s٩�j�H��A��E�0"@�UV�E �P 
@P`c�����5$�g�ԓ��z\K�rg�ۛ�dԟ�G�b@X �U����~��jI���?�RN���jN�@?A� �?����2���L�j����OJ�� " �X��w�����nhޔ�/��kg��mĤx�%-�-���C'4�{6NN�r��\)��i<��z�_fN�9��<�G�Қ�w4�g��/� � ���$����5$��잊j���MP�%�gr��DG�@�$@��J&Of׋���`gݬ/TB�$�
$��o����9*���#���`{6�X��,��M�r��7smX�fL�̍U)je��Q�(HQ�_�~��`~�W���̵a��B"��H*}���&���aߦU$ө&e�M+>�a`~��	/�!"K��ߺ���~,��V{�ʕ[�*��^p�z�fuY�Oax-��a{rX�m�b�^��s�S-�lffZ�3��ٙkRIz"�_H{6�X�ly9��H�N����v��QȄ�ɞ��Xͯ{�j�"6v�b"�̍�x�I�@��s@�����n�}�M�_5�U�x��$CR�؅	�e�`fnڰ3�,5%	�wx���[�M9������,�2Ձ�	F�/N��j�ϻXX(Q	v�j�j���q;���z�-a�t�S`�����l � ���UJ�F��z]+�.��ͳ��a����׋�p��n��ىb`�0�ϊ��Zٮ�J6�gn� k�Z{\n��g&޽Т�Nu��u۷ h݄��Ǣ:��:�ce.!؊*йɹ��l[����;�Go��<dK�s�a�YG�K+Y�D���>J�|닲����Ju���j�
��<]���V;�����儮�nWM�Ve*���>�x�33-X��?Д.0���v�m�ѭٙ���JeL����m��e��!(��������{����w��8�c�B�Y�SjG�$�����I.�b���B���D+���_�m��߮Km��Y��2�I$�L��>q��^P��w��m���~9���s.Kmꄢg{{��m��_>���L��i9����OߒJ���I%}��ߒI^�-I%휪�<BzF
U[\q��V��&!w"�e���:'=�9ذ[��p�;���Ÿ��e�p ��or��m����|�m��e=��L��2��ovjZ�5��T�MT�6�}=��I.����+������%�m�ͮ/�����_��	~]�y����MTӚ����uO�m��������;xs��yB_��������m�k���6؟VeR��*���m�˦�y�\]��l�2�m�Os�6�Dz��o=N�m��׽332:)L����9����[-�ިQ�H���y�������jI/om?~I"�R�6d�N7@���8�D[ɻ4Q��]�DphM\����t]{V\V�n�Hn�ع�� ������m���sum��s]��)�s6�޿φ� {������Nix(�� >�=����W���&��}�����m�ޯ��m���c�m�N�'$�)Rn���ն߹�vov��g��V� 4�PcAU��'�!�?�P���>�y����v�o�0����s,��-�����TG�H3?����m��O��m��=.�m��qv�}����L�L��@�YM��g�ݶ��/� ��L���f�m����M��s���m��BQ���̽�YD��i�:y:�t���7a{:�ti�x��u�(�ݹ�N�yl{5��}���$A"�!�L�ۚ\�9�s��<���_��m���Üm��e��re���~��������]K�2� �� ��osT/$����]����l��y�������P��K�D"��y�^�332:)L����9�����l��|�f>q��l��m�����m�.�lS�%8���e��$�����|�m�mz������f�m��F+����?�?���]� ?�����</���Q�� }��gM��v��m���e6۽��v�m�8}�����!*��v�G\�+!�P��p#m�ˇ�Я�s���߾���^�Ô�\L�m����v�y�6۽����̄��>�RIzϾ<_7bHi�����{�%�Q�)�o����m�+i�m����9�BJ�US�L�y���ER�DD�M��???"��l��m�����m���5$��;r�)��I�G��/�)���;m����8�g��um�%䪻~���m�?-�R��*�u$��TU���v��m���1M��;�.�l͞&�mϹ��o��~A���k�o!�[<�f��v�d�L�H 4P�� $ �  m�mKcO[qq2W$-N��=��Ht��c���7XM����U�\^��<�@�Ź��w�]�U���p���nh�ۘ��6�u��˥�Ƶ�"�gn3�<����9u��a�o���[m��)֋iU#%g��뗭�;L-��eظ�����]Ձ�h�q=d�g\.�����/��,���8�ю�g��v~c���:��S���7m��m��'���6ٛ<M6�������\�lS�2����M����d󟒄�����^*�m����6���_�$��ݶ�z?~�-�UMT�T����������9��=}TԒ_�Z�~I%Y|���&Lm��o�(��	]���8�fϿ:��|��O8����/�%w���;m��~�C�꤁�H�!ėm�do9��w�m���bԒ^�m?~I+lM����'(�z�N�2�ɽN�ٖ��kg;r�b�9�\��f�!/D	+�|B8*��ER���:���g}��m���v�o�������;9�������y)��I�)��$��b��ǡ��T4A2��P�?�D%���s��8�fN�ն���d�(��w{������˫1�Q�{�~9��>��o򈄦g����m�/�� ��w��⌼��o��?��B_�*���m����<�m��YN�m�v�����Q#&1�6(⚒O����6ޤ�G��Y��?�m����o��� �����㘕�)G+�����u���cd���j�nh{m����q�E�	�	���3m��g��m�ݮ.�l�{����(������<�m�I��rJ�L�(�6�Z�K����y�cm��jI/_�|�~I%�K����O�4�	�n$�co#zb�m�wt]�X�������!JD)Ʊ
F�H�ɥ�HAT�F���s���J�L	XIJ�A �U(e��͑��dP��U0 �b��H$M��Lѥ"Mkaŉ�rBE�5i�\��X���@�]1D���}�a5� �/� �B��t�� ��9d$�S����1�`#��E`	!�U�$� ��"��3��ą��p�@��b؀Qҿ�A^��~N* "��!��&�L�����U�xC?jw��gV�~�ޜ�m��L�cUI���(��m���3�n��w+J��}�oq��IL����I/~.��E�F�'�dJG��I��i����m��7�)���wE�m�op��7,�p]�S�͆�Ů��/\�-��|4��o1�(���o��V`m���y�zs�����M����d�Dy��$_��5$��,�����oA%�m���m�q��v�fl�4�ow��9��e��Z�lT�.�#���m����E�m����m�ݮ.�m�oLSm%�_-i��A�F��?ߒ_5�~&�m�{�M��o��s�[G��x��B�#s������Ir��L�%%�	
����4C+X#�9'�j��s����ݭ���8"�J�(��i��n�m���ͩ�m��wg�m���m����L{�ԐD�ײْ��9"g�9���vx��㖵�����\������6m��$�m���LSm���3g���y����$�u�2���)#Ԓ_�{����z"�?M����.�m�oLSI/����X�jy&E�$��JMI������y%c����y��v�m��U2G�AD�$��Ԓ^�m4޾�@��ס~�<���h���m�D7��r���@��נ��h�N�I:)�����,U&#{���}������Y?[඀j-�b�1*BtRB�M=��h [@p�    H�l'[v�=�㦋�)�1Ip���t��x��8,b���E�4Ƶf��vzm��/�%s8�Y�"��֎�2zM�8��k�����M[q�;s���n��������ݵn4�j�.�@�P�<k/�#Ԥ�m�k|W=s�ۇ����>|y^�����{���?B(�v���b��뱏�cFi�Aq����^�`7��v]��FLCRa���}��~���=���!q�Ϲ�`[��rʢJ����� �ޚ�^^M��?=���z�Ca�ljrL��Rt�L�U��������@[����->���3�&�ܷ4XlBO��l�<ݛ ��ʰ=��/:�VI�xI� �=���>��������-��P���.ف�8��v՛���oG\m=���mxNs�Xμl]3X�<�MP�����zhݞ(y�[}��@w�'��UJ��鶛n������5��X�@�H�EH�J!P�#X�d"� �TX �+�@H��E�W�r�@?{�o�bA�/Ѵ܎	6�9���~]k��ďz�4�|h�C*�FDc�b�F����	B�*�� �o����Ҁ�ϻ6�w���c��#Xԋ@?{�h��ߋ��@^F��m�)jq1��]�x�خ8թ��z:���(nc��됷cMč�ɉ��O&(�6��?{Қ��Y�9������Vv^�l�!*�Ḓ����@^F���/6x��f����T�(�R���>�� �ޚ����%~��f�=���Wȑ"P��1F���Ľ���;����W�{�hY���#��(�Ē�V�ea`#�Gk7����; ��ʳo������ќ,�qm!�;��]���Ei��ݎn&C�s��ع��.R��PB�N&J�oE�΀/7��߉y/X[�?��������I�E�@̎�@��@ft�@[��Ŀ��������UK���Ӱ��X}����{k�=�ڴ��q6�Jy1D�9���(�Ng�����zl���¥(��<�$������+�� y�N�ɰ=I����s}V;�����~񏻶�#<��n^�V�"��Q{6NK;p�bq������7��e|�����=���31@f��@��@^���V���@{�f}�H�(I��9!���4ݕ����rl����&�D�ΕT��N[i��f�������@fF�����GX�m�F<o���<�<�r���̝�}�V>������X��Nds���ty�4�O���@��ݒFےI#jb�a����ݖ��#�X*�5R�j l H  \����f�q�]�\d]P�klu���ݶ��	Q��P�&��yu��ysĄ�Z���8�|��kvD넱ZtIǖ�v�4��'3`ѩӮ{t�x�2\i��:Y1�����r�'=��)�n1p�`��@���z{K�&[74q�i���fV��{�i.z�8T��z�hk���cT�S��=��p��;8�r�&+u�G&�	�AH� {�}4��M�_U���s]�f��9�-��N��3U`s:x�3#�����3�h�9'�1� y�N��V�ﯪ�}�h�]����ʲLC�Fa"�9��v�ٕ`w���Q���`n�g�D���	�r- ��f�����=�ڴ��Z[i���0k�rjؔ�!7Z�\�����{ԶJў�^�n�c!zJK���d���K���ۚ��V����@=�٠�����P�y�Iq�RO��{t���XQ>t��T_EӠ��77�W�^�lנ���)28(��=�ߖ�{�O���+���������ui��A�"Ls.�3;���ޥ@fGs�/�y�S��m4��b��nM�빠{�h���m��GS�H`'q)V�s��
z8���l�OnўNwn<�lG'�y��(�iA)��^�M�}V�_m�{�s@�u�2���8�4��Z}�h�]��Jh=y�T�a&Ba�@/���릥 Avis��Y�ԓ�㝺������#�2D�$)&���s@�Қ��Z}�h�H�M�Ǎ�s4�)�~�ՠ�f���sv�����Ų� 2� ���-ٺ�M�N��z�"vz���A�X�]�V�m�lz ���
C@�]�@/�����{�4�w�Zƛ$$R%���@�빠^�M�v� ���	��SɊ'��4��?Wj�m�.�%95R��U�LҰ�������gu�feX(P����Wf������(X�Rd��DM9���Nc�=��(U�����=�~�`fea`}�Nf[�$�N(�N�h!���7a{:�ti�l������{sԞ�yv��=zD�]k���m��f���s@��h��h��]T�R�*��l���;�����2{ޯ?���4�$u��ڄm�t�̬,d�;5&��ڰ33mX\ʂ�(�&G0R��Zm�@�빠[e4�w�Zbh��H�Ӱ�ʰ<��K37��n�i`s'���mr�|b�
�Y�%�*�h�j�A,D,�`�&�P�$������P"%�e\����P�@��P%H#VEʌ  0�ul!p���`C���9�s��   k      �mD$p3{i$k�d�nݦY��{K� ��^V�C���kp�,��5�,�)K�\��ҽ*i�Z��z�BT�-Xfݭ�q��     ���  ��        �          �     @     ܐm�           �M�im��Ut+���ڥV�k�vW�T�Ω3���.�����bU-����.z�iإ9ym�p�#��q�YL��UV������*�\V{n͒�;�hga�t��:ivK7�������FgA�$���Ӌ��re<���;���6�L:܆�êY��������ef7���l2l���-z�|�ڦ�P!���m6��2�,��h��[N-y۝ד�+G/N݇��^ZݫcT���LNle�NN�4;s��; =�v��7#�q�X� /\k.�ʽ���:��Ը̶��մ)Љ�S���lev��^�	�so�:<a���T��Cg�G7�g��� ����1��,vy8����������-�ka��l����jh�����8'��;/m�� ��2�;���G��66t3�'5.{pzޮQ���ю:ٵ�L�,��"��h8����m��g��7@@H]�Z[�1��;Cn�)%ʅݶ0�Iv��:���4���x�6��7MY&�#��4�T���C��qs��x��n���A˶1[--�y����63�n͍%�1l��'��'$���x.7��h�v���jy��tA�mόk����2��r�71��*�f�M�Kj٪ݯm�i^0��RA�cMɭ	.��o3������&�)@�,!ɴc��CUS�*y6��e�^�I\��dX]��7VD�jW�+Jm4��U$
��	N��.+�;��w{�������(��P�
�G��Gj�:\��8"=5~�s��j���U��QhC� �%gi7 pX`m� ����T�v��:�-U8{�z�%�(uu�����������R@�ۓ^'�-	;2���d7Q�ۮ�q�Cn��X@L��O;�����x162jbkŎ����f����m����j<<�/O>�[�Ɯ���]��M��3bqS7=�������q*��q�[���u���Pyu���l�*<8�MՌ5�6� ��!���������-����Zm�@���:�iA)��[e4��Zm�@���W��g�;2��U&J*�DӚ,~w��4���m��.z󼩓L�UERu5N�b!Bowv��m��)�~�ՠr��&H�L�%�I�wu��-����Zm�@���x��K@��v�G�F�	W&�����E�� �#g�]��;Y���Kɰng�>���~�ՠ�4.T�D�28��4�ڴ���`0R@�Z�$`���Qb ����I���;޻��S@?gyզ&���D��Zm�@�빠[e4�ڴ���&�Jx�!1)�h�w4l����V�[r���쑤 y�nf�m��?Wj�nY�wu��ߟ�EC���5�]����y]�7�i��X��Ϟ�;���]k͌�c���GW�N���~�ՠܳ@�빠[e4���*C��I䘣qh�,����M����ݭ,d�;���qҪ��H�ĉ2M���m�����<� T���@Y @(,W|�3ɽ��Zoe�p���H��24�6"�ޖ�;��31eX�w4\�/""Rdq	Hh��h�,�;��h�M������*��8��PR�WiϹ�W0<�㍐6gc�����S�k=����n�nl�X��� }����;��h�M�v� ��Cnfe��RQI�UV{ܵ{
f�ύߟ�- ���w1�# y�nf�m��?Wj�nY�wu��?s�U�bDF`�p�?Wj��YV{ܵa�b"�(S����ŏ/�!�S�I�7�[r���恙���̜�`l%w59\�L����!�=v٣�m�]�&�)�F���6��d���:��S����ͷ߿~v�m��?Wj�nY�ʸڒ��Kd�9�`fea�>��v��f���s@��ʂ�dx�Q�%!�~�ՠܳ@�빠[e4^�΢�&i�U*��sN�RI��[Vfm��)�~�ՠ�|I��SĦBbS$�;��h�M�v� ����O{�����:���Io"f�gD�Hݎ�GI6�&@� m� H   ���h�׮k]&ц�r�N�7F{�0]X�M���țqn/SI�t�n��ܥˮ��]֞f��Y�=��!N��G1]N�^��.��qv��n�;�ٶ�ql��!��F㎧u���ڋ�%�k�l�cm;[\��uM�'��k�幵MKr��L|��x�{��������ޟ�����ZX�U��d�<��R����3�gdu<�s�We[�$ly&1)�@�����Zm�4�ucʲLCȔ�Q8X��w��Ca��j��͵`gg1�=y�T�1DI�x�qh�h�iQ~�}�ā}΀���a��
 	�4	C�{�Vvs]�̜�a�P�__��a�/�mG �6	��/Nc�=	G�[�������j��K��sЂ�J��s�;�t��nh��:�vù`8�qX�mǮ�Z#e��oϮՠ�Y�wu��/;V���Y��*d���T�i�wU�J>P�Q�D�Z�w����5$�1�]I7�w�@=�$�bSƦBbS$�;��h��������sVՁ���2�d�R��JF�h��@��V�^�f�{����X�𘧃�@��U��!�j�������;�BY��x��f�z��V���彞ָ�{j�&SF,wؘ���̛��G��z�V/�_��^빠^v���Z�;�t�#�2D�$I�h��o���f6{g�v�}�`�YV�}��*j������tdw:/�o�z�,� �mU�Q�
 T#!P�"��F��H�G.`� �$h�3�RA��
`�H�,	B1��L��R�́�A�A#(r�Ux �f{z>Τ���s@��`��9Qqh�j��,�/u��/;V���Y�CƊ��UM�sN�3��������7'u��j����bƒq�ԉF�˻)�f��b����a3�*�w[^�v4�P��m�O�	�L�@��s@��Z��~�����յ`fNěU2J�e)���`gg1ޤ��)��>�o�������?s�U�#�b�h�j��2��M�fڰ7'u�����ɬS�I���[K4�w4�դ���Ps��[��}y!�w%�Zt���ɢ����-XQ佷�?����@-�����iX��&�R6��}�k���X�[�	s�v�;P��4��c���J29��Nf�yڴ�hf^I(�0�͵`fe3DLRtMEAZ�ڴ�Y�^빠^v�������d�<�,�Š���]��h�j�{���<JD�TP:U6y��Vd��9���[�����#c��1�d�f���;�6�_ ��[6s2Ձ��2�h�Փu1����|�F�mYf�� l H  �\  Li(�p�]+4n�7<��]J��+p���P��9ι�<Z9��v��#�y�$N��6Nם\yCr]C�N�v7K�vs9�� hܾL���'k]k�v�]�ד39d0;��'b'&���{:�:r�n�ۙ:�����uG�fyU�zs&�w����{��o���#<��n���dSs >'%���\s��}�q��r��d磨����d(��~��@�[��m��;��@�;ʐ�F)<�#n-�nW�u�s@�v���h��b$x�H��������ڴ�ՠz������#��Cm'3C�[>�h���@�[��m��/tE0~LP�D���:�V��+�:۹�w;V�~��.MG@2�AU���rqיJ-��E1դ��l=;!&/H`���V���OPt�Z�ܯ@�n���ZWj���8�!7>"T����J�%�_����W��sX�{u$�q��I>��zs�2���D�1,���;��@��Z�ܯ@�n��uǅ2D)E'H%��a����:�V́�̵�w;V��^w�!̌Ry&F�Z�ܯ@�n���ZWj�;�m�/�i���|>D�]	�n�Qw,lti��b-.=��Z�%���&%��������sB�ի��>�����;��@��Z��@;NU�F�4�I9�s�h]�@��U�m�߱#�b>0~LR)�
�vl���<�;p���HJ���6`�d2�#1�\�\`���ȄS!"h�K"H)�Is�4�@$p�� :Y!���AR(kx�v`�3LF#0K�w
ġ ���,f!���Bc�8�n!.0[$$@�p�6X�3�GHmF�c
�����(� F�0�/��&(JE>�#�(�E�!�x���&Ћ
'�8
q6��C`  肿/nmVR�7c���5�'	�$�Y�@�[��z�h�ա�b�K����O%<�@O#�:���;��@��Z�ܯ@����ɂq�����Ω�OFv$Mҵj�{xV�\��yٶ4�nD��?$lx�S�H�h�ՠuv��nW�u�s@���	�
E �ꝁܜ��D6u7vց��Zey�T�21I�qh�r����s�h]�@�pg:L��d�,Q���m��;��@���RpY�DȸA�5ܝƤ���r���8�m$�h�ՠu}V��+�:���/��(ō$�r$�m��8�f�s�k&:�	��#`GdmŞ�k���4�0~Ln4ŠZ���nW�[�s@�v��qgS�"��AH�U�^�o]��ڴ_U��_O%<$!<�@�����Z|�{����ճ`g�r$ʩ�]7JF�TҰ��+5����<œ`fw/4޾�0�H��x18�_U�|�D};�g�n�ڰ;��;5D�W�{�����_~�VV��:��w��{�[X�y���q�
ڀ�  �.�h,k%�������3l�ڲ	�d�ҝ��ι�GV��C
i#��\-XG���mͻ��m���ATg������L�c#��t^Í�ۃq�0���"�A�Tv��I�a�.�$z9�YܽnƜ���
���6�auȇ,[�4$C�B�-vvsf�b�;Ʈ1�w�I�	q����m�#��h�'c]��ý�ֺ��I}4��X���Hs#�I�9�r�+�-�`w��z�Dq���瀲v�U*������o]���Z���?+r� �qʹ��Ɠi'3@�}V�k��ܯ@���{�)��cp�i��-��h��^�o]���Z��Φ6'�E�F��Z�nW�[�s@�}V�k�����Us����W��m֣��\ۑ3����v�l�e<H��8h7UxG�ڵ�����grՁ��q���z�.0�z�bM��%�t�mUM+��㽈Il"R�Qe�ݻ纶l���OqV�L�0�N-��h��^�o]���Zey�T�21I䘣�h��^�o]���Z���?z�1:L�Ib�L�@�������j�?+r���fF$�7"L[�J8^���$�v����E�� �:1Z�vڭ1a��F�4�I����ߖ�k�vb��.0�͵`ne3DLR��TK�T���;�	D&Ϟ�ٰ7smhϪ�?+�:��ŒF��Z�nW�[�sOs3Ǟg��}V�k�h���i�ħ�� '��۹�w>�@�ڴ�ܯ@��2���JcȤ���Z�ՠ~V�z��n������~9�Q*�؄[s&�E;�;^������{d�a9�l��{K�蜎��x4������@����m��9wW�vW�ʐ�F)<�r-�+�-�s@��^�k�h�|�&E�!
52=�w4]���V��[��]cj7<q�M�������g3f�ݝ�`q�,��Ⅹ	Bꄅ�|. ����MI9�3g�0��rH4��@�ڴ�ܯ@����uz�%UH217����"��#��m��I2ɰ.��<��xm��t\V�#PR-�+�-�s@��_�g�|��h���ǍO	@O#�-�s@��^�k�h��^�<H�̭�r�$ʠ:�ܛ��tj�P�7ǘ�l��V>��P����PKsS`ev��+�-�s@��^�س��H�'�b�Š~V�z�w4]����vؠA�i(�@�C��D��$bR�0�(F%`�	��]�) p��?_�u�T���٧[;�h��f�m,��H 6���    m�Em�kqc-n�<�+zKu�8��gf��vŷ:��n��b��'q5�:E�Zγ���<'��n�+��t.��=R�u��th��Fcm��[��\���Ƙ�x�L�Ƽ��	tU����x��9�k]��L�;�cNĳ���[l��b�[$�T����=�wf������!�6�f�k]�ۡ��)��LSۋ��s���]n�K��ۆ�G&c���z���uz���?+r� ���Q����M��9wW�Z���1d���W��M��)h�%U�h�G�}�-�+�-빠r�@_!oSR��r���rDʠ��$�F�ٰ7smX}�M���j�;�r&\�M�EUM��{��V<͛3.��[��ޫx#I�I9"�^��M3��4���8xκ�vx�'T疎(���7��<l�LbY��r�@����+�-�s@���d&c�O��ԓ��tk*f8�*kS�ݝƠfw-X}�M�ًv�����O$�#��z��>z��h���-�s@��L1:L�Bjdz��h���-빠~V�zC��6��������r�@����+�-�s@��m��ȚMĤm��@y������n�x�9��N��q�x͓�^٬v�zݗ�5$i���z��h����hwW�z�,�cƞ)��5&h}�*�6n�ڰ5�l����TB��^�y$s%<$!y&���}��U��52��h�|@��*IM��ڰެ�:�"L��2St�K$s4
���-�s@/�,�-�s@��&�L�0�'�o]� �ܳ@���Wuz�n'�`8��O<�oV��s^p�v"��۫l�M��<`�n:&��$cO��O$�#��ۖh���*�@����ތX�4M1��J����Z��ٯ3f��͵`ۖh]cj9Fcm$�hwW�[�s@/�,�-빠{�L��ڑ��DR=޻�}�f�o]���� 1q�w�o�9�S&nK����EU+ ϱeX����5�l�����xe�I��R%o&fSn�U`:�;���-\���y�hu����qJީ�ħ��dI��w4Ϫ�-빠ۖh�w�Y6D�1,���/t��o]� �nY�[�s@���d&c�O7޻�}�f�o]��Jh��R$&5'�b�����4z�h�S@����ތX�48�$I�h���/t��owF���t�u$���Q���@��5�0���2�dHD 	 ��!R�0c!�����mҍ�t@�B� ȑ		F&R04�RH�FAciL�A�2$�Aa!R H�$X�!0��j�(P���E�D!����+�q�0�$$��R0�Ct��2Ĥ���EH���c)d�"1dL����0d!5 b�y�7jĂ����0��0`�$!2�
2��HBM�!"cD#0�3�S��X�d�	�O�&�*I9!H	��Q��JK�O���l���r     l      A2N�	d�kt2M�js���`���郇f����v��m{9T��-�2�J�s�d6��*�)<m���b�K��Z�eu �Sj�V5-T    �d�  n��K@       ��     H           	     vS`           ����kca�j�ch!&�4��6�.K�-��W��W�Ԅs��'��J�n�U��nx(.z�s6�e+fg��h��< ��\��UT�L��V�.�m�UeiG���vـT�#8C]�,�f�Y���e863�۲C������j(�ɔv(��pm��7C��� ��;���*��Ԛ�J�2Y)�K�B)z��&�������d�I�*��܍;��&� g�f4^�^�wpݴ�X0W��R�@/&e�S�M#�<�}X5ꓱ��`�s����vN�i���f�ǌL��@��u�v�D�s�j�]��mg:�%\l�L��{:c������4N����Z�۵����k�=�ک�uR��me��WEpn��)F��/�sΕ[v�5�DnL�v�{�)2ҨN��p��r���̭����vv�L�T\u�N|[ �$����F\IӒF�P�c�K�Tr�`^�C�{���Vmùe�k'�����8��W+��Xln��[!=t�M*�5�+mUUq��eY7��b��� �Nr�MrY#���S��"���l�qkH<�ې��gH�L��c=�[��8��P�rG)�a�5=`q��`�`���R��Kv�*��x�1�*�l�wC���Q�n+�!����tj.�b��j4��0��U��@,�gJ�8X�'U�x1��,PX�R[ĖUvUY�͸zyK�ki�j���ٻ=�h�,lPYA�^�mUUe�3x��C�̃g�B�Q8�A��E~P�ED:�U�d�>�s�ۜ�SL��PɃ\�RC��T� 8$ h �   l.�7�u����������훶�<�Zb&iWm�vzӲEn�n�;���u��>q-�ڴ�i�l�nÝ��gt�cv�6��m�;8-��Ck؋m.�[8�o:"�/Z�u�\�i紻Ƒ�A=��jѲ�Qdູ�;����������{������������~F��`�S�is�]K]687Kq9[��;V�`9����lp�)5�;�U�������n�_{,�=��h��)��6�m4�9��� �ܳ@�۹�_zS@��e��d�S$rL��e�����Қu���|�9��E�'�h�w4�Jh��h�������#�Ȓ�$L�/t���n�_nY�{m��>����������3M.�Wn�V��N����9�l�����Iƌr��&뵭�t�*	&h����>ŕ`}���J8�s+K�v�Z�TR�T��UM+	;�N�P�/�DD������ѩ%��4�w4��kr7��2M�n�{�4�w4�r� �ˬmG!"km�3@�Қu���bʰԒQ���`w��T˪m4�9��� �ܳ@�۹�^�M �kS!�	8܉4�m�b�&ܝ;�J��W�:a��s�;@���`���VvTS$rL���4m����;�������bƧ��dI�����Jh��h����F�Jc�UR�3��{�j�P��IB�>�[VwrՁϧ��(����̹��T$�y��V��ڰ>��V��e�a�$HLjLd�G3@?^�4m��{Қu�����m\WFp�D�]	Ot���9.�ѧl�.�s�ݺ�Թ)v��89��<��u|��X�'=�l�n%�bX��u��Kı;�{f�q,KĿ{����K����~����)5�NUV����,K��4���TX�&"X����4��bX�%�����Kı9��+��!2!wL��T�MKr�s���Kı;�{f�q,Kľ�OgI��?�����~��I��%�b��~.L��L���5�,&X�2�����p�Bd&y	I
{�^���!1,N���Mı,K��4��bX@4��ӊ.w]��i7ıL���ZSuHM�T�UU��	���';�l�n%�bX~H�����%�bX����4��bX�%��=�&����{���~�����e`�Uv��{.��<B��ٶ�+L�bs�6NǞ�:��2S*D2�R�\!2!2w/K���%�bs���&�X�%�~�OgI��%�bs���&�X�%��3�9&sL�3&[�\fi7ı,Nw�٤�Kı/����7ı,Nw�٤�Kı;���I��%�bt�C�:UJ��EH��W�&Bd&Bn-�Mı,K���i7ı,N���n%�bX�ｳI��%�b}����Tԧ5#�J��p��L�D	I=��Ɠq,K��}��I��%�bs���&�X�%��s��t��bX�!�����֡9T[�{�7���{���4��bX�';�l�n%�bX��=�gI��%�bs���&�X�%��	BظHN���UUL��UUT�4�m��g���n�l]n�[P �`8@ � �`k̜a��u�VL��A��[J�7jN�e�s��k��6�v<���/;�y12�������/&ӻA'��j��,ki�ӓ$�5��,��#t���)��]��u�6vDo= <sㄅ�dy۫\7:�5s���e�&D�#�z%���ו]p��qtk\6ww{���w��/�[,r-
���voY����ɝ���GF�6:]�Ӎv1Z�=nǥ�L�������oq��{f�q,K��9�{:Mı,K���i7ı,N���n%�bX�OS[��e��*�j��W�&Bd&B�9�{:Mı,K���i7ı,N���n%�bX�ｳI��£��Bd'��⛪Bn����s5W�&AbX����4��bX�'y�zi7ı,Nw�٤�Kı9�wΓq,��L���bMR�)�"n�R�\!1,K��4��bX�';�l�n%�bX��=�gI��%��P�������Kı9���g4�c2e���f�q,K���Mı,K����7ı,N��٤�Kı;���O~oq��������T?Z��,Q<����s��7F�秒@�7n���t�����M�SN�R��QH��W�&Bd&B��gs��Kı;��f�q,K��;�M&�X�%��w�4��bX�'��p)٪�3R1���U��	��	��svi7��ŨJ�x�� -�x�p��B ���B��e�X�)�C�(䎔���L����N��Ȗ&��}4��bX�'=��4��bX�'1�c�ҸB��RBd'�7}U.����jfF斓q,K��}��I��%�bw���&�X�A!����w�?gI��%�d-����p��L��]�-h�3UR9x�9�Mı,K��i7ı,Nc�ǳ��Kı;��f�q,K���z\.�	������a$�I���9��M&�X�%��s��t��bX�'}�l�n%�bX��u��Kı;��f�q,KĿw�{%�r�J����O�6�a��q��v�+gp�S�ҩ�6��������hZ�����x�,N��٤�Kı;���I��%�bw���&�X�%��s��t��d&Bd-�j�D�������	�bX��}�I��%�bw���&�X�%��;�{:Mı,K��i7ı,O����3�d1�2�g8ɤ�Kı;��f�q,K���=�&�X�L��T�T�`E↍��N�\٤�Kı;�k�I��%�bx�SԹ3�8�˒g8ɤ�K����N{����q,K���~٤�Kı;���I��%�bw���&�&Bd&B̬�N�PԹt9���,K��i7ı,N����n%�bX��}�I��%�b}�_oI��7���{��߿�9u�fZ[�J��Z[��������$�'�^�)��-q�\m���uUU4KS274��!2!o��4��bX�'}�l�n%�bX�w���#>���%�����I��%��Y�mxC�����c���p��L�bw���&� ����Ø$��~����H'�{��!"�'>�r���%�d.�&�e���&UT�T�L��N'9���7ı,N��٤�K�0�LD�s��I��%�b{��l�n%�d&B}�Z�t�J�n]U��	�X�'���i7ı,N�=��n%�bX��}�I��%��C"����wgj�p��L��[�6$�.�������n%�bX��{��Kı9��f�q,K��9�{:Mı,FB�7x�L��L��f��o�UK�4Q*��(�����;�]�lឺw<p�[jJ�6+���j:�m�
�������,Nw�٤�Kı9�{Γq,K�����&�X�%��g��Mı,K�;����fL�ܹ&s��Mı,K����7ı,O��l�n%�bX��{��Kı9��f�q,FBd/�.Z����T�$s53Up�Bd%��}�Mı,K��}t��bX�';�l�n%�bX��=�gI��Bd&Bzf�K����Z��9�p�Bq,K��}�&�X�%����4��bX�'1�c��n%�bX�w�٤�FBd&B�kD8���I˖UMM��
ı,Nw�٤�Kı9�{Γq,K�����&�X�%��g��MǬ�Y��;���?����`+�S�ݝ�gH�(�a�#�� �` I��| 2 ls��x��3-������z��v^j��p�3:�`�F{C��n�N�ͻ&"9���q�ook�ջv�n�)�ծp�Ý�ۉ����;F���������۠Zx�"]��#\���Qr��墮oe %�gj`GF�&��ܖ.�&��qڋ������o����ۧ(�`��Ş�d����i��l.ɋ<\m�d6�ĢIN�*�j��]��!2!l�kI��%�b}�{f�q,K��3�]&�X�%����4��bX�%�|xR�5.�t��9����!2!}��4��bX�'q��Mı,K��i7ı,Nc�ǳ��O�E1S�G�O)tL��19�T�L��V'��~Ɠq,K��{�Mı,K��q��7ı,O��l�n%�bX�s>�g4�c2e���q��Kı9��f�q,K��=�{:Mı,K���4��bX�'���Mı,FBřhZӪ)S�QH��W�&Bd+��q��7ı,O��l�n%�bX��;�i7ı,Nw�٤�KǍ��������q�Z8�l�]ke벻X
nx\v3�	�<�s�Au�\ɑNf�ْ�G2�j�L��L��n�\.��b{ﱤ�Kı9��f�q,S!2grv�L��L��ͪ�S5E�̡�+��!2!l�6n0�m�"b�@(VHA"�,�@�%!�	ZD��q3�ｽ�Mı,K�s��t��bX�'���i7�*b%��z��8���I˖UMM��	��	��w�Wq,K��=�{:Mı,K���4��bX�'���Mı,K��N��I)�eUMQUJ�p��L��]����n%�bX�w�٤�Kı=���I��%�bs�צ�q,Kļ�
\����ə��\!2!2ٻ�I��%�a�V?��~�O�X�%��g߮�q,K��=�{:Mı,K=��www����89�o�X�*�J�{)�WIɫc�^��q�����]�u�pr�kqaq���O�X�%������Kı9���I��%�bs�=�&�X�%��}�Mı,K�g�rL�fL��3t��bX�';���7ı,Nc�ǳ��Kı>ｳI��%�b{�ﮓq?(8���'�{D?R���H�5N�p��L��Y>��\.D�,K���4��c�2JO�RF��`�q�Q×�@�@�v@ �؟/Tl A�Bxh4H�H� ����3A�S�+(�o�@a��F6A��w�F`W���T ȧ�&�؁] 0��](�T���$ ]� :��-D�D�3�]&�X�%���u�.�	��쬖��t�9T9��g:Mı,K���4��bX�'����7ı,Nw=��n%�bX���ڸ\!2!2�36�:��IjfIq�I��%�b{�ﮓq,K��s�]&�X�%��{��t��bX�+���\!2!2m<����L���)Uy�rs]�q�7nlѺ��N��q�xHNњm��vz���\"fc��{��7���s�]&�X�%��{��t��bX�'���i7ı,Os=��n%�b�gY��e�H*�j�T�L�ı9�wΓq,K�����&�X�%��g��Mı,K��}t��bR!>��MK�n�ʙ��\!2�b}�{f�q,K��3�]&�X�%��羺Mı,K��q��7�2!ohԵ��K�uJ�p��,K��}t��bX�';���7ı,Nc�ǳ��K��F�H ���E�EJE�%����Kı>�{�$�i��d�q�c7I��%�bs�ﮓq,K��9�{:Mı,K���4��bX�B��k�\!2!2��r��A.�X)��7o-��9�b ����<�6LRQ��G1��t��BS�ы���=�{�K����7ı,O��l�n%�bX��{��Kı9���I��<oq��Ϸ����.�p���w��,K���4���X�&"X��}��7ı,N�>�t��bX�'1�c��.�	��	��N�MI$�3(sJ�q,K��3�]&�X�%��羺Mı,K����7ı,O��l�\!2!2g^J�qS5N��,��zMı,K��}t��bX�'1�c��n%�bX�w�٤�Kı;����p��L��[8��%�H*�j�Ut��bX�'1�c��n%�bX�w�٤�Kı;���I��%�bs�ﮓq,K�ʟ`�	bR6%dh2B��D�B2, N�}���*��Պ�W����-s'WI;k]2 $8 l �O����  m�y�m�]{f��^%�3Z@�6�#=��]0N	�{H�޲=��\��bj�F+X{9��'�;��ZN��m�i�W��+$�gu�3��k�xA54�M���16���#���;b�d����Mt���^�1&�tgZ�X̱�.�\�F�n�Y���`nQR�;���wwx�|��2�A*�ݔ�ڦ��kd�z�[W)�{zN/[:ݝ7�[��%�.�bk�r%�bX�{��Mı,K��}t��bX�';���7ı,Nc�ǳp�Bd&Bd-���9�@�bsN�i7ı,N�=��n%�bX��{��Kı9�{Γq,K�������	��	���f�"���)�ff���X�%��羺Mı,K����7ı,O��l�n%�bX��{�p�Bd&Bd,Y���:��uJ�EMU�n%�bX��=�gI��%�b}�{f�q,K��;�M&�X�%����L��L��S2M�R!AC��c9�n%�bX�w�٤�Kı;���I��%�bs�ﮓq,K��;��p�Bd&Bd/�6f\���N[���T��Hc���Wf�������nx��1�e�v��;f�&s���n�����{��7����n%�bX��{��Kı9�{΃�R},K���f�q,FBd,�=��qS4U"\�]Qp�Bd+��s�]&��j�b�DX@M��2�&�X��}����Kı>罳I��%�bw�צ�q?)p���^�Mo�C%�*����;��,K��;����Kı>ｳI��%�bw�צ�q,K��s�]&�L��L����S25.�n������K���N{��&�X�%���_��q,K��s�]&�X�%���gj�p��L��[�Z��K�A$����M&�X�%��w^�Mı,K��}t��bX�'1�c��n%�bRٻ�p�Bd&Bd.�c6�&�j
^�p��v��{9l�ˀ�;��e8.5��r��&�ڎ���{�7���{�Nw=��n%�bX��=�gI��%�b}�{f��>���%���_��q	��V�y�J����R*j����bX��=�gI�~�&"X����4��bX�'��~�Mı,K��}u�/BP�\)!2v��x�H��1��7ı,N{��Mı,K��4��c�PO(!L��N�>��n%�bX�c�ǳ��Kı/�36�:��IjfP���	���P%����i7ı,N�>�t��bX�'1�c��n%�`~���~���JBd&B����q3T��)�%��'ı9���I��%�bs�=�&�X�%��}�Mı,K��4��oq��������K�Q��*�ܞ�[�x撋k�ªlt�;s��N�)�$��v�S�UU5C�|��	��	��s��[�bX�'���i7ı,N���n%�bX��{��Kı/;��G(��ICc���\!2!2ٻ�i�~ 8���'��~�Mı,K�Ͽ]&�X�%��s��t��bX���U�j�tK�uJ�p��L��w�צ�q,K��s�]&�X�%��s��t��bX�'���i7ı��lR*����19�4\.�	��Nw=��n%�bX��=�gI��%�b}�{f�q,K��HB�	"@��)�"bH �#!'�	�D�u���q,K!2V�kN�UUB�T�;��!8�'1�c��n%�bX�w�٤�Kı;���I��%�bs�ﮓq,C{����~
���k��|>D�]�<Y5�r]��m������m��JC�5�Ӭ�	�PP�jf���!2!2w��\ı,N���n%�bX��{��Kı9�{Γq,Kľ�w�ͧSRI-L�Ҹ\!2!2w/K�Ȗ%�bs�ﮓq,K��9�{:Mı,K���4��bX�'1���L�H��ꋅ�!2!w+5�-ı,K����7ı,O��l�n%�bX��u��Kı=���"Jt
j��uN�p��L��]���Zn%�bX�w�٤�Kı;���I��%�� �;�{��n%�bX������MԔ6:����!2���4��bX�'y�zi7ı,Nw=��n%�bX��=�gI��%�g����}�����Qlt�Lk,�N�7�$(�1����( [@p� 	�� ��ē�k�L��M���<���xD��խ�G��۞����ݫ�6����ȿ�[czq���ts���46���!�T�"�Ǯw;���Gj��ݮt��nN�5=�kL���޵�: i�ذV{�y�q��dv�}�.Q�k3�����G��yG���e`�Uv��Z�3��1s���m�� �w<&'8�l�5�==�nD�rn�'�Ȗ%�b~��M&�X�%��羺Mı,K����7ı,O�w��p��L��_v�b�T�D�u"s7�Mı,K��}t��bX�'1�c��n%�bX�w�٤�Kı;ܽ.L��L��`�Z�S$�P�L�9�Mı,K����7ı,O��l�n%�bX��u��Kı]��w�&Bd&B�
Y&�B���q��Γq,K�����&�X�%��w^�Mı,K��}t��bX��������	��	���3i:u5$��c�ɤ�Kı;���I��%�bs�ﮓq,K��=�{:Mı,S!}��W�&Bd&B��jt"��hUm�[�u���6K��;s���6�gzy�!:pb�gl���Wg��[��{��,Nw=��n%�bX�ǻ�gI��%�b}�{f���D�K���k��p��L��^�-�"Jt
j��uN�n%�bX�ǻ�gI�D6+s�>QӸ��bc�����bX�'{�zi7ı,Nw=��n%�bX��<zA���J*f��p��L��_f�.�X�%��w^�Mı�+D�N�>�t��bX�'q����&�X�%��*Ե
\�		Ni�\.�	��{���Kı9���I��%�bs�=�&�X�%��}��7ı,O��lR*���n�Ne��&Bd&B�Vm�n%�bX�ǻ�gI��%�b}�{zMı,K��4��bX�'������g�*�O+��C�ڱ���tk�i�]���s���*i��K��G=.j�v�7I��%�bs�=�&�X�%��}��7ı,Os���mȴq�Y��b�
t�D�&�'*��2�k:A$M��j'�%��w^�Mı,K��}t��bX�'1����n)��	���3i:��d��̡�\.�K��;�M&�X�%��羺Mı�b�D�"�t* 
7q1�wΓq,K�����&�	����7[�34U"S�T\.	bX�';���7ı,N��ǳ��Kı>ｳI��%��&"~����.�	��څ��-S�SU5#�zMı,K��q��7ı,O��l�n%�bX��{��Kı9����p��L��O��[zԎ����eWN;o4�۵�^ݎ]��X6뙶��%v]v��`7/=l��9��3�������ow���&�X�%��g��Mı,K��}t��bX�'L{�Ɠq,K��ѩjr��'4���	��	�����I��%�bs�ﮓq,K��w��n%�bX�w�٤�Kı_mn�"�����D�sN�p��L��\�{��Kı:c��4��c�!����~��I��%�b{�}��7ıL��`�Z�S$�P�5N�p��LK�=�cI��%�b}�{f�q,K���]&�X��A F.�K�*TZ����*���\!2!2t�B�:��AR���q��Kı>ｳI��%�bw�צ�q,K��s�]&�X�%!b�͛��!2!d�)�f�K&�hUn�+��փPua�؃�6Y��+��d�f�5��ϭ5�.�C��7|�~oq��K��4��bX�';���7ı,N��}��'�1ı9�߶i7��	��8�ܩ��h%9d���p�ı,Nw=��n%�bX�1��Mı,K���4��bX�'y�z�7!2!2�o)j����S�\ı,N�}�&�X�%��}�Mı,K�Ͻt��bX�';���6Bd&Bd'�Z�0:EI4�EMM��Kı>ｳI��%�bw����q,K��s�]&�X��I��3���.�	���G��r��'5s�I��%�bw����q,K��s�]&�X�%��ﱤ�Kı>ｳI��%�bo�T2�O9�	� (YaT�I%E�ԔP�e�DdL"c* �I����l��	DԙF��m��0H��ā���0n̛܃0n�BI	��AXÜ�����"dL����"1F p�&T6A$B���(�d6;#>�5�     �      mVm��I\�6�ف�����M�Mu�&;# *�v�
!=��+��6�K{.�\�52o
�\�4k��U
U�R������-�     ��`  �P        6�                @     9o       p    �6��$I0mE�a$����3X��:��v+�:�^���6�;kc:$9�MARl�貼t�楪�!�N�ўSlp.v���:ۇ]	h�tT�S�c��;,�KUf)6^�K]�T��Ű��Z�n�@ӑ,&���]���< ˅�Ȝ�%V:4�{d��9�g.�F���2��9�ɳ�	�m;g��W��@ܚO[i�l]K���{q���u�VyÛg9�m�[7\�%\�O:M\"�2��<%гqur�b�l�����I��H�}��.�pl�\a�4]h�'m�8�"��m���=��{-��M��J�Ѷv�iF�@����nƬ��K��nܜ�ͷm�5@ݞ7i`�$Л�����"P;i�:�A��aMc[��"v��$�J۵m��3�����uqR[#�V�[�hUCb8{aڠ�.��Ĭ[R�n�����^m�cۓv��p덋;qdwT�Cl�n8���d���ׇ,�����]�f۰m����6��-Ta����z����ܶ*�rvkC��9S�z{�X`9�f���m��t�r�K�*�\6y[�n8�@�؎yN���f�僕Z�b��Zm��ں��G��V��!83� L\�1���ԛm���lH7\��\�wq�lh&�'��e���f:�ƙ��eN��;2�t����.#�ʀ�r8���nt�-EM�"uﾺ��ӧp�k"�BC��r�x�]�����*��S; \����U��먃���� �S ڦ��9Ά㱓9�q��T^�Q ЏQzQ6��ɕ؁� 8�� Р06��C+���9�1�g9�s�g8�)����	��]X`�� m�  8� m�Ydu�Ē��� �d6N9q��a,c�㋡�S3���0a'9mV۞u���l��'�/F�75SV��Rc&\�;e+mu����+�q�>g��ۄ�����䍩��M�W��ul�E��gr��Y�~��_3à���:�nW��l��a'Q�w{���T�,Q*�؎�]:��Q��.�n���s�3��K�+q�+���j:��c��}��{��"{����Kı8c��4��bX�'���i7ı,N�>��n%�b2ك�-jUL�UB�T�;��!2�=�cI��%�b}�{f�q,K��3�]&�X�%��羺Mı,��_a��:�S%T���\!2�b}�{f�q,K��3�]&�X�%��羺Mı,K�=�cI��#!2Zfm2��t�[R�i\.��bw����q,K��s�]&�X�%��ﱤ�Kı>ｳI��Bd&B���d��&�S�MM;���bX��{��Kı8c��4��bX�'���i7ı,N�>��n!����}�}\����
Q��9۹�6t=�㍲fpb	��"��$��FCc�5$�N�MTԎ��.�	���w6n�X�%��}�Mı,K�Ͻt�Ϣb%�bw����Kı/|yx��H�&�h���\!2!2��l�nQ�"b%��g޺Mı,K�Ͻt��bX�'{�Ɠq?+��!2��%�1��)�Ni�+�� �,Ow?�]&�X�%��羺Mı,K�9�cI��%�b}�{f�q,��L���lR*���eH���;�� ���D���I��%�bt�~Ɠq,K�����&�X���������	��	���;B�R�d��I�g7I��%�bp�=�i7ı,O��l�n%�bX��}��KĤ.�f���!2!owS�ɤɦ�C�z��6��e���m��xs�&c�����6�k�B��p��v���f~{�7��������&�X�%��g޺Mı,K��}t��bX�'s�Ɠq,S!2Zfm'U.]*�ԹC�W�&%�bs����q,K��{�M&�X�%������Kı>ｳI�����{��7��~��r�\<&f>x�Kı;�k��n%�bX�1�{Mıސ$� �d�R�L)V(�E��(P<Ptj&�c^��&�X�%��羺Mı,Kq7�$�N�UT�4\.�	���9�cI��%�b}�{f�q,K��3�]&�X�%���^�Mı,K��V���*���:��\!2!8�{�٤�Kı9���I��%�bw�צ�q,K��{��n%�b�����=��!�j%^��ًUe93v0y�9�V]�GW#u�5vU�u���s�����n%�bX��}��Kı;���I��%�bp�=�h? O�b%�bs��l�n%�bX���~rL�L����p�Bd&Bd,�^��'ı9�{Γq,K�����&�X�%��g��Mı,K��!�aT�55����p��L��Y��3p�AbX�'��i7ı,N{=��n%�bX��u��Kı>��c�4��((s3UUp�Bd&Bd/�7��r%�bX��{��Kı;���I��%��� �P�T�0$bG��VD�BHE3��η�cI��%�bSӽ�K�����-1p\c&�q,K���]&�X�%��#�����%�b{���cI��%�b}��f��g�U}����)�c�8X)Uy�rs] m׀㫪ۮ]dkQ��{$'k���mv-څ���31����?���o@�z�hޔ�*��ք���$r�@�}[�?^����4��4�˔i
�A6�o@�z�hޔ�;ޔ�;�V��.e�	��bc�4oJh�Jhϫz��s@���L$Y<���N���oDP�Ԩ�(_~�UUH�D�q��i�ڛ�n�>�$ V��  ��p  6�4��y���D�Ү�9��m����.輻�A��솧1�����ذtu����J܀��v�uֹ��<�nt�
8�b4�݊Y6��{Z�_��@�Dml�>�v������\a5�^�z�G�7N�w%<�{i��:{.vth�&�����xm�$���]v���m�wa���Ŷ\�8�ۍ��C�6�e{2�ts��^�Uoͷ߳�3`s;�����������Ic�8 �nF�׮���M��M��o@2���ML�,i�nf���M��M��ށ����?*ajm6�S��Ԇ������홰9��V�BO7/Kuv�Ij�H�#������~�w4oJh��ީ'�T�`�m�"Q��x�vڪm�K���C�J��{z@Ş�u�:n):�nU!@�PiHށ����:���޾�@�u�h�\˂p1���&h�<U{�O���ީ�r7��7�h�w4�Ʉ�'�"3i�@�_U�|��Uf�ۛj��������Bŏ#�$�a�@�u�h�]��Jh����b�T��X�nI�s;���	f���3����s*�ߪ�}�\'*���,���7g5�7H��[�c�9e��s��A��1����^��;��h��M�빠~T���mȦ'����}V���d�?^��^��-�-�ƲLh���ˠ1�t�}�J���
�I?<�N�S@���@=�A��	 rI�~�w4�)�w���=V�4�.e�	��bc�4zS@�_U�z��h�]��3ߧ��@��d��Wn9ޫw�8\�s<�yN��8��m`�Z��o]����Fߛo������3*�gr��(�0�����dɔ-Y2<RO&ȴU�M�빠[Қz���r������rM�빠[Қz���m�@2�֓��M*m�r��
Ow/K;���I��{��N(���b� �!�A1�g���I>����1q�eƓ��Ԇ������ɠ~�)�Z���<��w_��<�H$�r$�m^���c�u��#Y2�1��6�`��+�jL��v��2$n�����4ץ4_U�w�)��\��m�a28rM��M��h�Jh�l���2���l11�h��@�zS@�[d�?^��;�o�	q(�M�������ɠ~�)�Z���_&�ʱ₎0�C@�[d�?^��-}V������]�LII$����Y1�
��X6c� $ � �   �`��/��5b��l��5��44X�\={uMF� 9����=Src>K���^�z��.���y�q�>,��V�(90�r����]�g˛&�
�VL��ͻH;��6I��".(�g�q��9�6ok����)d2���j��#7i$)[(�uG���o{��>t��Oƾ"S��c[�����F/d�rq	�����6{f���8�@�8�&Ӓz�_�4_U�w�)�z��h^]f'Ȓƞ&�h��@�zS@�[d�?^�����a�ɴӎD�0QŠ^��@�[d�?^�����-�-�Ƥ�9�n5&h�l�^�����:���{/����dpiI$�:���-}V�׮��ɠ<�ښyG<���U���W�;���Q�NŶ�nݮL<��7X�����L����&93��Hy:P�b$��TdozQ30(���"%��<W*�Z�����%vS�d�=�w4_U�y�x��İ��&F���$4_}�����k��Jh�׸�G"CN2	��g���P}�;6x�1�t� +��,q"B$��������/�)�z��h޻����6d�N7"M$���-ٻ�k�ڔ������p5������c�;����RF�&�Z��4U�M޻�����gV���9�m�@�[d�-빠Z��ޔ�{/����b�4��h���-}V�l^�"��p��A` J&Q�HiR0"@`aHa!�eE``1 ����.7GA���&�2�"H���UҀ@�6�0�&	���#c@�/Q��$@�/�!X,F FH4L!Ha���@wK��
y(H���d#�m2A�N�~�,`��@R$I�� ��8���:��Ba��!p�DH�E�0(`�v$3��Y��>Ch#�;5�h�\���%��H$b�Q���#,D��"D����'t� zv��ޗ��7�ʪN(��>DڀuS���P���|Wj/m�/x^�Uo*x�-���}%�bn6��4_U�_zS@�[d�/�)�r�ǅ�a���qhޔ�=V�4�Jh��@��m/�lveZ�W��q�n�n:�0F��/bLS]���O��^%�v9l�=t�mϪ���l���4_U���}�|h߾{�$r$4� �NI�_zS@��Z��4U�M �Ƕ�H�!X���4zS@�����ɠ_zS@�����i�#OCR��4U��u$���f��S�R�&Pp�WJ��E����{=�Ԓ}��(���0���h�l���4zS@������fx���4|�(�R69_iǹ��4`^�v-����
��]�]��ˏ��m�dB�4��~��@��4�Jh�l��˙pBo'��&7ޔ�/�)�z��h޻�+|xX��%<M��Қ��&�}빠[Қ��,8�&F���$4U�M��s@��4�Jh�׸�G"CN8�6��@����-�M�Қ��&���<̹ݶH��UH��j� �z�ݖ�C]׭�
ڀ��  t��U��ю��z�4Gf�.�Ӳ\"�mJC4�2���q��۰�c����{�9�n�jMغ���hmAZ�KɢKI9տ�|�G�
�cY�,n�r�n�s۵���k-���ġ�&�x���^jv�N�;`�A8F�ڎ�[��`���e�������鍓2� �ݲWe{D��GM���ƿ��=����	�<�$n�F:��-��볿2O��kŁ�v��>y�U�P��{�j�3��&�MIx���/�)�z��h�rՁ�����-�cs5H��7��}&�}빠Z���Қ�|�i�)�
DҒI�_z�h��@�����ɠ~���&�x�bc�4_U�_zS@�[d�/�w4������C�tD�D��e�t�M+G��k�&�n���Χh+�+���{Qd�Df&ۋ@�����ɠ_z�}�~A�����%�>y24G~I!�z��s����*t ����I;�9ۨޔ�?u�qd�D��di�4�rՁ�=�fM�r��:�v��>V�O#�ı�������/�)�z��h޻�ެV��MIx�qhޔ�=V�4�]���h��W?G��X)G+�3���E����q�ፉ;Ll���ؓss���ݎ�Ɂo7iP�4U�M��s@��Z��4��h�lS"��$�@����-}V�}�M�m�@�Y|�!7��j$��@wF�;6x�J��/$�1��h�����(5�!OmŠgݬ,�fUX�rՆ�J�f��İ��&F���$4U�M��s@�l��}�M��渌q'ip]�fٻ�[d^ЂG\9�#<��6rq]s�2�����G�N2		�h޻��e4�Jhu����byH��)�Ұ9�X^�6or���Ҭ�]� �V+D�ڒ4�5���/�)�֓@����-�M ���$�`�Cp�m&�}빠[қ&Ԡ�H&AW� 6c��Ԓp�A��2!8���/�w4��/�)��&���Icĳb���Q*���Z�)�-�&���]Y���uv2�j]�WeY3&$ۀ���	&h�)�_zS@/ZM�n�՗ǅ�D�k��{�4���/��h�)�~��a�y24G�$��^�����>K��|h[>4���H�Hm�P�ꊰ؈{��+{�����a`�&�g��̏$ix���_l����;{��;;�PI%k^�R�UTH�K��$�rc�U��Y:;@�]� � @ ]��V��qi̹�.�fm��j �m��\�9��Z��k��ɖN��dݎ�p`l�=�B���XN7V���N��a�3��(=]�y�84�=�^-$v�X�yy��ڍ��\��^���/B��۳�;�0g�s�D�����c��n{Q9�����U;�zX)T6��s]��#pZ�puf�[����g�;\5^�c�8�EJ��6kzקƀ^������e4�3�BI������&�}�s@��M�Jh�|�i�)�	���&�}�s@��M�Jh�I�~�ı734�Q4MR��{������@/ZM��s@������pQ5���@����^�����}��6��~�����+<�]���Sn_<�vN�w;;@8qϳ���M��^�֞�M8<	$4���/�w4��/�)�~���Ǒ&���!4�]�Qb�U ?�5��{>��}���RIz���; �Fб�����)�_zS@/\�@�����Ԛ��R�S�TXyB������75mX޻��)�ᖴ$���hn�ŕ`j�������ZX�k6�?�ߠ=�n��PJ�y�MM��H�<���s^�s�s؎�,�ζ�1[�VEqX#�&�}빠^����4��4՗ˉ6�!�D�����/t��^�f�}�s@����dx8:rәsE���a`��Y؄��E����H��{�jI�s>��}�"Xq^L���I!��M��s@��aa�{�����6�SN\��A!HM��s@��4�Jh��@��m4���MĤm�"J7ZR���6�P��]`��� sG,⌞�c�i�=��hX����ޔ�/�)��M��s@;Ԃ�1��Q�hjC@��� ww@voR�;�x��^I&�uvX۪$��e�i���V}�y�[Қ��he�ѦؤN&G!4;��y��ޔ�/>�Bf�c@e���@�
�$ȅp�d�9sU*� [�@(x���L�I�<���0I�D��ޔ�/>�@-������u@��diĤm%.�s�V���$;��9�\�\�;<�Fw\㜵��Ϝ$PMbm8h�U��M�n�oJh�bXq^8�8c�9�[�&�}�s@��Z��o���${O�oq�X�m�d@�ɠ}�}��Z����޹4?^vA�"��d�M�+P�{�����vgqZ�ԒIC���Xu���2�]Jrɩ�`gg���I���n毗�nm*���u$��(����Q_��EW��(��DU�EU�uEW�"(����*��(�*���*��QDU�EU��"�DQ]�(���(�*�𢈪���"���(���(�*���"���"����
�2�Ή~��I��������>����a�B>�%H/�       @ � H!��ˮ�Rی� G��bk��q�R���R�ۀD҅,f��ҹi�&��X�4ҹ� Х1��c)���q�� 0��w �a�      M(���UA4ba�i�LF��� b)�m@��MCSL����0M4d��0��	��i� ɦ�����TASP       3PR���F�FL@ddb�@B@�=LCD�S2'�5��]�w�x�^Y�`TDtD���"=��J�P<��"#e	�������+�E�,"����ਈ�Dps�Z�TBHBIc�N��S�/�������y�m��x�@                   q�q�x��࢈n"���{�<�ů��J�O���4㺾���}=�jߕ�����Uj��ZH��ʭjJF�(d,DiKF0)A-Є�kt���;R�@դ*,l��ti$H��5��d*���k�T�T!z|�b��-F�`�
�U�®�.S��*�1Z!��Y(�WQ�Uz&�M(�Dٴ2o��r��b�
�O���ҷT
=��n�HcC�4C�
K
lƒ#L���!�Q��HʱBA�$ Ġ�0F�Mn�q��B�F��\�A�j�
6\��j"�b�"��В�QUuj���Z���T��)T��j��� @��H�1�5�$�4F�T
H�FB� A� H�#���$ V�D�1�Q@Z�I� F��SA�*�UJlF5q�ԉաR\
���M�M��IfUp������$uK�@�]�}��iR.7!�[�fY8�"sw29�y������yu-Of�~)l����i�j�.&bj�)wwKׅ�U��s���mA�ol��Uf���0���������#�EF�;�W�b:�(݋�q��Z��{��                                                             ���                                           k��7i%�Ij�6��fۤ}_K}z6m��e(�mm�Ԑ6Z [L��l�� 6�E �I��6�v��.!�r�sl�                                 A�                                                                             z@       �?Co~����-� M�e�5���m-�` �j�n�m��dI�Ý��h�ޣ��sj�$�涎�@ٵlm'V�[rA m��'�&���M��$k���M�6�	 �U������p �� ,�i ��mmm��l�l4m�����ձ*AĒ[@m�E�L�z�C '�H��m�ޡ�$K/��=z��,�my�m�ld��k�$	t�` �d�n�ے� Y@�.�GP5��nu�Z<����zJm�],^͛vt������e]m�m-��E�赕��-����n�L�E�ݚ�-�ؒE��RȖD1t٧$� �uZ�F��ju���6�\4ݻgk����]�3Ӫ�Z����m[""�ߺ�aU�'�qH��ۿ?���"�a�a|OC�K���x�p.�A�<�!�l���P�P��m���	��L�6'
.�P�n�L�B�.�:L	.#�G	��DcA�}jt%hB%@�TF �]s���u��8I
�\f���{�          m�        ��mmz�h�tQ&"�i�      m�              � 6]q6���:Rk��*g�ɻ�d�U��[�5ۚ+��Z�,�^��۵�'k���yl��-�n��u�%g^�Nt�.����y-x]�/W��{�B������w��M������ m��m���m�  l���q+`�Mf䮻�.�;ci��ډii"'�?������?k��e[_��+�}�t�mu���[}��6P�
fX+}�s�E���E�����NV5�o�u~�}��¬�?`)	`�F�+�y�t�m�w]+����dY��-voqb�mf��6 L7L�	��NR�yX�o\]��9du���}e���� �Cd)��m��n��V�'+zr��s���s��      ��-�`   vi/5��m�"k%��;`��HK�����gW+�����я�V���,����6 LKDL���~������㏣���望Z<���z�n��{��V=4����Kcn[���ݖ��=D{�yc��yו�k鵷���
BX �%�LLwV�{{#��F�+�ß]+ǜT�����	�l ��J�$�f�V�7��X�]��ۜ�"� [�*o�    �FY6    �뮤ل�]ڦ�jr��	f�c'�gT��c���md��u�ݽ�\��9���C�	ʿ�G��.�ʈ��޸��纹\�N;�-T�ep�HK %�$�<vv�b�o�}�EoVy��͎�v���GfPt\�/kF��D� ��W`U��Rܲ�D�!sb�p�jUWYƵ��S&�v.� ��GDx�*����^@�_�`�^m��D�6 &�`#kA��+��=�n-�6���=�{sK�&�i�}y�wv���?��(�r��`�N�S^��^E�<�yU>�lebx���ʌy�(��     �l޽u�n    ,gk+�-�����&\6�b@�� LKD� �_u�ff��6�^o�sκ�k6����y����6~�	������舼���_�d &\EIi��,�����tGwڷ�&���@ku��sε5�����m�L����b ����?G�/��ͻ���L�`5��~��*k^	��'��_�"<���
�v��M�<L�����w��&-�]l��#~ŵ������ )��Dg���n3�������z��W � ��A���ۍLn�i;�uֻf�i����Z�q�/��;�\l(�+f����L�`�p(�cCV^G_������?G|�5}p�����dwy�]h���)~9��0Ρ�o�����    si�    6'6u��sշ5�n�r�`��H��#�%3ue�}-4������I�ڔ����Ɲl\{;�i{#F�=g�N��}^�HK ��w5EFU�c�o������}{�nZ�s�e=��Tn��R��.g/�&���| �1,�;�ʝUOv�k�9U����{ϻ���Μ��=齊s�ln߻���v ��l�t�kM�߿m����}��k�8�d׼g�wo��=:V笶w�HK �[i��oskf��kv�����l^����YS{�}�݇t����KA4�&&�T#�b!
�A�9�ݡB!2��_��t|��{�~                     9�t�����-�miK��Ө                       չmd�ݬ�\ӪV��]&�S5Y���l�֍����ki��Z��맒�]�%�v�KI�Y�^��L��lӷY�곙'[�*ަ�y{u�B����:D.�����x�� ? � t��[&�   ��݈��z*�]n6\��M�l�/ S���W~3���>��M�]e��/ߨ���=jo��c����{� ��C�ݭq�e�qG�_����~��y���VR�y�]�yn����R�`�SSQ�x��;O�}�-��_Ӓn�ڒ@ӈ��=����vw���B�3�w�&A�bY3(f�w[��ǙU�g��nڛ��6j�w舊o���6�u_����I��YW�O��-���]{��ݯR���m�m���mN�T��o�    �a` �z  n���gm3�f�n��~/<���^��6��������ӅfT�y���9�{uY������ڟ9��� KN���V�׽��O��=]|{6Լ�[�o�}��mMw�
̥��L�`m!��笿��24�����|wd���/�_}q5�f-�{~�m+�6����/=��d�l�3#��;��o��yt���ӅfR�^����^�����k6/*�Ǵ��H7-���Y疱ѕ�����=ڥ�ajc�j�{ո�ﻭ�#+�     �i�t�    ���TJ֬4�Vr�m	���;���Zl�s�����]k��w6�}�k�߹������nބ��啘mux&A�> jf[M��{-l�{�4�wz�w��ko�;�ͫ��eGQ^{w�ή�)	`��-Vu�㝛�uz��5�H��Sa�JTJaE� ��3w��� XR0@I@ @"E� �Hmz��>�E^�?g���RI�i%M�_'��m$�$�K�Wѻ]�Fٻ'g��2��S��2�]�ӻ[U�識����mn�.HM�!I/{ﾈ���v.���w� P�@ ŕ�{��Y���R�x��FuR�TR�g�j;�Qj9Aӊ��Gݶ    ���$�    ��*p�۬���k�n�����wCעR�J]�j&�K������k�̏
>��Ƙ=��}���^.a@��7	�X�_b���?{d &S� [�áxvY�gĽ��C�$�0�P�������^�;8���o�M%T\(�x���j�rdƯ��΄� 3S$�U�B��q����^�ñY�ѸC�H���Q�ÅY��kÑx���~O�P(Ő������ S2���ׅ�ㅂ������"�������;�)ﶁ|x�/'�����E��ʣW֣(��޹`L�uUU
&� ��!�x*�n�r-x��^
�����tZ�mG������Qj-|�b���     �d�    sc��4+��U�L"��Qi�:�3���g��i��O�h���
Ǔ^�1_�I"��]іBFB��}ݸZ�D
*�b���HK���0O�X��آ���:-iT`�`�z|�'���s��z+W��m{��^��m�X�T=�v�)	`��B@	�b�IF/�Gt�)�#�P��p���I�׵#�O�J�����՝�o���d�s��(l �n�D}�)}�����1}ii²B{(
ǂ��vqkGFE�,Q<=�?b�~�O�����Jf�4Z�ȴt/|K��у�};�ŭ�GB���,�<��t��yW3����6 C�����|W_�[�Sﶳ&\��                       m]T�e�i���k��^��                       ҞE�5�[-�*Z�ۛ-�n�ɪ�K�`�4�mA.i9zۦ�eM�K:�.�w;!v��.������.�&�ɸ���5[(��SiKIb�K�XӴ�F�mUUP  I)���    �KmvIlȳ�k�];o������%.��z�w`�V=7��Z<���d<�f³�un��"�мM�/뇪)}���d &�$�&�ԣ�J=gT��j�GB�]��֏"���hx+�+wo�*0Z;�pL�`|Q2ا�P�֠R����F'SR��P�V�/EB�[F�����شt(�:�x+`�u��"�&������*��֏��Gt��ك�X���֋�E�ث��!ડ�-0�ﾍ���ܪ9|�b�P��x&A�b&��QTK�Q��Y�e�Z�شt.��jG�܇��E7�鵃�h���v	}���֠_8͹��      :�et�   �br�����tݚ_;�(Zl��1��{�{��>�ق����G����ۅ����^/�x+�p*��E�ءX�x/g\�TUE 
Y.\11��E/�@��7�F)���8X-8V)�����q��Z��/��隥?]L�QK�}� �1.��UTZ�ȴt.&������X�9�kG��э�$m�I�Ma�"�E��P��6�PG"���UUUU������x+~5
�?}��<����"l����FD>����9�ZM�X���^��WEc/�UUUSUT�eMMF�G�У���xx��qw�Z<��'�h�Ǣ��;�*�_{�qƯ�Gx��      :ɳ�&�   �ē�n�,i�[�h�{�·�D���r�_>'i��T%�}�Z��xv.',�
�����t]8��Q�:�x+
�
c��d &Rd `�1}j1Z�P��C�[O�T&i��QB���kE��E�b���!�x*�}�Z�ȴ\X�b���nHnS����b�Q�u�kGb�У�OL.4X-_��)R�\J�Ei	� J$H!�J,�v��ݪڮw�s�"�V�ü��G�����V8��^E�*����v~�����!, ����\j��h�]іC�	(X*w{^�h�^&����X�Yɲ���a��B��~��i�/mΪ��{��y�ry_?]6�\h�X�ɾ��������8�}�r/�te��R<�ھ�7��  ���`    �]w4����l͵�k�y�6���N��ة�V�E�мM�/C�Qb��赞����QvOL<�C��t���B��Q���� )	r�ME�������8��ojt�*�vG�����K}ۅ��t-����[p�VI��d &�$�&�����R}0��$у�X���֏��5Y���m�,7�ŭGG�2o�d P�K�lS�(k�P/��-T`��h�^'8����VX���֎���O�4��}��0�+,X+�^���� )��5}j1|(����+_h��)��Z;�E�d<��rWn)���F/�}��      K(��    3�J�&CU��Y��r/ǝo�^�M�z嗔�ω����󺳋Z:��Ƒ=��0�V=+����6����x(���V>�V9��r�  7U'�Q��R���?`$�%=�6�HW�{K^�áu�&��W�X�)vFqkG�r�9��J\2�m�|�;�����>~��GB��x+�_6��{k�ŭ�z/�}d<�H}��QS ĲT�u'�Qy6�(����m��^�kGG��d�Ş4Z:$�^Ml��ޛ^�axv.Ϧ航� �,$lHQj%}j�O���1Z�Z:8:2�x)�+�}�-xr-C�ls,��ax��A+)"�pvX ­B$�٬���;�կ����||�                    K�Eד�ɵ��:mpf�LH                       ��:@�*M�e��X�R�ͣ�Nؐq�4Z�����5��[��kɏ%.m������i4����CK��qmnȖGiț����v�Ϗ;��<�=w���   j��@    ����-��ܓD��v�+����������QG���z+
���6�x-
;����X�t���h�_��_���� &$%J S��k�ߦ)}��������Oz��N�/C�P��g��Q�_�)�'釾��݅�����"�f���4����^GC�vP<�C��qkG�$ѣ�wF�E#�P��-Tb���𢫝p)	rD��
^�P�V8��x���1X�;v���X�T8�w�k�C͏ �����E_V	}�)}j*;|<!, RH�C�-h�Z:te��R<$�E�7��C�h�G�o�x*
�g�{ů�=<�;�y��{�   �s,�    l[�g:]m��.��.|��O[עd &�$�1�ڢ�ڣ*~tw�F4v~4���P??
��|Z�����G�9j~�Lj����L�eT�&�DEM�caмp�_�K�@�	���&��"�@���-���m�;	�a-��d9�w�k���й>�R�!.Z K�QK鹎��^�-xx/��d/*߹��h�op�;���x��x*X���U������Ū)Ct�9�����%���{��GCÓ]<O�@�V<�t�{>-h�Z:z��"�f��S5Q14B�EC�+�n�ra���<K�P�t>��-h�Z:z��1�Z�R�}��      I.剰    �t�WD�H��M2X��wl�R�J]t��I�����
:��G�&�}��~�0^��,��R<�ۅ��h�y~}����/)7���s�ϯ�qkKiRJ�G��i=0�V./a`�s�Sk��i�T`��h��V>Ͻb@ �i���������ޛ�/#�Q�tv�kG'馄ݴ$�! �$G�|Ã곜��[F�|�o�:M���@�\Na/EC�m����U�.cԢ����!-�b	���਱M��mxx/��@�Ut�h�k�뉃q�5
�%�*��ToMb��|�֠_s����	�d�UUE��GB�7��V=�.��-h�Z:z�釂��q[�Z<=>g��Y���   :��0    �Ni,'+Xu���vi�����-0 )�,r6%�(��L�T�f�*�]3}��2�x)+�n�r-�S�OTb�_b���I'Հ�%��!�)���~�*z����L9bgz]�[]���Y��*�s��R�	��$��𻮕ͽ�\��މ,�-[�������mpL�`��	d��k��][Y����w]+����we+�o4���j!L�n��V�����am��Kν��}x{��#�3     KVɰ    �7FN�����4�6�u�`���L���|?{�J�p��J�o��.��h7j�cƳk�d &�$�1�_��5����z��򺶷��վ�W6�+k�d�l�3#Nz>=����;��c�٩t�wWdI�����z
BX �%�@*�)��WV���\���\�G֍�|�������	�h��A^>���O*�{ޗumv�(̼6jk�տ��/�pMڭ�� :#Q�c�:�f��<7]s��m�                    n�n�}m|�8����tĘ                       �ͦ�v��u�;8����ʹ�]ִ���k1�n�4��4]�msV�B��YfӳI�����k�e7-H��4�k�+�Ǟu��y�wϞ���װ   -�ؖl    �M��0�l�M���q�h���-�b��}�]+���y���v��d ��fW�HK �[h]յ�\�GYY"ܮVU�����">���[��}o��[3�3����	�d��A[���˱e-��>��\֤��w[��\��a��Ā ����>�.��n-��7Εͽ�\�����lHbȍ=�{��k��T�N���*���������SET��6�i=O���9��J�8λf��A�t���;�9�5�u���b5jQ�"�s�9�A�A�A�A�W0Ny�z�A�A|5��i?���`�S��UUUUUUT ���z�    X���^����RNդgW@J\�,�ם�|O<�BED�8�y�A�Y/uox���aQS�b � � ����A�A�A�P�Dc|sV�'��i=N�����"�j���S{U�{�F�D�@��dKD��0�����A��h��y�fumuoy�faQL�ou30G�1�fw8�"�#�]�x&A�%�L}�/�>�:�7�5�q�aQ1Q����6��b9D5@ȃ��\��� � � �j � ���3;�9�wy�<��<���}}����	�Q�P;(E5�:�������B�uj �穄D9��;�8���J���D5ou4��$b��:�8�\�XA�A�K�MDD�u{�^���{ފ��Q56�^�������[y'�ك�W7�=�e�������      �V�:    ]�sm#h�I���v�Ġ`
BXCd)�`���qb�ma�7W���^U����վ��
BX ����
��wuҳ��n�_��g��b���^Ud��\��'6�&A�bZ"I9X�y�_�}���ȏ�z"�+f`�S �m��*�m"�0ݪ�JT���ő)$8lp�/�6Ub���IɬM7.Ӷ��'�x���ݖb���WUD�`5��db�y�>���Ŏ�s�+wd�oNE]}�	�]��Y���HK ��hW�������W���m��t��o+��X����`      y�K&�   �hg�[�h��Ր�d &%�&	i�菡<�����5��;�y==q}y��[�Y_��< ��lm�bɷ�z�M��km��f1^^��Z��Ӻo/�p)	`�Km1�ښ}qk�'��.�/�G�J��{��Y��՞/,&A�bY*`�X�	�\�oMյ��n����Uo6��H  Q-01]]ݖ�w�Z�m��s�'e���ny�    ٸ��    �Iz��<e���T���A)p��n��E��.�o���쌬kޯ+�����M���	�l ����c��}վS���\��[���麷����D�6 )jXH�;/ur�����_>�]"���}]��v��b�������r�M�`��\{��]���}=��=��=����ꍕ+��EC��f^{���ba� p;;�)\ݣ5�#;�r��c�9��gW��=>��TC�MJ�I$�X!J ��UH�>ߑ(�QD��_;d W�[E5&Q#D�=b堆?TJ"�"�B ����C�lR��P-�!"�T�{R$���1� "� P��%�J�	g�v!�Ǵs�Zs@U��;�{�  *�C��	ͳ~�Ҿ���~'�����_��;��z��|E�Į9=t`�&�~G�s��PǛc<O[	s�J��%�G�'/������>�}�~��A�QO���h!�,e��������K-'�8�[6�8=@����QG���U����=��|A���_�B�7D3��4�
#hy���>��T^����B֭�ǯ!�z?dY7�{���������x� V��Z��o�tBD@E$P% 5  $Q@�	$dD�	�A�dB@dBBD��FDF@I 	�d	���$d Z6"��-�ҁ�҈�?����֨{�Vϟk����p|{��P�D;U(H�"��(F(H�'�׿��|������A��q����^����\X}��}_Q�A�;(�#z;�g�W���~g�%v�1�\��_�}��g���<���� {���}���l��/�~��"�p� tר�}C'����6�ڐ��@=]¨���D��~�byL~��K�ߘ-�0[���6,�abŊ�o��q2 (�?q����rpxY\&L����pZ�UT?=�(ɭW�@�����B_�`6~� ���`�2 ���D��=j����x/���)���������şB\^��Fz�Q;�Y��Ox|��@�������=�-��"��Q������~���">�?e���~���8�w��{ܞ��>��;������QE�
)�b}���0>T������:�@Պ��l�,rM���#��J�ɷ>����X�q��������M�6���\|��>�~V�X�
3�ܿ��}'y�
���P��x��Q�\?���!�U#�`~%+��?�.�p�!C ��