BZh91AY&SYF|�]_�pp����� ����a�?      ������K]���Ǡ��U�3wa�UJ�6��jR�خ�T�Æ�jP���҃@��Ҵp��           �A@(          � �        ��  8     w��)UI�.}+�O^��:�+eY�]J:f���7jx��}fU�뽞����۾��n�������5E��4�HP �vV�pe�h���	v���l <��=w�M��P�����@JP�hY�����
P*�(Q�K�{���z[ս�\=;�{]vm��uUv������Tk����l<��x�Ǹ�<�o^�� �-�eհ � R%*� X���szYޠ�ޭU[sq�;u�`�ү{nһ�T�m��nҷR[Y��z�����F��ݶ���� )X��������W]��U�)uv����5�Ij�m���Y���.�����W]=x�p  ��T T+��nH��='���ށ�v�^��4p/{G���p��{��ݫ�z��\t��Pk^@� �J�Ǫ��^�漵��oP���pk]����x�^�k���r���P3/u.���  <zH�IIV=�ղ���Mo{�o���e{d)�ݩwP{�I�y7T��euMv��4��R�/d]y� {��QB���
^����Ζý�g�h�ʚ�z�{S:�7��6w\v�u�z�{X�=PP/��� 1�v����[��`myM��]髪W��Ow�]�[�؛�δ��{zs�N��^z����{��      (��JR"6����@�2 T��J�M0       ��5TTȚ�      S�ґ
J�i��h`�� *�E6U)R�0&� �` !H@���m@��ji� m&�d���LQ��a�����?����n��p׾���U�����*���N* ��������QU]!�����?�k�����TUV?�ʷ�TUW����?�E^��_���?�*���TNH4*�!A?�Q�����'!T9 ��U@�ry(-"	�NH�rDC����T�'%T9 ��Dȇ%A2P���䀧!9 ��A
� ���
'%9 )�EJ
r�*��
Р��䈧%P9")�@"rS��@"rP���P���$NH�9j ��CR%yr ��C�,�9 r@䡸^J��!���R�9 r �!�^B�9 r 仔�H�9rG�� @�9�9 rWR%yr ��C��,�9+�C�&�@��9 rP�r�J��)�C�!J�9�y
d�!NJ�9(r^H�%J�9(rW�'%N�y+�P�!H�9 r �����$J� ����%yrC�$yr ��^B���9)B�9�C��$y�C�:����ԁ�ܨ"!�AMH�rDS��D䊇$9"�S%�'$A9 ��QBrS�����'%9 &H�PNJ�rp���"�!9�;���w|l���������j ֯��F���������Rft���mf�tj{�˚�V�޸sXh��΋z{�w���wa��J��\��BfHZ0tuI�P���{η�o9�:��~[�5h׻��yч��ݧit�8�$�02t�7��tr\2G��ӽj����2L5��/�kÐ�^��C��v� ����3z�5��5�m��ph�!(K��n��B�8=�N�pru���iݏ��6ը�h���:v������:�o*el��L���y������A`��l�5ֻ;�Ay`k}u�i��İ�!��a��Y�>��<{�Ϟn�C��r1����q�q�K�=��#4ga��{�{��>�]&��n��J�N�������*@�m�7u��ܛt���c�׉�t�깅����q,e���A���f��yQ�R&С���S8�n���'�VdԔ��|ߞ�޺���sAx��n1��ٯ:so}����8:��7	BR��	I����Ij�z�A-N��#S��.�;=�}c��z��x�<��NRD{qt����~��<��H��鎛�f׿&��w�Xu��C�1��f���Ȉ<�:ǩ�C�$������>��;�>r�zv5�j}IC2��V�t�8��4��c��u�䱻u�Od�{ׇ���s��������6dsZ�٭��4mrLLÔ�di#!:�������h7��]��]%$�	�Y���c8�~w��k>��{�d	>3�	|�7
�I-t{�&�Ӹ3}y����}��+7��#�܄���Q*[آ�@��d��˒���~vvڴj5��Y����儞�x}����k\��'�ʪN����-l`Γ�%��H��O���oݎ�L�7�޻�z��˽�8D���{�4sGpa���|6���t�Տ��R�Ƚ�ȫ^�<S�#΃c����X����I��y컅8�B�0~���g�AB^O	�䥇dC^���LN]�>Ih��ҕDuԲ|�WA/i�U´��b�{j��,1(����)��s+" f!��7��dx���:�'agG��yގ2]r�N���;�mz����g9ֺ﮺=�u&�5	짱��7��r8�5�3���b� ���9�g�rQs�b���Ms�ٶ{���o���og#4q,�w!�C�]�=����K4m��q�O��=�у�y��oF[N	t�=��;Н�o�ug��P��u��N��;�tg�������;�8�7���A�=�s7��aN����ֶ��A�\�ތ�u�ߜ��7;�nQ�]�y߸:vo4k��*Ѡ:�hNN��e��4����[�O>�e�"m�'�2u��3��0��&g��E)f�Ɋ+d �c�X2��M)�naL��`�3��G�D���|y��j�Z7v9����-]i@�M4�G/
�����QZV�mM���OR�	��B�g�ݴ/!�595�ߍ�{n������:����ޯQ���T�y�x�L	��T=/�8(���+N*ay
!B�H��Oxӫ(X&����V���)��)/,�����c�Y��ΰ�O�o[8t݃��=�v�V&O2����҆���W� y�UU]�'B"ZЕ�!�i2y��[a�}��={ͦ�y�����󮍎�Ѥ�p��Fnw�{+�9�ú�Z��B���Q�â�ah'$�
4%)�BnS$)MJR��2s4�c��G��W^�٩��d��y�8u���V����asB<�7�7���Ws�,�z����}���w���Aâ��ӕ�<,B=��&�z�JQi8!C�r-��9�nN�4Y��Kk��va����d�iVNSS�ҝJ=D	Ɔ�w���g��k\PA�Bi��ڔ�:V�����f��yy0	����w�|ǩy�u����Z8�gG��yyo��|�V0�;'��m���%�l�D9��yjCp���c�ǒp��rCP�<t5���)�S*�]�*U�<��I�%���W�o7W�OI�Դ,X��y�L��zĻ�9Z�c�O�ft�&�4���!4	�˽Xy>�.|�BL���M��0�m��t����;���ͶAb��,�����fB8[ ����V6���r�'�³��p,�%�1��;��HI&kV�������Q��g�|Q�7�fb����{�
UTCQ54Py�L���Ue7�U	�R���Aa�V�F�����Xa���6f�����Y��9�u�n\�H��:�N�=��)!)N�<��)
��2V�<��{�v�p�#w�������/?o��z{�&����Pc���1�D�3|�Q�x�$�$�f[��	�IJb}ARɁ���}9����Z:��ëƺT����O�wE�@�ԥd5/b�ׁÑ��F��`h�n[���3��;[N@��=�ӛ/L�*J]B�X��&��1
SN÷'��+])��m�V�����Y���0�i���N(	Ęo=�	.�$�%�!�M�r2"�a�'s��G�f�vss�s
i��[B�bG���c�*=��$Ѿty�oέ��Of��:`��1�8k0��^h�K5���x��a�ĥ<|zu���wwp՜�OK��
�	'��������^��$}^M���{�1y	a%�y�̲o���a�����NBRB����X޲O���Jԙ��h̹Iт�il�I�띖���p�-OG|�w���"$Iё.�0�<�Ɇy���*���ԅ~����R���K���)L�>mVR�,�XZi�2i`L&$�����{�5�_�R��ȁby�ޓ(��p��==��f���ɯ4VdX%�gv�G8��'r���(M�P���A���Y��{<fy���$���>�����*2���*�_��5�� �a&F������gq�o�}8��c��津���s}ke)Be6�F%)tka��G���D��w���z��f�]s�*9߼�is�5��ߜ�PkQ�>*�M8P���-m��F��Xيӆ��i���9�|�#��[�uֺ;,�\�4mٝ���n�֞��ko9��;NkgWwu�촘�3S�y�Y:!�PF}��9�p���
����[���9�u�04hU�8p�5ٽs�y�� ����i��r]]`��ϳ|
� ��WJ�u�����{����z�|��{^%c�9[8�Sꡬ���T��Ǔy2d���7�*�#�=&�C6A���~���9�}������F�rt��e�ۨ1Ӣqׁ�'� �p�5�;�+V�QJ��zyR�ޕOn�b�HC���:�vy���o��z�t�3��9��%Ӵ���X��8�$ϨAw��I�K]��զ��P���Ld���hI��y;��L!X�MA��t9�kg<��Z��'v����2vj�[�hk3̐����B�C�MV��MJt�~gN��X:yq�5U*qH�Z����kN�1������ód�`W�7����)��%&&BP�gDtN\�h:�<:�FQnݽ���w�o֠�
����O���v��<|{�u��=��}�u��7�]l킌g;:�-��v�r�h�}wu�Z�=�{��ֵ�K��'q�[�	��Lc{�G���=�/�k���|�fλsf�%�baUZ|z��P�e
j�;��2xly�����ϊU�u��k��߷Dg�p��;��
�$�L��Y��#�ǋ��"���x�j��o���^OG�Pc�`�;�3b
�,E��s{M'����'H] w1+�n�w�+�:Pz^[��w��sĈ����|��	�^B[O���}�Gr�m7��sg��F�<<7OCS����S������ǳG��/M�:��o�/o����7����t�������4Y��h�뽝w�ggq��}�â��9뙦��5�?���X�%���S@L� ;��Rzf �;;�o]�+T��xi��<\�"L��3<JO�(�l�e�3ħeuJ!E��F��T�:y���;�u��qӳuǣ}�:"��k�No��o�4l5���j|�z�Gi��d^硬۹�:��������� pi���Z<�"5��ӬL��0'��0��]ߙg�֝C�e��SX��^E��K���h�9L�1��xE����nX��S{�3�}wU�y#�d)X�ڦ�홋X��'�v�wL�X��]B�4/7�rJPvm�F��=���V\�޴vgv���u���^�v��]�j��@��]m�}�s�xs��ᆶp�3�����/g�Ē޷��oc�κ�5��ׁc�~u���{J�Ԋ�c�Ow)Ƶ�OWoo^�U^�7�s���]�ky.��p<�E�0܅`h�݆�mc�P�����6�}��o0�F���k�(J��%)�O!:��(NJw/�!�n�'���Q�%]*ɴy��]x�^}����# ��9A�WF��.9h7ֺ��]txt��3{��=�9�&Q��F�5���x�]�$c�J���O���{�Z�x'��o�;<v���[��N�V��\�sh'P��3V���!F8���1#!(u��u�����:κ�������ad�5�vA��o7	t�A��cdb�	Ha���gVIR��V$��6�V��;+^y��=g]h����\��n��k�����|����𞄲PR���J4��>[�gGpjWNC�&�;�~�<p���:)\zU&����ޭQb�-����)�L7��0����$����s�6sz�G�l��4v�w�`ݛ28u��j�5�!�N�0C<����'ą"jY�E�oG5�7��4`]��y��qq�D��ı�����F�NÛv:ͤ��lĳgD朘��u��`h5&:M�Ln6�=u���Ov����s��4�6p��5�,�X^��������	�BrR��M�u!�&@�&I�kíA٧X�ѷ���a;���ѹ4�l��jA�^y��d�2�яM�i�)17$՜�::6w��;x�bh;�Z��)�0� �F�N��l�Q��:�K+7��8�(;��ĤS��(/Dc��fͼxk<���Y�@f�vh�gFk��+�E�f�8a�w�:�aȑ$��O�4l���õ�{&<�ëXպ\���VNO'4p<��c���{�㭎��3��W���}np�|w���f�4y�>�#��0�&&v����IE�Zt�;��R!�
3���-�n��Vuc�����^�I�«�&�ݝD���G���j�J�������|_�-%
�츼�!˽VUjӋbM��B�$7�OlǕ�h�g��!�����s����|�9֣t�C�Z�d�E�D�z%�_��T*�V:!(�a3ͺ�TŚ�G�h���7��&�-:��F�oYѣn�8�!3��XG��'%_���ԗx�<��,��3a�̮��R���{ػM�2����L]:Y�N'P����m�����oi�����wu��]ݨ�I��J�kh[r+"���}�p�)��S~�������x|�H��õ�d����B}+�A$��Rp�+�JN�e�)�~�󞐬��	��v	��9n��|�ww�-�xd�(K��<t>nB�ô��6冴쵎o���KD����&<	9)����������|�d�r�\�ժ����VSz�����>,dٵJ7kF�-��-�b�nC���W/����]�q?No }�[$m[�4�-ˋS���$��"aY�z[����>�}��4��oo~ϥ)�q���� ����F��{�u$]����{��S)�wL��w.=�S)��e2��S)��e2�L�S)��e2��d��w.fS)��e2��~3���������q_�:ں��i��2�L�S)��e2�L�X�ڸ��)��e2�[Owu��L�S)��e2�M�2�L�S)��e2�L�S)�r��g.�ǟf�]���)Q�	{���)�˪�e2�L�S)��e2�L�����m=�S)��e2�L�S)�gfr�=�S)��e2��e:?��)��g�?L�S)��e2�L�����Oq��S)��e2�L�S)��L�:��L�e�L���&SR�L�z�L��$���)��hv�e2��e0��˸�Je2�*��f�*x�FS)��e2�Jք���I�g-�j��W�Cw��RfH`�}�s�㯨K�����k�H�s���� �2��y��wq�4;�{��P�����47����b�k�8��O��Cs�Ԥ vb�Q�;��	����I��ʩ�mRs����j0�$��ռ/Q(���:�oX3�n��w�q�����W��X�8���ywI����y�z�? 4�`���|�D��]zs�[�HS����.eԏ>�ؓ����f<�y�Y9)�t�"��0y���ҳ�D�-��݅����d�{��!�Gd��`\.��{C�ePzjx����Qn#�Ĕu�ʚ���e�� �|�{N�,�������/ϋ 
L������s������!�]�r�x���^�Jw��r 8�b���C8�e2�L�S)��e2�L��e2�L�S)��e2�L�S)��e2�L�S)��e2�L�S)��e2�L�S)��f����wt�L�S)��e2�L�S)��e2�L�S)��e2�L�S)���{�����e2�L�S)��e2�L�S)��e2�L���)��e2�L 
e2�L�S)���m=����e2�L�S)��e2�L�S)��e2�L�S)��e2�L2d2�L��e2�L�^�i��)��e2�L�S)��e2�L�S)��e2�L�S)�ɓ�$��'�[�y�8��#AEn���Q���LJ4\GxU�k��dnO�� ��ܘ��s*r���vv'�e��$�@�p^��LR��iMe��cޯ6�Ȧ�L�/j��}"s�Фc�C�}�B�,�N�����9A��	!C�Ot��������S�ȇԗ�Y��3�b@ﱺ LJ^�l����KU)��`���]� 7��m��\�n�q���T��6�O9j���rĒ$�x�%%$��5�àju��voq]���L�{BP�t�[�nsH=gt��Ù�������s�fR�$��ww�2If�A5���d���#.�q���/o���+|Im.�	���p�2��S����e�L>k�õ-��C�R�E�ͅ�X� � H���	.���� �e�O>�f  /_D������Ws���{B�t[����0^s~Nc�&�*| ��.���'sq���k� ��x�x��R2�^9�Y @v�����nq��g�
m2mCy���陫�n������d�˘��+2�k�y���^DXK\��}U���Z�o�����n�� �a���`n><8��I/����m�:��5c�w}��sds0�ܺx%�i�RA4��{��k�J�±1ޗ��R���:��8��N���I�g-gN�Pr�e3��YNg{R:��@��<�� ���q����V�v�]y}9y��3��׆M��{��F/k�-ޚd��������s%>�4���܉ M��Jsg�����T����{윐�)���R|S5��cc��v+�h�qܗtt}LY1"�M$��:�9zJ�G�r��l�k�6t���
�I`d5/Km=�xi����<H	KҺ��V�K��s0��`�y��s<�4E���J{���!��e�З��add�3�6����bqS�wm�V
F�����E�TM�)�G�f�q�<&`#۩f�Bp�h�G¸E��]��{����aFh���by�۝���Ǽ�wf	"跩~��7�]؎��˃.;@�2�Vi�&K�{h����aRr]ܕ�
�6n�0�>����Z����E;�էZc9l-�����y7H���;�j���2��>
`6�x	�I�����E����/a����6�g'�Q�c��ȷ)�'���yY�.y��>��]��ˎ&"_v��npKx���Bw�̎;��=�f��;[���9�?6����^�/#��#��H���8K:cIu6�р{���3x�oiꬃ��.##�sy��nI���Xɰ�f��F��2ܩ�ݶ�~�v]���n|�W��{1r��wq�K��S��^�x�f���(��A q�R��8�cݨ�"��e�d���}�q�ݤ��Y���N��$�yY��c����7��CRsFN���Q�6Fŷ��Z��L�!����]֯����1-�Y3�
wB)�s��h����\	�I�jGoE�7�,�G4IJ�Y�>�%��ߝf�����崫���w�0փUq�<P�^ggg���޼�Hxg@�0���3�ǹ���p*5�yvd��zp�4�6j���yP=g��h��}�t=��=���g��K� �+�M���1� ��J��y�qN~zM4݅��nV�y.l��"�� 8WOh�F�o��{��d�8���{������Gݥ�\M�s<�g�vp飦����Y���u�Ү�!�>^�|?#�G�{g&�g�y�������W�s���	X8`�M,/k��y���MԮ��$>~D{{���[m���=��7�\�XY"�6u�RH��(a�º�]��7ŲD�)�8I J���<����گM��jNq%�U9f{d��k8T��1��(a��:K�ju�#С�\�|V��	����B�$�Gwu%�wzA{F��c������D�ߦ�d1�#�s���:�f�F�]����c��%Ƈ:�O')��n;kl�٘�y���7w�� x�O���Oy���y,��7ړ�� ᓺ$�n��u`p
=ik�C�M���@T	='���gGj�oA�=��j<W�)�ՠ~����3���zS�0-�R`��=c�K;�SC��G���A��"f`�u������UOx 8�h2.;��C<<'��@o�=��7��q|�h�]�wf^n�K!2����淹�Ny7����A��X�������]���y�rdeM�!p�u���wc��>�~,f::�|�}�}ɦS��-7�q�]�|I�%�;D%u=�S)��I׾WǾ\6���ԝU*G_�*��3ğ�b�I$�o�M���~mT�Cs֐-㳱�^�  px�(��x��ڭ~.�#,�ĻP��װ�O�z楬W1$�2�=���7ys�֢d0�VI6N��fd���a!P[0>���L�u؏�����+1��ZWv� g��u�㠰b9n�շz٬i�B��$�g��۩4��`׼t�C7�&�b��=vR��;Z=�Խ���>v^��i�J�<s�<�i�vB��2�I2�L����]5Β���<�q��H�P�a���wd2�L�S)��c��ׅ�j�ȭȰ��tn�G��i[����+����pʡ^Đ���3�
�M��]5���e2�L�S)��e2�N�)pe��-�&�wR����2w�C�v(�oGF:���;B�_$ŧ���zBO%��鵶tbb}9ow�^Y�5��P��$��~��s��6kX#�+�q���q�2�]�,?��s�4x�&�|�I�EԞk�%�Nt<��{��[�U=�֎>ś���1����\{�̧�������g�t���4	#w͞�����I��C/����c��vS�Gc�t)9�d�J˛�Wr�x����{��KR�e�fw:��2���#��N��a*k�=oj  ��� 
�g��SI��n�C�D�&�@<ݢ���;�].�n�W���w[�%sݼ�Ywwvs����l4�z��xOD�%����� )�;��L��,�qm[z(s_��Rӝ+��)�˅����i]u�π���}��G@���Т�E;w��+��@�i��t�����[#Z�"�uJ��+���ݣ� )���;h��t��ޠi�n��4N�4g(�㫦�7v�S)�^ �������$�rJG�ߘiqx���=ǥ� ��I)"@�hA�+��_�����p����mXO"`
�L����6k�bS�?���k��P�Jb=Ox�ZGnz��EG��m$�I�w�3 ��	�o%N5��(�7�3�;�l�2�w	�wr�\�� _bj�<]K^���[&#)�m6+��>e��L�D˛Gn���S�xnގ���%7^���yâ�-&���^5ww�]�p�.��H�L)�9��`(�י���'H��f�N��₄�/L��cȍ[�QT��!�1ۄ2To�S:�Iԇ�0��Ȓ���gv�=��b��I�2 C�(I��$	$�Wf������w���{�uMi�{#H�������60zv���ܣV_q�G�Ê�0��ɭ�/&L^@�)�f�uI��~��Y�4�pT3����)gc�wE*c ��?tr�@��8�ڷ3��a�06��gnT�t�]�B<B��&��C␽aׯ�v��Y����7��	 :��B�������%�+�0��~/#d�Z}c��ב	��<ٻ�E��<l&qXF�Y#�%����hG�f�����YM�#VB<[�^��㛀C��2���xG��w�������7�0"ٽdl�Ξ�I��SMd��;�\�v�7=;������+�!���a�n�6"9����	&����B��̨�2|[��	���2�u�`jƪ�>m�B�o�h�xz��)˱<�{���|6�ߠ�s̙���,�+�=�[^�b��D�>E���Ö�1#!��38��_$D�� K{(k��H�����|I�v��#�:�^��=�u��Ϗ"8�~�l��0�噇�cs0 ��@>��MG;����O@��+G����S7e��<ɲ�
�� nu͖mOs�����	�E<��;�A\k/�s4������bS}"F)��/�pI	�$�}P��-:%I!����dw63���^�AʭĐ>8��놾�[�e1��]Գ�&�K��d���Ũ�2s�M/쳶`�{�a�����@Y�/e�&��o�3������/�a��%�����ӽ��y�Y��P֙��M���n���z�=	�ٻ��E�N׉�w4VMI�;�ː��Ʉ�j��q���/n̫��<��<Ll��j$x%3n�U��R�/�ȮHcՃ5��%#���m��4Y�||tM3LpH�Gݣ�(�y���s��T�ި���I5!�|�;�^��.��5��V�d�XQ��l+����-؂��f�*рy�{���Y�"7&�P�{����7G�"sr�y)`gP|!�%���7�s��t\���'�X�rǄ�BI~>��o�w��]+��g�)�3	��/�U��!+�{�^�@�_����8!��7w�����)���zA$�߷��ɂh����-���jD��é��g�����|;ͮ*,N���9n��e2�q.��q���)��uۻ��L��i28� �O��lZ%�7m��T�9%Jd.'{��n��H<�J��'�y(e1��IOq�����I���M����e�ܺk�E�a���_��gf�&��2F���O�8�I;��ĝm�<��Oa�+x�ʕq����z��)�С��mi���e�3OC)�]f����t����?
�)�wt�aw��n������W�������@�� $$� ��z ��%\Pstz1����y���ҋw�1�ܐ��IN�E�Kzߊa��w2���E�v��u=�S)��}F�7u������ZK�����Ŷ��Ru�Cl?4�2za�N�΋$Ixf �rH�����aKOIǉt�e2���J8�p���)�� io[~x�.=sn�Vap��,��NAo���v<�u�����w}�k�o2��ξ2d7��@��\S[���*�i2WK/!\{��SR&Q�d���p���ΛL�a~za[�,{�l<N2��V�|n1��D��6���/��!��wv�1�m�y� +Y$�$�p�lę����f���{��S���frr+p��=v��l.i.��$2��;@|f<�b���/o�>&����Eᅑ�8y�f�K�x��w�s=�q��f]�w�(�˽-Isp�Cm�DhQ��{s�F��d�� ��y'Q)t;����(1���ElG�O�X�70�<�q�G��S� ��2�K��w�1�7p}��8}���Iҝխ�Ƿ�"˦��J��g=<��ή5��'��&S�4P�aU�R:*�+UC���G������0T�:k �x��jv�RhږnhMo��G�)-�27ǪP����������\�r\줝�w��N$\.�oʹ��$���������*���Fd�v���ŌAGvc : ��E3�3j\�$�3	=�2,m���x��{��z쓤��W @�ꩾ��M��L.ޒ-60 ����U���ݻ`˱~[u�˦9���]�/t�'��+� �yδ���L�\D��2�L�S)���>�XO;��t��#��9@o��ڂ��c���|I)B6�[)=��i>w9�����-'��d5��(��jуZ����J����n��a�&�ha�s������<ǩ-�@�w��J=G�RD�J�r�z6䤣�鹻���;�ŵfn�j� �(m�"Q'�[�7�xdZs�G2��c,j�u�򇬀^F�����\(]�_x�S�.7pn��x������C��w��I`�$"��hz)��y��?��� �����Ш ����v���������=�?�?�?����?��"��&��?�C��E��v�� �)�( !	؈��x�W���\;Dt�z��h$I)a� !"	���&��fR�� &�@��d�J�$�*`�$���� � XiB �e��$h! � ���H��$��j�����"�@�N�@�N�S�%OADЉ�T.@���L�@U
A@3�0�IA10ň��B��ID��- � �T�
�����;]�z���� &��ک��(�"�Bxt�t�������LD;P ����S�E}H@�Q����"�*J�zU��S�ʈH��Oq;;�LK�JDҫ҂v�t��1q0���"D� = �*�AE(U2B�HJ��)B1!BB@� J4�.ٙR�0 e膄�v�pU�<��C4Rv(� <U >�� �  ��b�L�x�*8"�(v�%|; � ��D�P��;Ы���h*�
mP�����U���?�?������Ӎ��������uJK�H�
2�J�2A2�I
�P�BR���2P�%	BQ%R�)HP���%	JR%)HP�� )T�J�("�$ � �A�����]��������N�γ3-�s�V��y�q����yҧ~���~�R%t��!T�*�6w��W>�pp�k��hW^����.�n��U\AP*E�����[u۝���U�3��m۱���su[�Df-XLJUh�B��g:<It��]ְ���W
��a���r��b�K��:�n��v^Z*��> 3gL��O<.±ݡs�Ca���&i�ڊ����3D�svs���[l��b�85C{:h��X���Ɨn��:�X��K1,v���B��p<�Y�m����ݝ��Ա��SU�D�[t͗k��n�ҙݮ�H'��8���1	���W@��f��rn�tß���m�1�i��+���7�%d�ɈI��Pm���1mģQ�ĵ�c�4�Xl\���L��~TE��E�C�E{%_��@�#�y�\�~���_��0rfd6kO6��٭�}�Z���<-㳵�^�mv�rVJh���#���!�,-ݗ#��Ϋz�3E�"�U�����^^pժt:?�I��0��jߗ��^����W��Ҋ�4u���r!ƥ��#I �m�p�u�.�H^g��Q4��V�������ｷV/����{h�E}�_�I�s2X�,�)5���cM�p���@*�v\��Z�r5v���Gl>ݚX��=��y�yNn�m�[��:Q!��i�2����|���ｷ]���>q5;��G��\���I�E�D�E6�M˰7�{h>�v��������^�><{M*p��K��l�r����y ���(s/7�{l>ݚ{�6�Y[�H�	�ҵV�3�<L��l�����L�g?K�tՇ�x����Z�i5rJ�_�g��۲���l3]n�7�4�S�uw$ut�m���vXŖ`�Lm�T�W�V��%p)�[��N�'��O~a������l�۵
��6�N���6���D�����H"h��{۷V���������J�F|�W�[P�w�i+�+5��͇6X�ؐ�ݗ�Yz��Ԧ�c���������}�m%YK�^O�yC�d�-�ZC��D;�&wS/23��ʘ;�y$׻+��[v����m��饇�+�$m2�9c.@[�~_�z����&��,R��u�й�&�m��hB�&����/{]�o�v�Xyj�oT]۾����0�M1��`M]�,D4���� U�,�e��3^C--�C$e��]��*;�϶i`��v����a�zia��zڎ1�n�M�Z��m�e�/6T���&mm�y1��F}�1딘�;�P�Q"�b���n�e¯cK�1//M¦v� �xd�*�S!tX�m��ݠ��uZ��+f&�XRZ5�K#�4�'�yr�;b�g]wjR��F�+��D�3�D����{[WEn�5�F�`���2<�����M�6�ӣ]�6L�۟d�9�)tcD��6)�$�A����و��t$�-�����]�������&'}��4�.�i����'��*�l�&~E'���������zV�+��l)";��+�@d�1[�,�4�@��ᶃ>�[h1{��׺�=�y�=�B�v�����
7V����/���h�-OD�*�A+-�Ձ���X1�e���Z@��[,Y����*2�YV�P��uX��,}綀���j����V\�q�X_O�z�	���h�	u ��Km�i��!�	�(nBP����[��X1�e�b�����&i�gc[�l]H؅��&�!�v)Z����rp4q{��Z��L{)��������0����c����,[7)WM�9$�'#רv���m&�G#��]�BpMP`n��A�Ƕ�f��`Vo��{ߵ�DӦ�w��w!�K{���^C�����߷e��W��lHQ�j�:��E����@��ג�2�vٲ�^2ׄ�9"�r��RH��J�@{�{h��,����W���V��h��ý�~f��y`<V̉3&�O[t\�W��%
���~?��%�4�>_{]�|�7���Wϕh��� r�Z/[�D�x����l3_�Y�-���`{����]�6�~�yv�D�n���������I�`�X��I`ⅎCF(D�Df`�a�3�X@D!iR@H������j����`g�+m=�f��Z�i��n�l�,�}��������G�C,�7i�Ԕ�\$m�$l{h<��v���D��vٞ�P��(ڴخ��Cv!�ϛ��:��2֥���K+Jm�fn�:R%s������(u�e³#I���/�8�췬�d����&Ω5��?+a��v�g�4���m�ګm���H�r���H8��>^�N��n˅�F�fF�Lb��L�"��.�ǐ�
̍$��e�/$����:ݶ}�K��4L�I�i�L�5�l�Sf��[fˆ�����(6%W-�I�������)?4����M���,݋���9�:�
V���6dU��ۋp��M���ڎ�"ʎV�j;Dx���whP��a-�͟e��/y2��믷_&��r60�M��߷n��{�I-^ys������#��n��+�i��37n���%��������;�3��P�=�$7v���Ӆ�{��$�N�\��Qr��=NI��J��vQrb��4КY��k3]��Hs���[x�g[�+m���5m1ݸ���;���5�y�;tki9��й���zxB_2�q]��nn��᷎�s�����1���ܹ��^6rs��$��h�v�62w��L�����OO�lҼK�hT���DI��[�\���2�9�"o>{���ẫ}�۬��:)l���)ӐHt�T1R]�:Sf��]`O=�����.y�տN�w�׳(�p��Q�C����u����Ta�ʶ�ea���gqφ�#�f߶�Z�/����/�����=7o7�l��s��k[՜>Q��{�=��Ү�֕�%�|hظv��<At��}����v���e5���.:FՔ-^�8uͻV���sϯU�x\�[Nn <з���=��w���AF��!�v�*mn�s����wSZ�o~�>�㥩ps��wS��f�s�ڔ�8xwdcq�p��
�6��B��[9�79��۾lR�����T�<����FOǤ��|���z�קU�O^��;��a�u:�xvu{��K�i���{�ջ��L��tn�5i>Ax�%zN>vZ��{T37�u�mi����(ێ(���~��mݛһq�
n�eQ�kUٮ�ވ&ڝ�f��<������WV<��9�05������G�<<h���W����KW�=mäh�?�=���K���NG�L:��~�y��[:�9G�Gݻ�=H���ܖ(�7=徕䗔�ɝ�^�³wcg�\���#G�x�$�����|ݵy��\�\��|@ՠ!��f���Q�Rڼ��7m^�������4h�7E?��ۢB�)���H����I��Ű͢�-���S+��~|��)z�L�G��;��O��W�pn �d2JFi��̣�EE��|�h�36h/]h��vU��!DB�C���ǀM�4#q�[��*�N�K�q���w���I!�+�xe����@?����<:�M��l,������c��a�f:��|-h��Q7��I�Igy
�;��n��IÝ4Fs��[  �� �m�
@��6a�N�����JH�jL�/}���o��pV�٩�!$�sE���H���Y�u�"sYf:v��j20$��[�vSJ����'�w���k{��#	$�bxa�a޷�"�ĺ4��f둢y�\ޝob��;���3]8wh����<���
�2vMtoN6w���`�I��f��<z���;PS���4o6h9���ge���*)�s���z��y�^���$��$�C�f|y�n���9��ёl��at��dl�;�8�a8ak�I�ok�l�l'���Đf�4+�Ȝ�y+���.��g���&�1(�"J
ʓ9���o_����;��m4�L�\��U����*fU�/�3�ͬ�ʃ�0.c]	%ŮH��Mi��2.C8Zq�&�1�CIj��Ƀ":�*`ffff�ffd&f�Fʳ31���9��=��6��L� Km�2�ǘ ��{F��[j��ONјc-�1��(�e4uۉ2mr��v�:-	�L�M'ew2�.����.ֺW�uq�a2�8، D
�Zl�+ʳKs���k����Ax�]�k�&��D��D�H�6Mv��Ź�k$�Y��c/oGbH������q�2�^okFP�]����]�Y"�V���a�<�����[K2T]3G�;Rh�(���vs�$Ul+[��l�k��	�%��ۇn����\�n�R���E{nG,�;F.��]uK��6���]v"01�r�[r�ۖ������/����wb@�s��Ǚt7=E��-e��g���";�8;e��6�r���d���L�.Lj�4�j�-�:�(��؋SM�&}����(:X0�cYu�F�n����lN='s�mի���z:�&��[0��*�:�i:����ِ�D�Wa��{úp�1<�>�:;��\1O�M�Z3� �WDWeO7�MK�]���-kl��JGY�#��o96D��s�m��m����%e�nG��SZ�+
��+ڷ��Fe/��'@��*?�VP?�T4���(��>�
������ �D��H@�z�ԧ���Bd�'~y���)��=�fk_o0�淽뜵����)Cמh���)N��~��);��}�/P��-�}��)���߬�32��twk|�u��8o��	����P5�7�.�f��z�c�5�P��^��r����Z�מ����)O3�}���)I}����y�v9���f���@�2���vp073l��(i���	I��������Ϸ�� i:��}��n�)O3����	By���5��^�N��Q�U�vO	8	9=~~���N�(s�}��ԥ)���f	JG�n:�d���{5i�-3:yI3���;�7�(N��G�`�	Jw���)��I���I�	ߟl��d���~��,oy��O<���s{'�9��}�~ބ�i;��}��%)�y�}�rBC�L,Ԅ@Q$p�VtO�-�=(��]	�y��/kgt�7��v�C��6z��8wQ]�6�k���Jv:�E��z�y6$�ģ�su�ZU�-6&��ޱ�M+mqn�lxj��&��V�lm{m�,��1a�4f�K�LR,u͗��'E͚5���<*{�~���'Rw.G���y���n� 浭og5���(��_}�� IIޞw����J�n�RhP4ڥe�l��@SAf/|�ϟ�i8�ߺ}�z��{(zyݞ��{̶qu�ys��bh���H��t�A4�cWC��)�kX%)C�h��:����{�������Ͽ~��)O��}��y�k8����p��MJP�����:��<�߹�)#$��t}�R����~�5��{���f�=I�sG5�θsZ�����w����G�`u)Jy����	JP�ߺ���)��}>�������y��8�);��}�'P4'yﹿ�2��>�Iԥ*���e�K�����gw�G��:��S�ָ�BR�g���ԥ� 󭜏}��FjF`�M��Z�ao7�3v�-��Z�����߰~��=����L����4}�R��{���,ٮ�s� Jąu��:��l�I�n��bF��g ��u�v-�a�.nv��&�9��$l����v5ssc)�sa{g�hz.H��ܼ�"���k��C�PC�tk�+2�ek3Y�nKZX&UA���r9sￓ߰:�����^��j��<��`�&�����s�)�d��{}��Y�7�g��9ֹ͙\��JR�g�����O1ԥ'����z��=�o�pw�d���>��2�G�����޸���|��֮	���y����R����Z����~����)O3�^��j�<�>��N�p�Noy�GZ6}��=�R�g=��	�4?y��>��JS��ߵ�)~�$���Iԥ7��|Z����kv�sw7�k�n�����u4{	�9��NI��ؿ-����0Kܺl%ԥһF��%��9����?�S h>�����nC%;�=�ք�[��'s���*��tΥT��	��snsv�sM�T���r{}�u)I�~k�:��;��}��C˳�8^�y�x�tB!Ԥ��!��woy�R�������G�4�
2k�x*�M�}�����j����_��R���}�>�O��i�~�~��N���ԛ�Z9��}j�g�JS�����r(
��߸=JR��־�ԥ}�����R������l�ֹ�k��m�)K��!���~��J��}��	���y��N�hO}׷���}��In�aU2:VJ�m*��;��o��(�o��n�e�[�q�և�1�H5.��Xp��Y�q��5��?BR���}�iL���/o?��U~
�{xRJ�$cW����=��tQ2��=F��n���׿bu)Jw����	JP�����N�)Os�s�)�{{��k�#�Rs\�W[�l��J\��w��N�(}�`u)Jy�����u	�y��}�R��מƳ5���p浭l湽f�&JP��y��N�hN��︦��bF��@�Q|��3]h���)O=�_p�(N�=�3��y��:��殷�gN�=BW�Q��_���!)<�߷�N�hO}׶���O��d�����N�)�}��kY�oW ���n7�����'�y��:' I;<�'�j��U��5i����]\P�uF�ܹ{�}�}��5)C��}��J����`����߬o�����2��Ŗ\�J�59X��s��n���@�'�?~�ꔥ��~��C����������(<�/<oE	IB^�i�-ù�9���W��]��ߠ�?�!��{����)JO��_�`�	Jw�^��?���3����Y��ٙ��u[�ι�����uB{��_��)�;�^����2S�k�R����t~��ԤV騈UБK���)�y��L�����~��)J}����)JO���O	�?=�嵞�[XX,f�i<�.5��u;uN��a2�d6���Fn%j�
vf�bu�.����NJl]��\��*{vw;r-���tK,em*T�S"������o��X�W����Cku��/0e*���x�90�f�,լ���ofk[ٱs�������r�h�눇b�<�)�5C�JT{�=���?YȜ�	�;,�:-�n�=s�Jy9�g4ogG}��~��R��<��qJR��>���JS�y��z�f���7�s�����v�z�Km<pt�W;���{�J|��=JR�g��qM@�w����)N�׻�X�!�}�f���I��,�u��=BR����}�d%'���~��C��N��^��j��=׿bu'�	r}���ѳoQ�7�k|�淜R�����~�����w��h� ���߱:��>�m}�ԇ~�}����\:�|�[3{����p:��{�^��R����}���JR����}�d'�V2O����?��/�����[ֳ�Z��fs[ݭ�Sq�&I����O I_S��"X16Ѩ�M�2jP��LZ��g=����D�):��}�/P��~}�����{�F�J2�
�.;��f]�(�?6�x���rB��M.����ϳnCG`�@u��q��N�n=nBnNl����Ɔq�ͦcP�5)sK�s��$������ԔcV�j޻L��n����{k�`����u�؝JR���w��B���Ͻ���BSٞ����5��\޳z���9	I�}����>���&�({��}�ԥ)ߚ��┇��}�lޝ�ǩ9��֮��\5�R���}���%	�����؝JО痿qM@Ю��s%G���ڳ���#Ԓ���x�Z�����=���BR����}�d%'�y������>���&�=��h���Zx�&u�s]s��o�ԥ)ߚ�j�' G��[-U��F���g\�n6rU�MݤW���t{�'�4'����)@�{�}��R9���s��՝�w-���v�P�Ʊ�����{{ݶ^�@� r{����N�)N�׷�!)>��v��wBg�ow�&H}��ky��3z�ԛ�Z���f�'R��y��k�x~$�a�!�QH�0P(Y��Hg��q�(������JR�����Bd�'�}���p�>/�8���9�f[�\����4}�R�����z�);��}�P��y�~�5߾��|Zս�Rk���e�}n���hC�~���}�^��ԥ)�}�~ބ�
��G�bu	O�y�ַ���6p���٭Z��w	I��{���=��w�uݙ��a�˂D�Z64.��L�&Zu��k7�}��w�`��]��߰:��=�=�\R���ߋZ�5�é:|g����8�1%��y�zG5�f�n��R�g���ԥ'�{����S�~��r��<���O p�>}ef��2�^Ǯ�g s�}��~�����ԧ�����L������N�hO|�{�0�;<��>�{�ǩ7�j�[ֺw����<׿oBR��N��G�X�@tr�:U5�^J{�]}�u	I��}��:����{���Zޮ!��{�ke�w�@���4}�R��y��k�R�ԝ�=��>� ܂y�y��$>���oXo3�Rs{�U��vk[��)@��p�99'|'��'��6�m.�X��Ĭՙ&�jImt�e���99>~�G߰3�R��=��oBR��w���r=�}/�ֽ�uF��G��!v��6�과�9��s�����9	>��}��	߿ow�&@�y���N�)N��{����^��[�ћ��;�3:�\3E��R��<�>�JPy߾��:���O}�����({��}��"S���[,�2�pf���[���u	I�~h���hN��^��jE/0>��}��(�C�~���(N�|���k��ÓoW��'d�� NI?|m�~�5)I�k�z��;�>��	��f��!� �����l��!�L)�@��01%� 22 ' ����tn�F*T㶒�tm��l��f���9+�\�F�ۃ(�Q �Vc!t`�ˀe��.L�2N6��*�1�\�\0\���5�1�3�Ac��m͞���e�c�a��6]����3�1����jF�Tb��陶��c�D9'�}����)�>�s�Y�6p��7��Y�8%)C߾k�z��9�F���Ϯyk"5��z�n�Vff��lˊ�}�k߱MBR}ߺ��N�hN��߸��:�Ͼ7lٚ��xI^���ű���kZfnf�(%oU�p���ԥ)������)I��h��N�)N��︢����:�_�
��^]ˣ'*UW$Q˫W�	���w��>��@�d��}�)@��߾���)N��^��u���߫�_Vk5é9������7��JS��׿`�����4��R��g��Д�'��������/����j� ��\޳���n⛀�$��t}�'P4'y����{���'R��份�HK������;��ja4V��N�)O3�߸�n��/:�����ū��%B�u��u��ّ�͛����oNn�P�ϵ��O hO��_}�jR������I�9>:��}�v��7�=��z]��!���7�����1Ǜ�性ӝ���E7|�ރS�٬H$���l�h�&Y���f�0p ��FY�xC�{:��s��;{� ��Y,��3;�B���h�C��vՍI��sÁ۸�"�L�X�uC0��Yֻ����}o\9ջ��4���Q�Ţ2�Z�f��`��P4o���G���"g���9���fK<�v�� Hci�m�bh��� h"��gq�5�ދ��3%$�F�XkM�֛7�I�	��;��f�(�b	���{��;��,p���Y��溍��w��=n�+z��5����k5�8�11������7HBu������<
�A��\"�#��u��f޺�Z���ޞ�xl깛���\�N����>�7�q#�N� B��"N^r
IA�p�+Q���{΍��d��<;��7��$Q�bJ��m� ��,Pq�4�Hfih��3�ɲ��54Q&��3�`iޅ�&H
�x�Ѭ��f��A�ͽI�(7;�N��!^�����o����N����S��u��~����u���z�����zN���@6���ݳ�X=@[G�{& ��6�#�\��v�,�UB5T 5Lɪ���k���
�j^��6+:i]�Үd�Ͳ���d mF��k�����<�q�Z�a��['������ն�V��h�Ks�7'�J���nó�|el��WX�F��p탈Uc�y��� 8K��v��s���<�O,=�s��x拚|�n���$4pV�����F�a�h��3���Y�:M��0��8׼E�w��כn�^8�'AЮ۬d�j$}tv���{4�ԣ\�]X�;7P-�CG	l�b�6�{/{Ҧj�g0�&ɰ͑bz%��m�ւ�z���l�u�&��[�؛������l��S��C�Q �;>
;S��"z � K�`�PC� ]�{;w��yo[ݼ��le̙˦k��t�M�av2��(p�,۽6Y�9�:}3�����sq�x(ź�b��5m�b���1�keu�rI&۝��!�m�f&[��F����|,�YqJ��h��R��y����5)I�~k߱�R��<���&�=�ϳ>͘�w���͛�����u)J{�o��P4=����)O3�^��j���׿bu�>~?cM��3����r$�$�>��}�'R������Д�Q����7�>Gr�'���8�=����f��kO�ι�k�pֹ������{��%)I�~���:�����~��iP�כ��J��vo�n�P�ə�$gx�yp��Ͽ��_}���j����	x˚j�ٵB7t����I<����os���>:����#di'�|�l+�t�E�](}���M
f�����p��]��m�� u���V����(�r[�$��U�����q^���̄����L-z-�Hـ�
eV�z�1�F�p8��R�&f���8u��H��-�6�Xs���u��Doz� �l�3B'��]y�/���o��Q���uU����o�N1;x�����vwU�^I���{n=����{_(��9VԺup�������^Gu8noJ��ޕ@y/%��t�Xyrk���W�\O*X-�v�c[�L�nmb��kƣ�S%'!Qa~�ϻ���/�}ݘQ^�b��5W.Ф��T�gYl*�8��y9�u�c�n��ߚoS��o<�ב����yy'����t}*CC{��hR7fe�&ǟ��
���uU_�gzwc��; �����xq�ⅹ#.5����vaA��u���Z�@qP�_�'t@�Q
%IB�(�0�2�Ҋ� ���%�yM����o���;O}�����:�o������]_�WO����`3�濾��K���Q}���i��!eۅ+.�:Sq �[��u��������L�v6�Ň��wN�0���{�_n� nf�Pw;�5����w��V\���~$4�T�J�nRr�Έ�Ӯ�+L��p��]>^^`/7zh1a�:w�y�xvyQ�.��z��K�m�t�y�4���H^^L|�Ng�xtT��C�4�H5���*�u'�K��K�����������ի��R�vܤգ6Y̿"��_}����e}����k*����Gt��r�_�$	����[�����zh�M�s�;��9��$��m��Bm�{Rn�ٻ1T�<�L�(p��α�D�(�	��w�[r�b��1`�b��Xsq뮺9��h6�<v�ƋqF��*j��=�t��Nj݅r�����~�����n�S�Jr�X�L�
>�X��$���<�0R[2���e����Yf�6o{��oz�l3��!"?Ͽ�����_�@��[���n�نxNL��z�l1�i�#�T噺VN��ם�@vl.�3��＼%��n��V��_Ԣk#�y��!�-7����^�ٽ���Gā����S�0����|~�~޳Y��9�$j;��]��5x޶��� ���v#�w7�)������V�0+���$y B���	f�|���O}n�osR~E�X,�y����~?����7%4���,��}�)�/%ڃG�y;��c\p]Y��ٻy�����%����~�U��}N�oK����ND/	��M���[K�Q���vYu��'>J�ά�ukKZ��z'��Ξ�M+�ݺ�����w��3n}�#�'��[�2V޴�%=��\�l��U��S���;zWZ}�ݎ���ߵ�+@��]�^}��������(0���*���{�ׅP~F�B�Ͼ�Õy��s�YG��+ܔ�RH��\�rX�� �����ٙ���y�� B����HH�3������1����s��#(R�o5����ef3Ͼ��]U�~�~�����/��#�K�>�K�v����(��Jb��]ئ}�)sӭPtWa����1� 2��0�Q�l��R��r�$p�w�Ɓ�N�a���y+����Qr�h��r����2�V�vI��9��Ӿl����~��-�ޔ�{�Լ���+>u��p�w'�I8L��c��A/�>���=x"�[�����+����2���y���3���7��y�9�ݾ3V��7_v��S����>�^���/1����౸ﭟ|{�$�B5Yh�Ӻ���u�l���N�Ҥ'���ϻ�5L.\���]E%\"��ݷ�M��c�8��n{v�oy��l=f��oF������!~�߯��������37�H`f�3��	�*���*C�S㰦�]R^���M��yI��}�p���/�wJ�I8����sog)����-Ӡ{�����뜒i9��~��})�35���n�iu��P�R�򙞨37�H���$���%����N+m7��3;�������ܙ��k��ћ�~IT?��R������7���R�GqN��1}ơ�
%<J�-9C�������f9Jt��כng��4'.�:!�""Ӂ%�{�$�ݽk��� �w^�h��]HN�dv�B8�4����p�ki{9$��`�]؅�wU|�� ����}�ć.�Y�_f����\淽��<�ݟs�"�#��w^�����gߵ���*��~����T����K���JR�۔����X}���x˚�n��~��s�Vn�$�T�x�a��zvj�K�_lq ^��P�1׿sW����	������f`���bX���j)�$�"I"	)`&a��
�����:,�Z�G= ���&��n�v�^w�|�w�v�/UX�%�fnltv5�j5q��q9���PnN�lo:�xv^�fL�|�3۷�m�[l����M\L�<�)]�����Z�ٍ��F�&���n)R�Z6�1�i�"���],�$y�rz��'��{���|?�Y_}���[w��4�v�����KT%'����-��A͙���*J�b%���3}�x|�޶w���B�����9֖°��lM�L.��y�_#�ޗ��!=�g��� ����}�Ĥ�����1����!�w��H���3_F���������i}���0ftq?y%�$�{�9�w��𜪩�z"��k|}�.���|�� �����W#�N�/��D9 ����l7���We�%�^9�;;��)̷/$"ʬ���3�,�ݯ'�ss��̽�vqQ�)i�$��ƚ��ou�P���u�����u�����[���3{��R�r�0s1A� 	��"�U�I�U�ZR��Hr��ϣ�3B�mv^.l��@��FM�v��5�I�&��.���s�a�]� �g:��/5v������儘�Tn�O�w�1�×����k�u�'��9��x/��1��}N�H��T �������b!�1DMS=H�3�z�t�{�H�������P�B�X
��������y�;��/�8��r@��w@n����3���Z�{� ��Ň���Hܒ�ȯ1V]�����8��& 
@~�߿��^����΍u�ߺ���U���,��^|���ʠ�}�~3C�-Ξb������A�>c��E6J�S�k����U��a{=k�����W����0�zu�wڙԜb�Zs/Զ��5&�'9?���"�L��:�Z�խ�;���o�`}ޝ��<�����]�ύ�ɶڊf&&&p�4�wn�W%�� �#Ǽ��K3��O�-Xf�i02�I�D��k2�RZ0ƅ4Ja1�%b!�p�M&�4Y���j
�� ���hH"K�!����`a���"��;��� ��`@�%b$D}��=�U�����u_g���k��~ �hQ$J��$P��7�i��c>��y"y�f��:��ޚ?���y�����/v>�����f����sz�kv�B��
 F� �	I�Qs�?l���VwB�X;�z�?����W�Ɔw;;���fc����A���`~R�C��;5v���O5�pE��o�o��۵��@�EeE��d�HH`@}�k���U�����������wTN0�$�'��~)!)%7��%ST�iF)�}�N�t^ߵʻ��}���� �3�	//{ ޘ_Kf�ξq�CT4L��l��Uy��>�Р�"$H`�^J?�S�7w� ]�wS��]�D@�e�p�� :��w� �޺��:@ ��N��v�i�I��ꂘB�<,��f��������<��8.vj��&���f�E������Z�ݛ�-�!�y`܋���N1ISa9�p�$�e��i�A�����E����ޯ5�Y� ��e��.xN�ֈt�f�"H���޹/p:�<Y7է\4vH��J��7�Ɠ�;��),7�m,�Nf-*sg0.��a��o�B�����#X�&]�h��.�y�q��o[��X��Č,u�E�;�4]�Oz$Lq�e�o�!�0֎kf���N!Ă	�pj��J7<���0�p�s\�m�n�-I�0Nｇ?|������g����Wm2��399��eY�Y��{4�6�L�l�ѹ�O�*�v��.���&ݞ�qs��q���c��j�����L������ʳ3˶���efffV��ۯ�놃t��d�]����g��#���v[�9�R���M�1\s�s�s�Ѥ�t��%
�e�e�����3yv@.� ��ZBl��j����<t���T�٣$9��^���Fk4���-���CT[���ya	�^gn��;,v����S	p�؋A֑�&Ԏ��1����HV;#��Yz�ˊ�wh֣n��vM>ŒCK[��h�V5
p�8�5҉s�ٰ3�ݳ�nײ��U_l��m����޷%��6�v�(KL�1��������"�!#΍��U2��G��ݔ�l����MY���59t�Vv4]v4]=�D�6��r�Xw`❥�w&���N݋V3sEp��;M��,8R����6�nJqڶ#��2aF%�q�fm��
ؒʚ�ƶ�]�኎-��0�h�d�w����.�\�Y�����W�nd���U��e���:�]��vƆݝ.:�P�e�ZPC,��{]��h�q����7.��g+�D�]�:�sv�L�+c��j�[#��%�:z�oM��gx��x��ܰ]�.�TB�԰��:{ֳl���-�'�!�Q�O�PЩ� |��A_¬�?�
��C�Q �&<%�/^M��N�w��wAߓ��L�UO��f�?RK�P��K�`����Ύ9@	�e˿��ߺ����kY��Z�7��vH8հ����T���J�'BWq��zL^�d1�0�b�n����@{�ӱ��vݦ�1s�</|,���+�pHL�R�Z�̠��u�f�����5]����:����v}�^�O�ȡ��~���΍^����B�v�N��$� ��{�4|�ޗ��k��{�����w���>�wq��Zy����b�7��t//]l/���_|n�J�r�r���X��^F�Gu<3vtq!׸���%�t)��ZG5��DX�؆���V	�tVmj�f�LMa����U���A��M]
)�kQ��.Ʊ�6�ͪdM:�����ڠ��m�L�1���k=m��h��XX+8ۻm<����[��uϋqZq�2J�B��=k���壜z��YV�Q���z)�4�>�n�+����@��7}�5{���|h�o3�淭sz�<�>�J�@�+m �ER4&�H֞Mӭ�&��'d��I/%��tN�[gs�{������Y6�77ʋf��1���/�}伓K��<�~��`��S���ݏ��޺��7[�TQ!�f[�Y22����}�/y�﷩P����ݝ���\>��]�)5i�F��ݾ������㯣��݅��_st(g��dS���>�� ����a��\^������f���L��˦��;ݳ�8b����H)T���S�fzs��3ٛ�{�����=L����-f�yraQ�|�/�3�������,�aX
G��u�̊��jծ-�)��8����]�)��A��6�ӌ��B��7^Κs�tn�oP�m�^6F(���ʖԻd����{{��F�{4�n�t�ٲ��G<�I�fGy�nw���fGu8_>�~���0���A�����3"$������ާ^K�y�*Aglu0kv�O�~����NDܔLq�*�EY�n쮴s�����ndwS�o��C�$hiO1�!�/x+7zhn;����0���V�5��8,X��Yj`V��ւK8���E/�%�%�/j��]�n���v�������tޅ���ѧSco;��hS1�M^Q�
�C,�s����)��$���p�u�)����I$�Լ��l���i��c2�ǒ&��>����:RQ�cHrp�@y�`��^f��~�U�{�}��237�����+5��4ļ�yx�Ԩ��:�/:8��//&n͏����}.`_qû�U2��P0�A��$��I/l/��ϣ���a@
[-�i��߇!;�be�H�hq�B�;��_/$���k�=Ã	�S,fu.5r��Q�q����!�����w7/���zWR{��.u�d���a�RlxS�l��n�M�s1��7`o}��������w<�yyw��Ni�q
A���wt�ʖ˵oc^7���wU �v8�䗂��˓Щ�b��$"J`��],{�Tu�7�����]�u޶{�v3����]I�mKv68٤��㯣��/:8�)��s�(l7��m{[K���]��<n�F`}�8�>|��\\^E�^=۞6���4f��a����[��\ESϼ�g�ey�+��{���Խ�'�R�V��]ʃ3�F˼∤�p����8�w��N���ݝ=M似�y�Ć{w�Q!y�n�"�J����0�͞�ݎ$��]M���$a��d𠙘�t<ǉ`���j����z������{��9�CY˓-���o/{�,Ξ$n��6����z�iX H`i��a	||�|s$@`'�:�kq�\��܉{]��EN�۵��u<��]�y��W���9��SV�4,�e�"���u�B+��8[l%�Ofu\k��i�;Κ�d)�]��h��t�ױp��awU,���{Śqs΂�3��C�d���$�4oGW�����7v��#�f��w]f YX��Jtrn{,�3Z�aN9�ݛ�q��B�i�����ںX/{��)�"�������`љ2����7K%D�t�J�HГ����A���`z�;�������۝�A�-\Dy�]�RV�ȢW�����k�Vv��b{�u��ߑ�{WH&9�K`�&��U��� |���m��)�����X�E�!�K�ivt�4����[n�FKǻ���zoc���H���'	Ƨ�j�po�{�+�%
յJ%F�`��x���/"�8���O�vR������ù��@.����g�_����^�:��98��X�%��!{v�gm@�wR�����]�*P�i�q��̶�[.]�Kv�` ��d�	xv���b��c�솱��f㮎�%�f[��u�SC:������@+�$�lm��e�/P���=�oJr$�<r��X������n��B�L}��/#ݻ¨�V(];���}���a��.��j��>ޜ]��_Pۉ,y�d1BiDU����}�@������s伒K�}��A�7|����
^b%�;�&kA��;�w*�Y�J�&A*|u-E�#Yf��f�s+���+��i �������N5����D_:�߷��/��b�p̥�\i�A�Ț�����8�>^�������UW� _zoc+C�SC�C���W)Ʈj�����u�}@Д�C$HHB��D�{���6u���g�o߱�^��W_ߒ����ɹ8��`��6��K_oU{���LwwҤn�����������vݫR����{��m���Wdw57�_���߫�C���_�d��V:ˢ�`}���������.\�2zg�3)�*O\n�I�ԃ���������Z�A�v�`O���5N��{f�o����"��LW��U+j���؃u�,�p��z\.�z�m���{���s��;�MLHD�S��G������v;>����]���ݾ0;�Zj����ӉL1	�%�u��Sn����L��L�g�dfXf��`���P�`���D``�`1�a6c����	t��dfG���ٟc_�����kms�&Z��䑋01��ޗ]�������e�wS��s�Jr�'�Z�Ӕ�p>�v����Xs�cc h����q�V�ݛ��j�{�p�!#�翳�>��~�A��*B�w��<*z��"�[Y�k����h�;�����m7�·;����y�y/�G���x���/����7�	�<@��ӴJa�/����]��w�<P�oK����ID�W/~����ٮ���V�ԹT���@[v��0ci�.��T��}���5�s{�7��5sw��`���aR7�o��?w���o˕y�����;~��#1��a�!hT��W`��Mm&n�VY�\��n�Mz����.���8�n���My9��q��Y]-��fIekLp�MISK����me�-ג�7oB��.��ˌy��s�V����@�㰝O���i��ޘ�@A}�_|}�j��߳���t0S�909RP�oK�缽�U3v���D1�ec	�r�Fۂ)�kz�,���a�7��� HB��$�o����7�Hۺ�Lf�W~^�'Xi����(Wm(��CIȣ��of���1w�v0�����tbc��ǀSˢ�Y��:��*���aA�y��s��^g�~� �o��n��)]ܗR4��V��4c������^BIK�����@{������'6����v�ycb�����ȼ��못�G�sP��Dֽ���������)*F��#vH�`w��~�드������T�j� cyj�T��U���k������_���׀{�N�{�zT����)x�0������-[Kf�������f�֔ݙ�%�t᳉�
Rd���"hn(8fi�!k�M���������d1œ��`�]o.���>���ߙz���m���@6���(ն�v��f��ceݒ�۪�L��n��uUW:��AJ�����z|��p�.�t7*�r���f������{sԜ���T��eK��6 ���{du���6��Aͧ�C��J�K�8�f�l��b\.�k�'��ד���Ŝ�8�n�NV�\܌e�x�:��k�R�j5Z^1 �fj ͸�E�0�٬監Q�1oW<n����7;�j��:�v띜<+҉�g��km��p��v+QuK��T����h70]2h�4f��3V�.�,�.������m��Ǫ���'�s�56�nqb�q���T�r�s���qc
JY�^4�0G<�yvt������5f����oV�P����*x+�*8���< h�=U�E������o��[����z5�5��z�6�mV�n6��Ur��+ͻK,4�Ҏ�b��2��e��Kl�y������vm�Gl5+J&έfzX��/m�9��Ks�XM������� ;1����c����=��B��g}�P{;��O��	�<�;DK����l�y�#��77�O�^^�_�K�q}�7߉����j)؄�@w?���ٽ�>׼���݌�ռ�7�k��sF�k\��"��~�����U~�:���
���Nټ���ɵqUD�ȋwD���Յ���N�*�ӡ5!��#J�&m��ԔN_����7^�h3�wcj���S�c}��;�vE�����Р�H�~�Nu#B��>�a�l���{{+ �:�|�͸GQcS-E����<��s���Ak0�"	���FK3)��h�hpČf�����Qb�I� ��)п��e����U����@/{gӣ'�r�JԨ�X�;�����b?UP}��bh��qt�uu4���B�R��=ϹX�+{%��l��{�0+�⹵)�˻r��`�t4�������U��BS���,�J5�<�H����:v�<�|{���4���}�8^�ޗ/p���i"Vb����t;�~)��GC�S��Br"C>ݳ��7���A�}��UP����wV��4���-�*`73z��/%��}J �������ϸ渎A�$x��mس��G�sUw���ί��O��ZS��5FӀH`)�F���i��@�Hؚ������`�3��;�N�{�~�}�u�#ڎ|�jU�%;m6�(�>Iy6�J��p�Ӿ��ު$�68��}���̖�*9��3�{��������\���4�;I���;G�Ҧf�!�gv���z�\���M9��HU�����UD�1���Ԭ]+i�VWJx�w����D{�������6�25.�5%)[�r<�7�8�
ϼ���������������WT��wn~���ٽ4���͞��'��yq����reʙV���?�~��N��������b���,������P�i����6ڵ��5�t#Y�#��S:���K,s��m���ݍ�"�N�^�n�ɫu*vdzIN.�]fᦙ�������'�3��^�j��K��x|t��z��Z!���;]Bܵ�Ų�Ys�o9�s��ϟ��g�[\��T�\p��nF��gl������A�2r�Z̠\KM�����:`��~���`}�w^}�*Pm�72��<S4E~{�^�E����%�5f�����y?�s��{�#�����ö:WS6�᝝�@�n�T�wr۴�9M�{�{�U�n;�p�����n#��-n�;ʈ�U<�QRD@�Ay�*A������q w{��V�k�%9�K*�J���~�/�;���g{�{�cf���������U�,�>\w[����j�m�n��.WX�����n��G@�@w��ށ��uaG{�}�{�ھռ��s[���v550�BDD�2L�AR^���� 9�sY��f��D�bɻz�0C�ɰ:�X
�f��[�1
F-�l#밶]Ŕ�f���Y0�b:�7�k[�3.�_OªL�\���&��e��1`�M��"Lt��KA�������փ����y'����|J����ʪ�wrZ�5P[i�+�J����o���;������6�e��U�9M���m�*]��g��wt���zu�}�T�A�i�y�(=����@3u��p��z\�^K̯�ﮁv�3����Ñ0��xp��ϻcˤ�R��Ci��(CB�i��4
&��)C����>������;�yv��x>�IS�6�w��dB�2�L]�b���Lf���A��wc�*��ŀ}���6��9��Bh*�!�4&k�~���I�S��^.Y�s�r��5��j�u��t�Cn�s2VR�0<�[���:x�=��}�R���@�4\ڔ�e�r��cP�{�ו�ZN����������p*%f)n��C0)��0:W��t�Ӓ1J֜Q3m(c��Qh�n`G}I^}�}\6��K��Ժ��Z���?*mޮ��9�ɦMHM�`�%:t�h��i`Q��������]h��� �i�l��\��nS�Y.c�V�R��w<���!&����p��>$����Q����r���8�w��W~�߳��<�,�.�)0�"R&sc8ek0-h5��I�/|_�]���^��ݟs.���V�"�jS҅L(&������w��/>��*ۻ�A}�䙯����wɓ�h��r�S�`}��� Y��U �$1R�ɤ��0]�W����p�<?��/�p�͕�n��B�Y��u���7<۳f��p��L��JEND�8���h�w^��{���ܰ4�+C�(ݧvڃ��~��z��>'�cw���5�ޗ;y��N4�V1�yFX�`k�V�v�{�+�n�^�m��.8Zjے+>�݌>�ӭ��݌U������S@�'[�u�٭kz��ov�C\ٜ�ͻ[EL��.�i\�%Ɔf�mt���m���V7J��@�5�����ҡ5���4�z�1ng��mM�ݶ0� �O,G(�t���BO����wA���	���䱗E��Zۤ5ҹ����I�$U�O
u��Mr�Ğˤ�Jrf�����޺�mfxM�hS�l
K�ڪ��H��'������5��`���V�p�(�fbn�n�˳:+-� .�r���L�>�8[n��}������5�>�,��!�7ު��N��&����~I3�G�S�6�� U�.�sQ������%IV�{w� =�uր�y�c��;��ħRX�̅IX��=o�qր��u��Xb�zoc4�k+��[�][�(Ձ�t��`�0)}uh��Xь����c�"b�A_���ݮ�owf�t��wԵ��+3��\�PH��n$I%Q�S�pW�-��8��sۄ�Fu�M��Fpg�w���C�e5k=�m��w&�B�ڳe�[������ӷ�3���B�L]��0ô&�a��� U�oS��B�`��^�F�iH]܉պr��3ޛ��I%v�|������/vKƚ�.���\���r�`�N,;�{|�y��N�eo�&��Wmʸ��d�ٽ4gG�F�8n>�H`^��TR�ǒ�U���n��A.�Ui%ֺ���z��א�k�yؑ�N�����-/v�Հ}�{��O�Z:^� FY��]7�"���k�������;��S�u�b��ה�w;�x�d��&7k�����4{�$�T�u�Y��{���]h;�M츾i\��feĳ��� ����m���U��P�?K�.���B�h��*%<EQ����n��77��i��m�p���j�l�Oɺ�r�ȓWR
�W{f�0Rŉ�q�j�wl,���5f��"$�Td�/{��<���c����}��Dd�V]��eJ�PJQ)$�J"��H��D� ���-�?l�A�����zoc=��N9��ӥq�}i���y`n��Q�zoc��i��}߫���CUK���jf�P]�}.{�TbHI/J�ԏ$#�$�geg:��t�G��HG("/�ʔ��	�j
T�H��]�T��e:��I�ԸᕆmZH9<�����.�����$�=Ν)k 5�1:�3l���������3'f͛�NGX�y��M/i1#�3,@#�3{˽��-�N
�Yd���.8�k\9�Z9�р��&��`��"�@D�35s39��N�u� :cSBd�J`�0N�]��)�PQ����-d�\:^�!&�$P݅�gZ���,I2�9)���NK�r�v��������N���[�Y�ih(�)� H�b���I P�اZ0"C�ƸC���0�L��o��Y�޶�oI�w��f��B�T{�9I%�A%*;7��3�^{��w�u�kZޙ��jܮm�U��s��fBb)�[7k3h�ʃ�*��<���J.vH�Pa�i7f�[��K��1\���p.�333L�ʳ3m�eY��kJ�fb�z��֠�k��9�q��Ib�	ۍ�ܚ��n����]���غ;F7VI�x�#��9�n�]�ntfи9�!�^.�ˇ[+���F��Q��\Pq�y�M/;wr�M��X0�3�T�ؚ1��>ڑ���t�c\�h.��&rsd�ր񶧒*�����xs����,,�lH��
i q��k���l�0:4�zRsm�`{���Z��cn{`�{c��&�x�[<Gt�3օ�fj��OC��Dd�Ɖ�tW$���<j�)`��I�-��u�z�.�6�mnh��/𩤲��P�<�ꓝ�uۨ�n��P����|��,Hk>����(o'�[p��ڝ��� u�	>C�d^.�^7'[�ۤ�C�[rFϛc��y�/s۟���w2l�x&�:*ZbL�"�n�	Uv�m��ֺ�
��j��Om�S+rvteR�Y� Ϛy{
r+��;[��Jk�Jg�����ݎ�za�x�i�c=M�{p��咹��==lr:�wM �B�[q��f9���ҎԖ�.g��u�ݽZ�־� FA�E>T�R�(RRP���� ��t*�  �> � �}{<���}{�Z�W}���Gﷺ�:%[�]JnA%|�۽y�yo[�� �vWZ3ګR] Qass)�f������v�8Ja$�����n�].ᇝ���E&���×��a�ݽ�yWf�Q���wR�h9��Pk�cpNFԸw�v ���a�����޶{ڻ��ThU�XU��i`sgt�?�y&c����>u�K�Y��L��[\��JE�Z�$��of��q`��؃Wj��/v�N��meۗ	���@��.{z�/v8��/{��t��1�2��̤q���r��%`U쵶��ۮ���8��Jmc��u٫K��LZ��G�V 45��ɵ�+	L��Lfi�1���r�C�2B�j��7m���ds���c��z����T�v�E����oh��@�ߞ}�Z��r���{ݫ�]�
R������o�LJ��.qmNƒ��]Wo"P��3�]����{}�Xa��gB��ŕvTR��ĩ�R(�q�%8��]��P{�{0ۯ�{ҷ��7y�R��˲ݍʈ,}��Nη�������7���Q�,ǔቬ���8���}�0�ں�}����e.�(+wv7V�_��y7Ѳ��p��>$vl���sn7�����;�*�rIw�<�cwK��{�����b� �a��$�Y1"J$��L"���D����s�� ߼��������Q��"��_��*�F��e�$�I������������MG4�n�ts�䅓Z{!�u�]j6��l�@�8�/e8S4t����>�v��5;�x'��j�GV�{$����<�Jk�p<��eHD6�9NS��n�f�ut�u������f�|H}�3�̇v�&;�$mg�!.7�&ϗy�^ w�u�/{o�]�6�����Wi��� �y�c/r�A�����v��ڨ�+&<u�f(���Ł7�{�0�������{����)A+�RR���wcW��bH��NJ��o�tn-Z.y�+v�2��;w� �۽x���g�7�&J˷3ˎ��K3
K�uJ�J���
�5�y���\��y��伽�S�n�f�x���J5m����i�a��3���I ��B�0�$D���:�g���U�߷���=�Xn��\�b�+1;�fRi�rB^7����Ŕ��o;>ݺ�Gz���O�]ˉ5u �Q��o^`.7����tW�ϒ��,>�y�B��U��c�,V�`{�8�?��U\+aV*m�.s�q�<qz�I��(Vv�����޶n��#�K����s��e�W���b�4,t�NP�$��v���]k�o�v{���t�����|�!B�������,'����7�~L�������� ��4��b�	V�N�$w�������\�^�����]L����ma��8��Q;C������>�>�`w�����݌�Q�t@N�V܍G`�w^2by
�H���%HN�:p	M�
CH�*�UJ8)Y�������r��a�5w&�H������s���o�.�\�F�<]c�I_� ��_փ;k{0��; �����;�W$�i��� ����ioN,9.��^ }���Ioj�)�Yv�%.���=��oR�o^{�u���݌��%����"V���������}Nݯ��vf�E1i/��O���d$䤒$�������1MkF�pv�sKl͍[I��խأ�zݭ:��,v�3n�Ĺ	^���j�,���sX�Og���s̙����\k�v0�7n��OǤ���K��5�p8��[���^���痝�&s����V))n�9w�3zޭ��j*� .�� �~��܏~��G�feݵ�)7e<�>��`9��BX�kH!Qi6x�V��R(鲤�I8���os�.�a�{o�;_I*'*���.��Hc���n���*��J7)�{���0�ws��~��/{޸}��K�7��С��n5t�������������,��ݛUQW̤�F���h�>�m�@f��o��%�������<�wkɆԬ��Hş�`���{�����Ņ�v2���M8�v;
�N���ޝ��]�	:!R:t�8*�/�퉝�faaldw�>_��!�zo,���ǊK�'I��L�(F;�	J�#�q	qĢ�� �y)��`Yy9}�%�׻[6-)��l�s���z�[x��ʮ)�f�i�5uC�lm���,�����n`�v���7{n�c�n�a�~�p��$vV^K[(cZ�܍/������݌�}�g�-��
��}@�'vD��v ;��^(���,o��} �S��m�66���5.��.������>����~��7}.���5#{����f���d�$���w��
mﾥ ����v7u��7�'+.��D�y�yw[�s�"lV��.v:�s��D�C�~qH�T�S��z��a۳���݌���WF�Q�m��cv��l�$�)E6��RSL���|`�_Z���v�]Xo��\�b�+��o�k[�Fk:��o~�")��(�^muP�oK��B�3k;���d��	]\I�ݳ�yq�l>�u���9=]h���Ғ��U���2�e���޺�<�u�#��޶ZϽ����&�4�����\��J�ҷ��<1'�./*7\�In��;>\����P��>�o.>K�'v0����~��Qо]�n�c/�6ۛ�D;G��as!TXcwK�ft�0{w��[��������]�R��H�y������ꀬ��z�3y��{�K�r��Z�\���y��93���}��s�G�6xRk-8ᬬ�B�$�e�5��-:KI�E��N�2!"�������:�^u�}�G���x�iO���ܻ�Hҫ<�j{��#u��Ͻݘ���Wp���V,xȌf,G��z�G(�l�������v�5�(����)�"GJw{��<�o[Խ�����~��������l	�P�Ψ��8�pq���;���A�޺�5n�L ��֨ϻR�)����d�%��U�w<���������w�},�ݘ�\BG�9�B۔;��zq؀�މ�#��/��H-Y���w���w��MYx	/o?�}�;�a�{���]��:g�O�;Y2�:��ݫg&�'IB\=�6�t)���t���2:��SXW�U�ƀD�x[�8::�e��(�fUb��k����"��5v�dWK!t��ܥ&�.��6\M34ʣ��E�]re�;<$����O^������
e�,��"���������J%Ce�C��1<�`���	��օ:K�����M;��������~�]�8�۬�� �t!!�&��޺�<�w� {y���zwc+��)w�Yr*�J���һ�rG�J�A�ov`η����ѠmJį$b����ޖ�齎���8�%��y�W��1ƛ���t���VdwS��o<�}�����at��h����D�v����z�9e��2��b����i�:�9�J��IF�m����{zY�/zwc����Z,��g9�s����i#��	�äeO�o���s|X��]%$H�lM6(d
i�K�Z�[�I��:L��q̷�:���?tGm�Lt�	c�-#�Ε���IHs��IQhrB��<����Ke�S�'I�3}\����*my8���J	�a��Zr
dGfiҎ�x	����y�&b�-�E�����dv��,m�R��*A2�bA���"WZ�Fk:�Ż�3���0[0�9��z�: �v�B��p3f<��l�JkM��F'[q\��b&�X) o �213%A�J
`��(Z
A���̱�j��XAL��j���/zuYm����|j��34(fP�U���uJ�A;$����U͆�"�Ŏ�9mmKƚꪬ�TJ �h�T'�;:ĕ3P8�TQ������YyJ�@���O�3�}��%�Y�l�������ƛ�.z��Dtɭ<��본G���K�Z�b��l�wZ-�G��2W�f��K���Y�ZG�-tpę��u�l��:R�5������mzA��m�Ǜ1nE�V����RWF�#�ݎ6m��cCKsgb�d�81=��zt��l\0�Љ.�r�2��e�n�Y;Kv\��6�#�K{x3�3��\�\1MGk��8��QѲJ���!��w��9z�=cܼq��]�lJZF.V����1�$n��9���,sP�-�=����}E}|E�!ڊlq>�s�����V�gw�����$�����^ֺu	ƹ7Zz4�������=�,Rtq��=<7g�n��u6�����3����]ea- ��#�?��I!�zSw�@�+�X�i��H��k�K �~�x�wKg�}��5x޶W�{�H�R�o)�U�Rf۲��ݻـ{��3�;�r[GNI�qʵq�J˓!ٝ�@^tq n��u0���4��4����H�dO05x޶w���n��`�힦-Ә�e,�
nTu%���ܰ����i�ԗ���E)���p�N�䉅&��]�û�ـ}�Xo�Wri<�o/�$��wݒ����&[�J6/�v&/x���`g�ocl7���Bϣu7���}fy��g���k�]�����pCmL��ʰ
 ���V� �B�p��)�z(�T��~�\���o, �-�t}�s|�r�U��]	�
�/68�5�z�Y2;�@��ާ/�s|����U�+�����}� ������z��{ɻc�Cw���1M7��,�F�|�����+*�I��Wu�{
�&i�y���Vf�h�Hf;oT�w�;���ɒ3LJi���%9$m+=�{%�N�a������WZ>�ʶ�JYj^,��MŘ�����J�`7z\7���,Է���'j�K�H�V/{�{ս�?��B�$TD� �(P�C
�D��4������Z����[3Ʈ�$ie��4e;�����W���~'�a��q��c��>���ϖ�%R~*~����H���v0p��ˆ��8�&T`��ء(�$��I��oup���0>�l�񫜦�K���*t4	Sm��~PQT(�Ԕ6f�u�l��݌>��,�m�"�D��r!�Rv�x�ˇ_l�_y$������p�>��mޕ �^k��ߓ;UDS�=Jv�]�|���]��G����o���K��7}.i����D�v���G!`o���{�N�}��yz��3��wC[<!��C6������x���\�W�39�R�Svnq�Nj�
�Y�p��rҚ8v,pE������٨���ɮ���u\Y#������;�������=�kj�eɟG���\���-y��Z�5��M�ڵkfH��P���ߵv��Z���HĞ5��Q�����W@\䜍�5q��\Ɯ%"8�.��S)[����Y�ϗ��؁�۲�Y��Ph�S�ވy&	�&���\���I��n���?0�l3�X���A��]h�w.��cnU��#2�ۯ�����a�������U��ԩ7"n�t�.�l>���-.��g%�v���Ki�K��̍�Ʋ؞`o�h3����!���{���qf���� i����+ ��l/��bIR��!s��tݎ.uN85�SM�()��q�=���y�+
���8�ا�f��s�b��0M��x���G;����X��cJYM�紳��g�s�"F۞�k�G{	��[���-n8y9tj��ʏ����x�x��wǛ7[�J���H���ay��X+3z�΅��J�H^RݒH�p�.�@p�,o��}�H՛�@��?{�yt�o����*�Ō��*L������ڻ��}�[h3�����*����u"�;�Ͻ�V����{}�؃�t��7ʻ�j��,̘^TLw�r޶��wJAʔ��������
�n6�n��VTc?!>�oy�����o.�g�R�ݷ�l�{�㵉.�<Ŏ���#�!"S�h3�������Ͻ�V���
�<��D��Vff\�%Vf��o�:qSE���JP�$��*�$�A	��Y�mi��I�Ri�� �TCqJ�I!5���&`7�(�Kn
a� �JA���%`%�5m��$f�ĳd�DBc��łbjA%&)�2��,L�ʃ$4B:jW���V�~�v�/[�f�c7���D��rU����y �n�q{e�I&k�{�;]w��w�ߤ�@Xܼ��)t^ }���V��J�`���@+w�B햻>��3Rܑ��}�{+�wMeBSr��v��Wnq���Հ.�-	 �vgspcf˅^B�b�9�7G���~��/��;[��BtF�q/�(����X�em�3�{h=���#�ߺ��n�ܫu!#�V�D�Vf�����8v>�,e����B%��3"e�ݕփ=齎W��s�*��1�%!D�H�P��1I��U����J sL�

(��AY�'N@�x�o�{�3�+m�n�R~*~�w;dV��^^m���3��� �m�p+sbB�gC�e��լ�h�^�ւګ��<�����-��n�Q��j�J)
B%�wLwem���۾�O���b�L�����15K,�п5ITq(��++�J�@g��X2����K�$��7���Z���;3�⊪v��NԂ���_yy;������w/�@{u������RU�q�jG%�ڷ�ާ��i�!t�^d-�*�mv�q��V��x���ŀo��������y�7�T T�0"�T��q.�	l��;�^4j�,lڲ.t������&��@��,&u�\+�]{m[`nm��f1�8����:��+]��ct��[,�����5�%ɮ�lu�
>C�i-�`�ٓN�۳�5�kZ5��x0����֧�o����j���"�o=�`\��Q4�Sto80X��{q`�̼OU�q@��mw �zoc(�>�a�w?�v�w־��?U��d-[+�Z��qJ��B����=�+�}���>�X�����j�T���b�t�.����{.#���A���X����E�N�I�ˏ�����r�H϶WZn�ڴ�ݘ�x�6��v�Ҷ*�����l�[��>��`r<��Ef��MHR�Y#/� ��K��<��P��]�]��LYa�M'B�:C��[?Z�������[��>����RݑH䒭˷u:qJH�h��u�n�GQ������Em���wn[��0Vc,*�&k7+r�fY�#�z+�V�mauV�2屩�w]���o��8m˻[��L&�Hq�0�[}����}��H[n�5{m��ғM�˒˧D��Odi���z�,�lH���y(e�q�q:n���u��l�,�Ҷ�f�N�a��]Xn���i4�#�Dǘܷ��}�ـw��h5v��g�jlȩK�WN�j���7��U�Vs��F�o-�mŐ���ܑ̨ʀ�i��z���n�,�ҶѺyiҤiR�q�Y0T�2~T��ddiS����m����vq`bԷm���n����aF���P�s���V�{����>�>�~ ��f($H&%JG�I�]e}����r޾���o_�~�w��HE�T���3z��]��N�H[v˞���]Ɣ��iK��{{0��Ձ��u�>��X}����)IE���Vf��z�~y�6�wN�J��O.x�ў#h��힙�6�h�����]�i V��圸8��N�s���_<�2˱Au���1�dTȪBJ&#�����>�������{z���Q�p�q<�Y��rf���`���3��
���^^Nݜp�J*~��+�G��������zwcg��օ@���X�H�7��qKGs�5�L�ll")�0�+r��)P[�3�7�N	�&2=^�2�b�9�1a��E���鱜��Jh��0��e)\ٳFa�͖�U+%�`P��Vٙ��2Q�j��q�s09�)$�Lq,I�03��th�1D���[w�N0�7d	`L��"Y��Hq�Z��\G��f���v�b��/L<����0�6�b�c����l��K
3(�1*q	+B�)���f1NK�ā�����Ȭ�l"7������MFʛ
,�4�I淖i�D��qa���Lk�w����zo�Ffk)��紹�����~3]�S�Vq�3&�m�fW���l�:�r�͎�gFz��`���L�Lö��u,h4].�[ōuv�*������feY���ʹ��Ų��ɤ�̳��5un{C�Zx��CY+��9ݣ4tn�)L�(Mfb�a�q�&�s����j+���6;�M���Sn{u��͵�`W���ӺCa;��#%&�[TY���Eو-�e�A@�t �d���+�[#Ѯt��0��z�F�d/m<��bv�f� ��z���p�{�;9ɱV���(EʴX�J�T)�P�%�xgc��;^.K\��
�R�D�+kQ��s���Fڝ�s�ӣ�����N�P�����ᵧ��F��muո��^��F���v�Z(�d5����K[���<v�p��Nr\��4�r��	��5ct��Ќ�iuԢ�ڑ�¦�����F3��9y�^Gg���]�Z[yGk[���lKq��@��1s;@f�+�추�5y������k�+]����Y���;�Z�I<U�\1n2�#`�%mㄜ�؝��g�h5˴ee�E���������kk��m�q�X���2��e��I@�1���c0�0�lS����UGQ��w�m
eVb��EbZ�6�T9�f�@��s5ͥ�Z������k{��{�����"� �iW� ��"�"'R� �Q@�^����SI��'�ayG��������ު���	��\��Zʺh���Ձ����`{uݠ��{0+�˕.����wM�ۿփ;Һ�u�j�OaR�)P
�R�S-�m�I��Gmx�m�������;1�����m}�p�|ʙ���Vy(۷��p��u�V7Bh�[��W��N�Ҥl;��3Ye6��v�+MH��}�����]h3�+��{n�2���Rq��-L�)L����[��u�ā��6\E^F�9��ܩ�D���D`j��l7ޕ��>�v{�/�Yk���"Q'I���$#Q��lF0-��b;k�EaŦ�m�cUZF��Fӻ8�ڣ��-ٷOG���t\�X�,�h�ҎY���lJ�6Ѭ(���iyuS;[�lV�j(�h�[��4��/!�z�grM�Y�C0�����f����B�q�z5�@��SI����=���`�UQK
m:Ŧ�\*�,v�h����'��)9>�o��0��o[��,+7w�v�o�t��NL��O�{q?��T����}齌;��V���a��+m���m�0���q�0Ύ'��1{о�͎$
ߣ���]i�m����*�n�N�gϹX纬�����}��
�wҁ!O4^3W�w�o[����X�+��[��8EWr��cWR�����1���}��ct�כ��r^]keh�6�)D77��ws���A�=֐��z2w�L�\�W�M��{�xDSD	�E�&15ΛK�kHB;]f\�-(��\��j��쑐�n ����"��=	����ڂ�8�mu���5!��W2�\XƌMo�ֳz�8`	❜f����R��F��$�u}��q`y{��R�ߝ{m��ݗ؊��sQ:n�wi~L��`f���[饁��ـw�o[7����iFc̴��]D���}����ocn�,/o;�h�{"���U�d�)���{o��+��]h3�M,7O-�*T��;hl�Y�_zV�0Nƕ�Q*��O�:j�)�sY�a�ɊGߞ��A��K�齞��|��I�?X�}�WF�L��7[�4��6o<�2�n˅^F���z�X�s�X{���ߝ8D<ne4�J�m�ι�W�(D$(j�d@bR A��@���Q�@n�ޗ!�㎟���n�Z3�C)V���r%�ݳ����Ӌ����ߟ�X{�Z:�PJ,�x'i�����y7lq��g��`���@����7;��F�lw#�t�$V|��@�U���0�ʓ3Yr�Pci2�r�B:ra9
��]�y�T�G�����c~-��M,���O�S���M�G�缬��v>f��;��{���|H^.�h�B�fJ"�"������/yKk�� [g���U�<��Nۺw�
���Ӵ�N�@g}����>^��x��B��eUdO����{[��\��Ӆ��y�L{��M���H���o�ާ��{��~��B�>f�ww��S�	ڕP{��~���^�.�*K-f�l�R7k�A�`Wa[=�����g��u�ǵSORd�v����'�{<z��dѹ������ާl;�p����K�`lt.�o�{��N1���f9V�F`o���߽��`�����ӥ�/�꠳yp���n;��(r�_�a��벃�zoc���g�v�#C��K�%+.,
7zKgGu8n>�H?��x^K�B=� �$��&������4�8t�º���mmڶs��Ħ�:��-a��N)L�5M��u�ez�Ł0�8�vʻ�l�b�;�lcVͮ�=)�:Ss�<нmZ��ڹFg�C�n�r<mrT��/K������9�n�o4f����.��>�9��~�V8�-'鎛�.��wv`
J�,��!�,�[*�!yf�T㖬�$S�d#�����5|n�Z{o"Zh.cg!�v�|��(�6�NSԒ9�1|j��l>׼�{f�oN�g�^�AҤM�\�I�K�0}Ҥ
��e�/�z�/7�mk�Ox�J�����1�09q�l>�wf/���a�u�l�i{c�jB�˴�ܘ	����;wK�3ft��o���^l��7���3���")�Q*S�������������n�sFmyf�-%ɗE�g�=�~�C﮽��>���
�җ56�ۤ���kQ��iK�vc6�/��z[/ga3v�L��K4̈́,���܁�ۻ9�����Ɯ�-m�'��bY�:�pv粋N\�.���nN����nA�f�rZ���*W����?�Ρ���Xo�������ޭIuR�5jS��*�at�3nt�S���Z����թ��
'wwJ�q
S��wex�S�s��p���Ct�c��q�Lɂ�Ff��a�{n�_��{�}������'?Yr[mB�/�v��;;/�bU�kC`� �1
�E��J�u��I������� �λ�����6H�x�Q�2��S����)I�SI褻���S����Ł�����������*׭A�g3�3�ֹ�vr�~��}קJ"�yw�"*����{*@��m���e��f�戅��
&���=�ܬ�]����_���zu���fy-}J�Tlt���K�	$�1��$�My� odwS����
�r�NSr�,yM+ȡx���`JxM9�ee&Ψ���^R�)I*m�Qg{��������뻩���v��t{�C���YD]�JI2�2�D�6�A�wv`η����V >���5:8��A�N�T�
1�f�א/2KfGu8����,W-�����s��aｿnO�IKTH4�D���g�IJ��{�+l9�6��9�wK�˚i��x��RSYW�}缬�齌/7�H}�I��~y3�ߝ�u$̤������c���HT&ӧ��qA\%2�g���(l��%�����p�^�i/}饆}��Jn��B3�6�o5HjƊ�N�Q"9�=�����t����Qh7�7����O�D
�J�"���9���}�\H���x��!��_�M�W��&4%*<��l�����a���U%�������N,+���NA;IԺbt<&��߲7���c��C�$�	 I�d�F^�����ך�f��7�S����9hW[tefL�wF��]��p��v�v��طh���y`2�r��,�^$;�Ǭ�]���G)@[�m)5HM�u �]Nݸ�x�^x�B<��f�,uP�ـ��᭗J�՛Fe,��t~Ns�������,;�k���˷��f2�`}�[��G���LilٌhnYA��2�,�"B&�(��$�D9����}�K;�}���R��8�ˇ�AI;U����b��*��Cߟ�Ifb���of�P[�Ă��9�	�
���i�X��X�7����r��yX}���iJ���� ��,���`���@���@�u�.no��B���D��;�y�āMfl�z�H~$���^���8�߄���]�R�I�M�缬�Z�⢔�U%���;F��7LN�8J�{w����׼�=�U��4���Q�=
�|����YjD��L/�D�N�n'[�قp��4�ؔ�ܤ }��ә�71�G,
j-�7�ͥ�2"������RuP�DOfGN��XZ���ێbXl!KrC�e��rb��P4�\�:5����̰& ��[9`�Bv�w���Z�F���k	��d4+����8��[
9����6�S�F1Ù�p����A�iFdh,jN�hB�9Bb�T0T�2�e���4@�D8�6!�Y�I�IE8�!��%:$�<���Q��+��|��Hۨp�
��`�F�����ݑl�vD�c7E@���euڪ��j���h���e�s�%1��p��	�\-v��[se��8�CV%�m"7H�	pj�l1��g�,!��v�vt�����;U�:������:ϭJ��Ϝ����|�+<�d�F��lmK���:�Ԋhj�㔺���)8�V�G�_լ�\�=�7���͵Ѫ'���q��˞xr�F���!�;��6tk.X���c�Y�M+O$�ݞQy0GqE[�]��T�.2��-6�GknwKL�d�K]�Z��8���^��ؚőh7JZ�b\%�`�j(�Kq�]3	�
ݹ2:ٚ��ky���W��C��]*��S�Â�Q��*��ڢ�����fs�w�w��^8�Z\�P�Wc���;��l�k�嬓��1��+��q���Y�[��p��愷�C�ݭ�������of�n��-�=����;.��f�͐�I� �im�K����>3�����`{�u����{W��&��vXܤ�{gv}y��a����G����4�Is|�m�˂�D������q`gν�������Z�T�'?Y�m�-/�u���=��սlϽ��IQ�񼱢��$^���g@�4���
X��icF�ܑ!A��\tS�D�C�����������{���|���GD�nU���:Z]iL5.R��]\�����TgG5���X�6\j�w'戅[�!���@��#ly/A|�\2�eH���_��������ɡӦy�x)�����T�Z�v\/��zf���C��˜Q�����Ϥ�/��3���3[zY��5���3�&��$����A`g����9_R��#��v�<�������R�&h܃<:r�4�`�Ε SY�.]�����w���B'iKSK�`m0_�8:mD�3�t����l<�=�������r[ɨ�Ԋ�HN�K���t�76$�+���]���t������o�9�*f"]�;E*>~>���߻�ݨA�l)�N�3A��ZH!dL̉�s8��;Cd�A�7f�*�7�'[Ey%]�H�f˔^�����Ԍ�;��v�ݘ�[��9�u�߽4���o2SjT���1�X��K���@�w��Z��`���e�bYn�r(EQ��m�������鶃�齌�������))I*�A6v4eiG0t�@��|��k7T�V�uP��Hj�5��PЩL�W�%u&`o�q`gzwckӭ{�ut���r���Z�&ԡ�}�}�;�+�$�o��_�fW��6�&�-KM5p��%�zXλ��[���� ��u�w�5n���U��k�7�n�ơ���5�Y�n��i�0�\�����R��3�6X9�u����&y�n.��#A(EQK��նW@E��n{x�ͣ�*�n��D�˷-Њ��[t-��VU6�U�f��[��󭶭���&�w{��{��ު�������[B8�e�[#����΄:�ҿ���I����J�[��w)s�LfiY�V��~}������`��],,��ge	����d]����͕��+����rӿ��k�쁫w�bλ��m/=��FU�r�\j�g{{0y�u��{��_{\�׾��%"��⬖����͛Hۚ�}�yz�ޗ�������I�j�Zi�|�Һ��饁����7η����j�D�l��Ǖ��V�;�WHWF���ͅ��<{t�G1�uðҟ}۽�wN,[�v���Ǵ�����!9q���N���&���4[���sF�5g��N.�)��-cv��Ӻ�:�uc6�]�F�&]kǜ�o0���q�{��mXp=1��svFť����ŽNټ�s��P�Ho-c�q�J+v�ۈm��u�r#=1{����0>�5u@R~�9I+N86�<�X�6_���:��9��C/{�I�x�~Vf;�����q`f�{0��i���^쯥�����R�2�����������J��ep3�a����\�C��ؕ�֪��!�&�{�>�7^@�|ѧ��s?�O���͛*gV���!�f`{�WZ�ܬ-f�����wc7��gRU;m�l�Vy�Ϲ��X�����(��ϵ��2��w� �l��g��7�J�f^AF�$P^�sH���%䙷_��`ߟ�B�����J"�N�M]+?�7����+=�]h=�M,>�MN��.[t�w��U����>��7v��Q���y��r���nu��@�D(�}��[��U��l��eo���,�'�Ϝn�����<H��I���wO g=�`gޚXw��0���a�ڒ]J��2�f7�Won��@���768�)�Η(��u���vyww���nF�8ft.��%�I!���A B�y�y'�����1�� fdi!W��4'�$��y�R�m�y�+=�]j���������
��?:Qj�J�5 �_���C�'9?�О{]���(�L34��֨�p򁖠;G�����̎�p�~:X�zk��S=D;�}~��jl+؜��\�@_wJ�;r;�Û�p��],Y���n9I�n[�C��b۽���,�1q�l3ηm�^�sI���,I�Q�0y�փ��փ�����WVֶ��2��Z.2:�ؿ����ϗ^n�,�ٽ����������8��>5�v�g*�f���0L�u&�1�#*�fU�he�M���k��ɕ���$�l��\-=�d�N��A��=N��Z;S>V�Z��'r[��UƝ�c٘W�`�<���J���
�^����}�{���j�Ņ}���*jByY��������/l�3�a�ƚ1�S8���Is�1��v���]��������t�g>�,n,}�C�C�F��y$:���|��GO#�=�������?S�6�P�<�fdi!����jH,�b����f�g-7m�y�����`V��r��N�7B�[sӭ���`{ݷ؃���g�j�\�n�k-Z�I���=�X�7�@�t���q�l����M�6��B[j6��۽�d��(�
����K����㵮w��sio �{N����[��=^���1�'��xϜ䓼�xj�mi	�6l]I����:��f�&����+���,��5!���M��]���Aѷ%�F�O뽃7WX�6j�b�V<���O��N�rI%���7t��.���Q�0�P��ڴ>l>�\*�8�.�4RwM�f�.}P�ʱ�Qn$�Ձ���pֳvS�noU��*C/���DcY�<����r�Tn�� ��z�g�8��-h�	W%�$����䏻��0�=:�b��am�|{m����K�m��$C�f{�8�$��ں��֯O�=r�pm�ۧ�5�)����v��}嶃����/~����F>v�~˹���k
��`�R��BQ�lm�E�=� �=������=6ћG���i���D�$:�����p˫�1K������W�Ӌ���Ef�n4�p.7hi˒���vy����WкX37eHZ�ڹ�n���X�j����]�����������۹�I���rZt$IX�]&�ܡ���_e7�U&%I�m�[���W`�t.��\����w0e��Pg?K�2wnM?~|�^p|�>�s�ۖ�6�Q����Ձ�齌�޶j��s���1:8�Չ��n�N�3�����Ł����B_j�G��sJS�pǘ�aԼ5Pg?K_B�l��^^G��D<��M�b4f����=1���� ĥ؆�N����X�DU����Ĩ]`h����h+0�kNk���o�O<;�#9�r|$Iܗ� �;ݎ����7E�Ӭ�ք&0�ܨ�J�K8���< Hh.����bP�$�)��3M!�F&��DQ�h� ���O02,�(F%&��Ⱥ��ߗe���;��`a��7&�(�CID���g4&��Z1��@�H�bI-���9,��ｻ(�dlތ�μ�aƆ��;5�:0$��sA��%��L1�1̙��`���Jd�PA.�D�AC��Ad�4FaMi1�'F��I5�L���!9=߷��}g�����m����X�W*���9�k2��[u�D�a��0�\]Ga�\�Ol���o[�;�Ę�h�W6��� �s32�������̫34��*��Ӝ����J��c�k2�H�T�J;,pv-�1�:���vPfn٦n��
np!6�s�1F1�{'U��o[�t������p.��uZ:�NV��x���ӹK�UaĢ�@v�ޛq����
��.S<9V�ԝ��e�]�'fw���YrW��C;tj���"]�Keѳn<�ޯ=Q����P���mv�\6��zܦ�z�6��dm���$��q����5�0����[���X2�WhxK��W4bw�u��Ӓ�5�X��G*M�D�p7eκS��ں��@�`�����ִ؉���횶*�e]�Zū��<�C�2�@y��v��F�v��o5,F�Úe�X��
�.�����k���fE���S-�O�%��-I��q��5q�1ֺ�aIn%�T�9h�le�m���L
��-��k��u����u�/!0�}I��mўw[��0��3Y2�c���N���<��gn06�T���	Ɲ-X���B"��v����v�Pm�U�RE���$r�ѹ�]<�ڌ���M����4�N�M.�l	�5���W�ƪ:vuvv]�Z՝ <|@� }P<T�@OT�K�W��H
x�x��(�D_A�z�=���߽߿u��߾�JD�5nEEܦ�/菗m����t}�y��eu�+�5�#�+3-�]�Ϟ����P�����B34�S��I�u�ȻZ'��C�s;�����`g�+���z�"q��W�L�mI�u��lt�G)�;��A�]��>|m�����z���P�F�.�;�'n��۲��b��;��a���WV�M��E���\dt��ϺWZ�M,��OK�� �]������Mt!���;�`kn��{��{��Xe�<���	x^0�Q���Y��̷�p̷�{z�:�j��Vp�Z�V�0�LT���[�8^	�8�����w��l6V]iNec�YJA��y�qŻKfb�u,�j�Q��?��l�c��B�c u�1��v�eK-X�vc���d�m���xn���޲�P)�P q��]�s��i{aQEV(QV��\���؂�ЌFD��M1�*J�䅚�y�0em�p.���ߟoųgD-���$2�w;�D8��K�v�<gIll�f΋i����J����;[���j��e��7_䒦Ύ��W���R6'm�j�L������`g�n���v0;���-�U˔I4���SQe���l�������޶��mթ�i�B�qZq6�ٽ�>�J�A�����u�e{C�c��2���dLy�w���r�-~�M�1�kk��5�rLXr$l�]`�&�Vn.���$
�ުk�� ];�w���s���5��3
�EV�����ҷ
^�ݻh�����bB3e���ʌ�5e���Ԛ9�ъ��$W\#��8�QrV�0����S�4����S�;��V�M������}6i�܈[,��y\wB��o�����F,�X�1��}ϹX�M�`v��A�����Z"Uܖ
�vX�;���ޖ$��綊<���F�W.b@2܊�C�0�����A��z�f�j�3ޝ������F��حRP���Xq[j��!*&q���T�U;���G^��8���0;���6�Q��kY����F�]�\�ѳq��N*h����ں�{{{2�>���伕8ki����s'xf��y�Mo5���<��뤀�{Uv�����
Ύ$͍$1Z�y
B�y�g"����z$�e�^�V��ւw��}�}�ލH���`&	�f�k;e�]���#���k�ޗ,7��A����d0ޜX�.�V3M�P`�0��X�j���Q��qO����`ooK>|}�=>��,���k�[/f�F:�d��Z��b�%P����������o]X/��a廮�>���jD�e���R�K0yo[Ծ�X�[u`gt�Y�#��Ҡ��".Ԩ�[��3cH�� B� �B! <�R����$�RI���@^o]X{�KN$t�b�e�-���\w[
�� �m�?<���������C�U˻LV9IՁ��;��q	e�g&�sظ����ޑ@��A������mՁ����k�鿥�m��N�y�	ؽ�^)� &�TP�J�����]X�=���M�؏�{3�=�0�"�ZEʊ���}:~���*u��~����ޗo�I����Jԥ&V�zu��۷��{�*@�|:X�M�" �$�v���;��3�\+���c�I �9
�
�
��w��df����kA�K�6�vƫ-�Uݓvy�`^��\V{6ۛ��P�ᬺ�z'O�:�٨κ'�1������&�m7.@����x�ަ�]*��GKAܢ�Lf�E��CpIN㚶�6�p ��Z�K66n*��^NI"�%�-��%Hf��wfPК�"�(iyNـw���S�Һ$(0�5)Q$.7q̎�bp�n�hX��߿g�j�ݶ���E{y*�"tݸ�t;�k�")���e�8B��·6li2�5���W��@��5٢��	6��efSQc3��u~�����˒޶��,>Ԗ��Ã�[v�j�{�o��޺�<��փ�l��R�C���ݙ�a�z������7��D�����vT���wS�����h�q5��H'p>�٥��9'��D���G�vXy�l[���ha�'2�����`��!{��!��<�o�K�-4@�͕�J��K�=�u�(�ե�65�^�7o3�a��d^9�����3ֹv�퇃J�fyրf�JGe䠺�X��rs��|�-��'�\�V-�]v ���:��n��`��޻ � �m�r�����w.���+�������0϶Vډ|��v���7��(�.<����j��� Sns��g�͎�s7�~�eS�����[���s���?:����5/�u�`r޶gQ�7�F�O.�\d�-b/w;]X[D����X�ĝ�D��̴T�#"[����=�����-�U�[j�s���ն:�fΕ����2"IJGh>�M�`{�����l>��K����Q�Wv6����g�s}؉���vs�]g~��U�ޛ����Nj]���^�9vcs!l�]�wS����k�rr���{�!�.���K͛�� }��U w-�a��[h���Ѵ�ۖ��F�$��p�%䞭5=�&�d;��]/����n�*�/<u6+in�u �����M�o�;��H��;��P��w��̷kD�[5ծ)ґ,�;�����l>��E�ý���[��NPj�]�Q�V{em˱mf�Wf�P��]�a2Ӣ4*��ib�٦��~�+z;���/r�$ iU�h7�@pC��T���_[^�v��Dԫ�#I<0� u��S��L�
v��ꥯK�aջ��FEI���WI��������r( �1��I��Nj-�˛��iep��p��/Ͼ!�{����;��QG��2�8�%o�:�}�KOg��І-I���9���.�4�+�g��~�W��&�������j]�^;�����`��ﱁ�]��}KvQND[N��ڄ� ^lwS�����9�y���$.���1dnfB��u3 �ޖ{eo2���}�+��j�s+��i�İ0��{-�r�kelM���kN�J�h5�x���M��M�a��f��͛�-)�t�	8p4���K���N�֨\b�Y��+Qػd�Z�d+)Y8B��V�����v9ay�\���Y�lb�qՎ5v@��ۮPZ1ŭ�y�q���͌��
��W�L��s�Dh�@�+�9�|y��s\g��7�w6�,��m�!�~������rL��:N�J��Q"���
v���M�۵'�sn�b;�/=��vi��1�����ݛ���.�fz���U|�7���m��e���T�%F6"P�F^�l�����v��3�i�1��;���i����oU}�f7~�����K�k��^I~Kv��!�Ge���yLW��?�_ٌ5{y�}�3�o�F��q%��xt�0��.}�{�y�R�5���w����6�GĆ���"�*��Jw1N��Yw���櫊�T3�FuPXY6�X++`E� "C�������7a��l�r��gPC�������l����TUW?�(������*���=���l�Hn?�] #�*�H  � u�����D`�D@� :Р)�L"!����D_$�P��UO�{�_����6g�?��24  (P��}�߲������Z����Ö���~������*�_ʕ=�_�6b]�_��_�߷�~����:��*��j_�K��A�G�����ß��\����G�C���G�������"�D�O��������]��1?�����<��?�����ڢ�����T�?����u�����tg������a���_�������a��*���D�TI�R�`�H	$�D�I�Rd�TI%D��VIH !D�I$eD����R�R�%D�%YTIBTIVI �RT� �HQ%�RUQ   �HTI�@d�	Q%Y%IRUD�RT�E�`		YB��H��Y!	��T�%B!%BB$��	�$RBa%P�Y	D��IBE!%VQ!	@��	BT!!E!T��BP  P�HU�$ ��FP� ��@� Q��P��%BP%P��	BTe	��BP`I��B@HBV�Da%@RP�YB E%	P�$Qe	IBQXBEX@����!E� �$T�  �$aE�%RP�YQ`HT� F���V@�T�$	BP� T	BEF�P�$�%�!P�T%	� R�	!	�	B 	 Y !	@ H a	aU`XEBT	Be�!V�eP�$@�$X �a$	XV��%�`!FRC��LH��P�Q��P����?ؑ�����������@P �֟��a�'�������O���O���_�l�3���F�������:������UѬ3������,�����������p�������|��s�p�����?������:��TUW��U~�������?�������0���\*����������:Kd<Hі�QQWO���_����A�u�?�8hw�1�����8�����6y�]���QU[������O����_�����QU_�?�w��.������|?��G�I�k�g��h�EUs�������_��P��QU\�=�OO����y��?����?����3{��bN�����{�_�_������W�_�X�_ޥ��e��~���R�w��TUW����+�M�1�{?���?����}����y��c��⨨�������w����~tx[��TU�?������?��������t�T���?���(+$�k9��P fC0
 ��d��0A���U�(�tu}o�� �*��q���hH��+�9P  ���i�A��^����t�	AI@�  }� �C@ �   C@    �@(  �@ ��(� p    x>�(I�M�:������})���^��wPݫ{�N��}���w�&�p���W��ݹ��k;��}E�
*������>�x}�;my���}�V��/���׭{oL��wj���Ʈ:f���F�^��G�^�N��"��Y���Ot�@{�����@�ܠ v�tP� tt�9(J ��
f]�CmѺV �7f��vm�  )IB	*�`:�v:t��L�@�$f�PM ���vP4�Y��ҕ��Vi�C�٠r�@P�vP�1Ke u�@P�A tk� 󷮯�yuN�+��gm�����ݬ�1��s��M�Kv�sn�+��r�[\ R/	UE*���w�=�\r�v������ރ�y��V�k���R���c^�<�������m�g� � �N�:��]�uMV����x��Μz9u���\�����M����Xu��  �RTB�($�y�P0ѷ�Z��\�2�Z�ח��s�=�5�p@u��G^�z׵�]�B�������@R��;m����;ڃ�������K-�]������ĭ��	�ӝ�vJ���  �ԠB� UǍPg:�m�<6�N�y�=V\�����v�=i�צ����n�=�{�t�\�     jy4��%Tڍ� O`EJ�  z5JF�� @S�)&R�(����*�*l�R��   �����(� �I��		������_�����%����.z���_ *����AU�
�*��( *��� *�� ���U9�v�p��p��8��?������D��w�tXIe�-�|7�>�O��&���=�f��a	ٻ/k�;�6P��¬�*I���!��T��a)��(u�w2��,v�S�<�4`Rk6JbA6nG3N�L۰%��qt��w��B�g'4^nA#�A�����8h�88 ���*cJ�틖��[U\ ����;�������x�d$H�捛�k��ǐ)Ě��_�����#�6
�����A��m��[��}׻�\"h! %"�%<le�V������ k��3��j�
1�➱i���y�u��qv�F+�g�l�40�����`Ew>�`�I �	��� �xxl��������MJ񷞆�7���!S�� �$X'�<�u�)�aS�p��<5��7���l�\���K����
V�t�Oބ�  t,s�5g��Qx�'wP!s����h���/��@O7)v�rC#\`S�3�!T��>%���3����f����xy���n�y��F�kw��c�B� !E; ;C�����b���B�0��.�O^>Now4ae�%6W���1�'��ԍL����oM����r�\�k�F4�Ѽ���i�F�;�g?M���aY�ۭӢJ����3d���i��x���K�=J�^&��	�"]�'�!V� �A����k4�a�4Z�4A���I���5$��O����tĽ��>��H'�6;vQ���g�0�B�5*b�g
�p&�-L�&���\���6od8f�=e��4Y���42(v��������RX9�wޔ�(X���I�'�A�u�n8��M�n���Fe�)=���S��h`Ъl�+�}5Z���'-ɿ1ᘨ�N���Pǁ xK����0o,�lu� �UU�����LPvko��Uu]_FYN��p�b��V��7@`�2�u=�8�Q���:�E
���n���Oo86v��_;��78�[}j�g�ن&��"��W��Bg,�{h�q��xb�7�Z
z^�	
g.�����1'	L���p��	y۰V�s���6��,ia�5��lU[��EmV 4�������4(R����|)�a吐�a�����`��cB���N6P�p�>o��Ltv<�3N�O<�xa<�84���V�~k��|T�4�Rl�\B�}І%ݗ��)�s��R<!Ny'�}g�$a���l*Aa���!��C=єә�puy9�Zؐ+��k|�&�$�Z���_R$�GSA� i=#�*�6OJ��(p �Āp=�����y��������h˶4����c������p������of�0'���܄&׆�xpnkw�ț���9&�}5�8`J� ��s�k,	]���e5����Jn�����тp�O��9G��\�xe�y��y�q�y����]VZ������������6BP�!��r\H6%� ԍ��f��5��l&�粙�/��w2����CE8�F$��: B��@�h���BHR��$i�6�K��bģ+���_&xL�c)M,Ӝ˭p��&�xk�%a|XFS<I�Y��x�l���|#	S(��qB\\�Bᤔ�C���Ѷ���M<�o�L��y�l�F�Z-���B=v��Y�`Tq�w8�K-ci���ݕ��A_xH"�G^J�ŉLYq(���7��=�d���
�Õ�0���b�z�����M�]�d�F!WJM.�ʎ�0a�`@�V5_G
(�Kyi��{�㿦�i���ӳ��G=d�x+;�[{���{�*��:6�U�� �B�^v�p:�����f�og
w�,�Rb|��,΋��xz�f�'Ftm��Uus��,��r��(-��`tP 
Y� k��gؒX�1$+�O�_��W�a�Xs��tng<�<4�a�¥=��}�$C�a2@��&����|��y�=�L�p%�kn���>�VFs��s;� x*���9��5¨�EP�;�#�;�$��Wj�Gt�m�p��B�4
̌_	D�`a�Z��AV���r�����W+}� �`(�� :n>�9��p��\�v;�G�~�*D���$$�!�HՄdV$���|�ap��6��Bt�I��&O� ��Aa�`�����1H\xˋ _z0��c+x
�WH��\�ѥ�ӡ.���1ܽ�B��b���r�ч�*��0�.z��O�08y�C9��c��o\xd�^��#f�SS�4Y�|�z}	LrM���d2�1�
���o���u
�F��8<5�zy�x����&&
o���y�{xNkE*��6�R�A;�\.��T����Vw�8���#w��UPv;C��gȂG�@��
\��)����ayHt\(�W�'Ǽ����[]���3w�����B<�����!}���p��B�h�F$�l)�Njg&�#��B��V5��S[�H#�R�� HB�BB�P��e	g3��4�5�g=�0ӽ��<200u�g<5Ƀ����3�i N0$.h���IM;#�s�rM_<>�,�n�p��c ZXeb1�X,vr� ��;���N:e�ORH�O��"����q�.�T�����+\;#�p��O}˹�/3gȐ#��a�`13S�9�k���Kٸ3z�n�B��
�M��� g�L^���{�gS���]o��0&�_o'��56V%I0w ��0J���]�᳛`x�
�F�l�x�aL�7����p���5N</��44����g���G
v��B�;%���}�ds�i��/7�u�B���~y�� �x���!3���_8��0�UǑ� ��fs<�s�{5����#\4s��=�o��c��`�#���ă�܄(i��	������k>OC��Yez�a�,8J���FH�#��D���X�Ah$��g���mEԒ,��F^зƚ>'f>='�s���y�y�t+3�X\�%�sG�Ԍ����4��9��]�����!P)����ͣ|��:����ס� *g���9b�
幮��� >� �]�&y`���~&�5�K�e�|���Og��s���L/��!�S�%�!YBR{1K|�<e |q{��6����z���8��kyy���~ܥ6]����&r��ӳ�F�K�k-�/�(SWWъ�S�G@  ]��Y�XN��+�t�d)��R��p�ˌ���d=��>��[ ��Ѽ��Lw��L[oGA�Kr�p���6�.���mXQ� }�a��4�T�������5������8na�p�	�M�c���Jy��J|H0b̈́1����T�3�����y�֔���`��-6g�{��}�q}y$���.���8y珜�\�!.t��o��<Ѣ�`B��Mko<5����x�+�+���G�&��*b�|4n�SA�|.1�7x0�������Ja&�@Fm<c\o�ݘ���NO3<¦�dd��{=��6}�G�C^>�� S7��洗�N|����"\��bS���dhbiHS5<9�y�Mk��9��Pw��Ȇ� �]��;���|��B�Ls;C�c�I^�[c����,�A����ݎ��q��(:��y@gptr��Pw`���β�$�-h@>������7�a		�������_��!L"P�I!g�Za�����U;Ya=F����U� �N] ����*����D˻�Si��5#{�g��`8�ûC7K�����e�'.��xUe�h��ˢo�i^���7�.W�������V��ߚ0#4��(�Fί5���4�i�
f�h�5���Q��4�%��5�W�
��f��)�����I��?xi�T�5*`�R&��hv��y�Ee))�>!�\�4z#)*L�4f�Fb�@ &I
>H)��|�ξI��1��-&� �h�t�;��1��ز��m�)�_�b ԗ��q�T �1c�� IB��S@򈀆��M��I�;�x7�ހm�J>��:i�ύ�~�����M�����>v�\*N�c�����Mp'9 ��]ү��!
��ۧX�oF� �'���xe�ˑ�ġ�������B��/��`0�*E��Y4l���M;�7�=�t`l�p4�D��M�%��[VT�[p�)�k���C�F��<��B������<�SfyzQ}m^y����~%
<�`Bس�w���$�r��<0䧆�k�H�Y�|O9.�S٧w��N��L^�R�X�eϑ���%6k�XK-�˸Lײe3����!�<!�B����j�-޶rA�5�6l<
�x���Ro�H�vW�<%8�B�;"��P�:	Ip�+Y���X�I	dυ����x�}�X����6�skpѽL4�7��=P�I��<�?���;�餐-�<X�#L4�����S���oL. مJF�a)������xħ3ݼ�/��^r��1��&oX�!��B�=E��1!X��\FJ���	a/{���hy���W��Q������2�Ba�=@�����Q��'���������SA�y乽��<Xq�Tt1�e5��d��8��6��� ǐ)�M���[��sr��R���5LF���]u� ��ٵL��l�*uj=���Y��3�����C�z��.�4ռ�{n�:����֠[u�Ov�*/�������y:�ws��;����=�U 
]�T�9Ps�>u�d/�����F���=�0��w���8�Sz޼�	�M�O�<>b��Br�47|�^�v2��Y���|I|�W��y^W��y^W��yY�${�&�#��<�#��<�"��+�=۪E��+��+��+��+��j��+���y^W�%X�<�#��<�#��<�#��n���#��<�#��<�#��<�#��<�#��<�#��<�#��<�#��+��5vś�M�^�h�,k,��I���b��b�����,ʞ[�B�<4��uc��꼯홤����T1/9ᣜ�o5���{c���x�=����.d��Ը,9kd��g��ً���Qo�O헦�`�{	+T���n����O�꼯+�#��<�#��n���#��<�#��<�#��<�#��<�#��<��+�򼌆(I1^W��y^W�d�wvI�Yc����yG��yG��yG��y7d�wvG���<�#��<���G��yG��yG��y7d�wvH�^G��yG��yG��yG��yG��yG��yG��yF3��2��[U�z�����yV�o��c��YG��yG��yG��yG��yG��yG��yG��yG�^W��y^W��y^W����+��+��mW�+���y^W�G��yG��yG��yG��yEy^W���o�r���V���G�̍>}4���n��uy���tj[wt(;{!M�{{��l���s�,��Ni}���*3t0+*x;�5�e���h��G���z�E��=fg� ��,}a}�t)��˙��`��J�m<����[[$j��[W��Y����ςOu�9����"�Ԟ�ʻ���-��pvE����9���Q�\:�R[��M76d�A��KD�ݱ����{�^`�[����G���gLY���pZ;iˮ��W��}lx��m�r�a���"���;��In}�]�oZ9�� ���a�|w3����R�%��wV�l�5������q[DvPpՙ�L���G��	�����A��I�7GNy����=�Ō�L {X�F<�o�2%TZZϻS��Xpi F�׫��}=�@�Fb�o����F	Yټ�>���=E�3�����3�>����n�o�m����>>+��=�?M�O�̿��|��z`0��2Cώ�[L�2S�6�K�M��-����٦��@����]��gLD��\��ya��s�ࢾ��8۵[E���RE6hү���<Iز�jd�6j�$�����i�c)/ؽ���.���^\gW�F�{'���2N�Cg�@
{��䍍�{5�mm��l.�-Ndʸ�<�x���uI==���f�ujZ���;u;�����sk�׵�q���|�I4����`�;��ңt���Vsd؅�/>�͓�>��|�N���n�}�j��p���mbt��oz�l�#���d�diS��3~{�g�C���}�Ÿ��$qz��/,[�Q��L��>тņk�d��xwL�V <G����OV��:f���x��I0zV�q��/='�&��l�y�F��hd=��t�'ulu^ݢM~���g�#�����)�f�1Q_��Xd`n��hؓm��JF��5�]7���V�!��,U�������i���mV�M���Q!Y���>��J)C��ܟ�{�,�$Vy�Ҧ5@ǆ����箳�	W����f>3�J�-���M$ȶH��J17Tsёw���
C�u��֮x��Exd]�D��n�)����'��gI��p�������˞'A�3�M<4k9�*�*]4�i�C�zK�,d���u^�8a�9I3yD �����F�r��y�xL��:wFd�P��^b�<�U<my�Fw�� ���~K4��g<�E�����[���St�$'ŭO����0]���Dw�����vr|��7�߽k��&�J�Sj�#}.�wM%�+s��7�\�m�֤�3O)'���'j�7um=s:�Ky�͵b��^���ڳ�YE������XV�l��C
'��_/��v��3�S����M��fg6c��6u�a�C�;3���o�vI3u/�4���i%N�3�R�.ř�{�Ӥc��s��[!�y|�K��k�W�鋺��%fm�rn=����x�[�7nH�at��v�}%��\R�<:�K]�ݥ�fh�q[j o'�������d;Q��M�]W��y^W����I�0�|y1V��$sQ�d���gX�: گ��@�.�m����wm��u�qAe�;d��*�W��R콩-���TԳE�y���ʘ�����3�{��\��kr/G���;��^T���.���i�.�^N0d��V�z������x_�d�J�r�/��](n���%���QD�dO�1���\�n�m�� �Xd�
�Xgq$)/yi'���3�ދ�V��\3ӈ��u�<���пl3j���Kz��#��w�;pwLy����=���u������->Ȓ�c"b׮ĵ��	��=��Z�WU�yz��$��"��S�V��$-��Z�*�\S��z��L,�NX�mQE�L̈́�˝�N��4���cͱ�6�WbQ�J��#VT]���&�u��k���_����M�f�fZ���)&,���Ξ�^�Ҷ���C�}��M�%x{����m�uo�L�â ��ˊ���mS�ԗM��@��ՀcŰB�)Ҕv��E�[Q����6�0n?4�WN0��ז���JK�n��H����17�<{MOU�s�f����a(7R��횑Gq�{2��@6GTwOQ��m������f^W�{�n�\�,�r�jY������wh�ˣ��U��`S�R�W:r�j�/)�ݲ�u1�h
�]��n��bӾ˞�D�Q��k~ߦ'���6�����³H:(̱�2�ZާO�#tM��rğ��ª�^��8=�3uf�]B�1�EO��X��;�i$/���ݦ�ڗf_M��3�<��y��{�ϋ.쒛2��em�pvl�xY�^�x;c��RΝ�����f�ݓq'��l���sO�Jх��w��6�.Z�U�7uGW!��ǣٴ�x7��;
���ĺ�4y���.�^ջ��l�j��ȷ�a�q�\okG���uޜ�^۩"}�֫{A��M^W�I��E<��,粶��uj�WU�'G�$:ƕV�#��6vݗfӫ�}ޛ��͐go���;|:�<9���Q�,�`T�>���o�:�1�n�ݼt��2�y�z��~[���r����R������;<7e��I$��mLkp�H�q��k2qBI��z\[�����A�VאH6 �j�}`��y^W�cƍ՘��4ψ��tq��+N��qv'F�X�~]c� 1��f�JԒX�S��!�X�r����@��7v�]�3���{F���f7�h�g8Q,n3��w�{�!1�����є#�n��ު��m^�W=����������u���r��-�Q��F�2q�<d��ʻ����������~"%�I
��n�:3��C�����ϥy[d��>�ɺ��.����,�:�<��WO[��q �=�!����v�2>���(��쩖��m$�x۾��=0jT�V�i�Ş���"z��[ۤ6j��;�#�{����"f=����Ө��ܛ���v�}��{"�ܗ.��~ٺ?Y���ZmO�.�}'[��,�b���p�&rމu��ϻ���Z�.�y�^thm� x��j����;5ł�a �Η�W[ۙ��}$'Ӄw���Nat^'|��|�N^�����o-���9��:��.~X�m�v�=��ݶ��J���RcX� k�~��x���d�7A�U|Q`F\E�7��%V��my!�w}���wj�5J���{/�yド}�V�Q���"�V��[���[y�<w^�ji�/��N]���t�ms\��ݑ�>��N�c�H��)���t�H��co��f7]Ԕ;�T�w����'"�u�C�1�`��?6�¹)�%�˹^W�F�]���j���$��Y���L�|�S4�����C��ۺvMZ�g����No1�nf#a#���myO��p��R|:Y��ڦl0�>���|�U^����V�����m��;�OS�DH��MKTm�S�L� ��DJ��&�d�y]��kn�r�W����.\ �͵�A\�k�v�5�je�Ms(�|���Uuw+���wN�6{�m^]�L�5�j\���wf���ܫ�l�Z��e�M��L��tǦ
��2$�3Q�u��n`�'S��m��y^W��y^Ǻ�n�f�����Gˎ��8�qnj���r�=����	H�͋{�8��5ndW��U�I9o��8��hI����9.�d�~��l�50�lIr�|{k���8�9��E�"Z�����9�����yn�dԘ}�v�[��'Oit��v.�f�$W��j�R�r��ꎢ�ԏd�׾����%L`�l���t�t|�<$+/�"պ�<+qC�`��9MVԇ;�rz�U�՝�3�|�-�{�S�Ey^A��SU�֛��\���S�I.�y^W���{�t����8��Ǻ�qɞ2�đ�q��)�7]V���I23��d3��v��=n�x��b�ꤛ#nJڋ��Kr"���W����m��I�RVn����'�*�$�U��#x'w�G��U72��u��'��[�A7vIpp�+���-�����$�|
��=�w$Rd��%$�c��%�ڮ��Clcm�m�vO����	@yAr�1$��Iy�m�l|1/\�1��6��;�7�Vn����Pےyܞ��c���f�۴]�6���f�T���g�iR8�뼻��Z.d���M�n����m�r�ҦQ��ὩM\f���r���9!��v�/�Sگ/+�<��B|F�S����?���c�w)(";q
㚫��l%�e b:2v�Eɉk��+'����H��:^��7���F\���Ik���ay�ZH�Gd��8/SmZA3foL5��������ˋ{ފ`������V�Y�h>oU��u��1�&�=���{�e9\�`������S���R�Cd+�f��KRO�b�u/#:%�Ns0�-����{��7ct�U����j�7=�Ó���u�p���A����N{+ <9Z�3��춑�[�M����F��߸�<tܿ�է2E�t;0?��`&�V�F��Ú�VZ�*�=��%j�L����{'�/���d��O�G9Z��U��~Yy�+�r�o��[�sk�x���٘��{���Z�$������%��5wt�j�G���D���̩�w0w��n��P.7��W��u�ܯ�����&��	���U�y^E'y�<V'�Cd2#��s�y^I/=� �WU�[O�R�*a(B����� (���!<.�l�4�դ��D�vJ�)����)��!�h oHwf���%d�5�]�d.��5q�.HOmǮ��J�+���L٤���p ��wF�%�%�ɔg`��5�۟1դ����0�v?Aկ��G��u�=�rI%܀�� nH��K�+�$d�TJ�\f�䀴��F�@l�����z�ʱu�<@��r����6o!�E���x;{��m�u��[�u��OՖ��]���z�O^��Hs{v�ݵ^�S�մ��|d����!��:��j�W�h#� z����d��P-G�ifENc8�ԻsykH ��z�z�΋l�ռ�"I����<�,m��V(�wo]n6�G��${�Y�Hٴ�S{|�wV���:��$�-+{m�1r�{���m��%n���.�7���9 ��jI%g��)z3�*��&��]��H�4�;&Ș|�+��K��@؝�s�G;yЪ�#+����U�i\�U���Z��j8����<j�+/%��-��$[q��!���In���'����g�fr���oV�I&d�^W�/;кV.$��{�\jk��$�t����{��}V��(��g����!�w����o�Jfh�IuӁbb@bOv.�Ep���{�]��,ӞN��4�;u%�g-Nz4%�o(��NZF��zj[�$!��{PȵJ���>#o=�����j���hC25�����Xy�Q�c���[�d�Aog�t�i}z�^���xpyJ����ޯݻ���/�Ⱦp1=&��6M����:3�;M����5�;��v��EF�f� +C��\8�P��c�&m���a�<��̙U�n��nM�����_��2�4e3I��c��H�Ժ�7q�v>��������zA�=����=�;��ɏ���&�7N�r�)�R�ӥ���ǔ�1�sbi��{�~^��>�z��5����hXwt�jvn��3�����%}o?�z͆[(��סQֵ��Hd��"� ^�fj>~;��\�ܼ�0y������ϵzG�}���y��SWn=4˖�C��pm�..���v�f	{���ěvH�v��z��GJE��gn�[��F��D����=ރyZ�fm��;�k#���!]�����?29"��+��+�>z�3��!?d.��گ��i%�����X�u�w�s�o�īX�����;ԉD���ٰ�]��Wj��*ꬺ��׫ws�M٤�yG��|�+ʙ�D��}���W�+&�_�*gxR�[���o}I �=�yfpr�&�fػI����<��k�wQ�gӅ��7T�\L�":�+�Wt}h��uv�4��Vj�+M:��ʖ�z�������xt��vD����'����'t�Kf��+��䅝u�N��r�W��yT��z�W�=&�xf��7᳖m�N�vC$�Y��z m��i���k�f�w:�Dzut>�TKy�
�]ə f��"{7uv؎����{B<��I�YYfZ �C�p�{���cKc�~�
� v��=�^+c����g*VŹ˟c���w��h�p;�3��5]����d黻�l���������"�0{3��ÝS���n��e�7��Y⾪����X��>#��L�z觮��y��QAO�P ƅ <��E?)TT:(��S�����(z�0T�Pv"�Pv �'�B(�PJ���@���$$��2aČY!�#d����$HF!F2#��F2B@�`0 ���bA����0#�$$0�0a!$$$ B0	1�d�� �"����c$B��HD����!	>E�U��� �� :����/�(O�GH��x��� "F1$�"F(BBF0�!22# �"� �� �$!B2,X#��� �$�$�#�b�	� ��lD�
&��QpDJ��0F�Pt(��&�"FD�T�N � ?*�ȉ�D���"����Aj���
'�TJ&�W� x��U�����|B�m��T�0 8�� ' |
z�DC��� ~a + ���0�! �����@M x�z���B '�i6"TAM��VC����4�����-@=G�R*�P�Q���x�qU*E|U`����H�_�t��
"�(���ҀTUJ�(���ࠀ����|��P�O��j�
�����,5F��1����f8\�l��U�v�D,z���Z�������6W�!��.M���2	3,/CJh���������F]m%��j�̪�˨b4]o[,�h]�Ex�nu����v͸e����c0#s�$J�e�!��tn�uR��vm%!@�u�f�M,̲���J�XXM��s���Pn�5�m֍�7D��!��-0͵rQ�c�nŻ5q3sj,^6k�[��ź�����f��V�a���7vXkY���+�E�d��c�- ��V��ݴ����dfV�cM5l�ٰ���� �T��t�����(l45���h�v��t�6�.��Yu�Ɖh��M{U5���$���)�u/��/
A��">U(���E� � ��U1~�nܷ��ԘWr�@�f!���f[�F��3!6�,l�1���P�P�����3LL�L.� ̂�M.��^��Tv��.���+��2�x��V����v0/��(v�(}�p�)�Z��fDd����wJ�lΨ>^7�����]J'k��&�%@�{9uA�=�@�t���z����S,��	Jݳ��y�X��@�͙�f����U^G\Ģ�>��TQd*����Z	���Ue��5xn� a��DQ��eWf��>׼�}�����]]����i5�үj.����G�q�1����`o��P>����z�|�|�x�H����ޤ���n�ȊQ�[����<��ʁ��r��Z�ID�1�]�{��Z&M�,�s��b�z蓱Og��S&92*ӵ��G���z�!�-��k��9�6]w��6�B�Af�7�8�S����	�NLL�]�gQ�)F�Y���A�t$���fM=��e���2h��8�|[oƧ��k�6��a�i6X�����޹@��7���Xn�bƞ[q��@��ެ>כՆ�g���T}�5��"s-��i6Ѻ'3e�$�lR��%����[�Xow\����L��ǔq� KL��L�k��;�6]ݡ����2@j~S,�"أE����wnc�FT�лDj��$+�!��D�<Q�бo��Tou��yuG�wH7B*�Yq��ŷr�ZB9�1]�;C����X7z��عP�[�>I���N�*�qXk���}����oVY�Z;�!����l6TŒOvGd��R���F=h�Z}룢"�T�ȫX�f�7�.TwzP>�{��� Fb[����5�L3L5˥�ۣ9��5�YX�W�q����פGV1��j{��W�]cɋt�iu�3<�yiU����Z�!y2�6W71fڢG9u [�Ym*��X�
�;.&����4�&
�k��Q�,��,5B�M`�0n��"o$䜿{���p�\��׉�6
���]P58���Mel9��c�U
h�q��u���͐i$��vI>�}+=����OՍ�4�p^r�`�ֶ�:���}���ua��Vn����3������*��v��fuA��o:��uA�o\��{�Ǉc����;&I
�ϝa��:��{�����7Cy��Ȕ,r�"�I*ݽ(�7�������t>�p�k��e�JcN�,��}<�q��|�f���+�Z�dy�\�su8����￯������a�.��%��تX�L2ź5jR��9j��^ves(4�-�[�k�U���{0�L�.�,�k`Kx$E%utP�<�pٞXF� �0N�w��ϥ�=u�v��J��hRUTe��I'1l�'f��=�ҁ�y�Yܑ��dn���L5V�����Ü�"r)�sg�Y'�����mE��ps#�=�3���� ���a��q�}��b}���X���J��y�Xo�gT/f�n���n�vFX��<r)@�}��}B��حu������`�����0m�蕶�������8�}缨o��x������1���ג���:U�˶��=�z�>ݙ���*��:�;�xj`e�t/�3)_`�~�wӧ'ԒIH@k`T �S�.p���s��G�d�Y�Z$�H���W)�$�Tn�i��P>�����wK$�IaZ'�uKG����㴪�@�!(�L��ػ��ޔ�ӊrŚ�(��,O+q�݀o���R����6��J�����]�e�
6,�"#d�ݻ��7�;��ޔ7�11�ˍ�"#X�$L�'�Y0���H�
���]Pn��@�tΨ��z��a��H��GVT��'@��8�}�3�}ܥݳ:��%��pJ��V�qV��(N͖*׬s�<�p6v:��fG�dﻦ9���e���qƪ�bެ��({��fuG���5B+-�׍ȕݳ:�$T\�b�~`�$
9�k̻�G�Q�Ts|�R�wN@Ӽ 7���o�?)l��oe�Sr����s�Zy���P`��$ �o1� �����I'��J

��{V�a^H�;���-[��0�O2����o_�[��x���qT����0��p`ux�`���!�4�?��>����Y�E�|��s��)�e��}��)eibZ��M]��B��U�m�����ͥD��]k�ۺ����e�A���f��Mn%�ņ���7ȕ�����e���j��-d�\[M+SR�����1ZR����hR�c--6^�:��MT��n�0���!��[)c��Ak3#������9$SX��필Dd��WmإWM���t������X�lԹ�΃[sH��h"j��L�,�[����I���$=�I�*]R��h�Z�v�y�|�Q�-��8-��[6����4�=�Ij�b�$�`cgz�Ei[� ��� /����/`M��K��2@W����� ��� S��s7�Ä/$n<"$��� ��s$���! i�~, �^ޑ��B�R��n�I&)U�n���� ����w�%����u����^��H�Э%��^T�K��w��7�޴��e����e�\�a�6`.��]m[&�(�I�(�����1$�Ǐ�i/n��ijH�q<Q��?fQ^�J�e��m�Z�栝�.Fn8vp�g%���E��U��46�M*�F��+q���Ԭ+��̳W3p+�'j�{����v�5����,\�[A�@4��Ҳ����o���0n���� ���d��4����S��k�*�K����K
� URR1=޴�������tw�,\҄m�:;1LH,I/n��i-[�I%��q��$-�q{7��F�/���牴�z��9�[Pߍ�E`��֒ݡ,Q���y_����mw�Q<U���"����ߧ��e�����-Yt�#�\�8m������tc���El��I-[�)	�a-����w��Jb��:3
�7"lo����z������!/-��I�ٛ�藐-\��"��娶j��I,�b�`�� 0 �mAK��S6�=�If���H��7���v�H�;�Ij�tl��`ۇ�I#*����׏�IrX�ntkkk"��&� 	���" n���� i��i�f^��p�I�bG�� R��U�β��&v�%,m�`Y��,bms�m�d#�&�����߽����(�_nm��G�O�RI���,��cAK(F\�b��v�lo>� N�!� ���� n���Fox�$��(	 6��m��m�{Ԓ�n%i$�������w��$�&X��D�!J��g_��O�������|,�c�Á����<�4<ن)4F� ����J�C�3D.�,
TJ� ��X0`F�$��)))++�!��ދ���Ȯ�����Pj@�C���K5Rh+ ��k���%OB�7�{���m�I	zBR��6C�Xy�HHB��h4�xQ*s�˶��m�%���
�RT�c+*DaL��;0*Ij�Z�
��	���Tq��F�h�*Q�tk2CA��M��RB�����5��6R%X0,Xـ�S2�(����#4'�̛�%�Ѭ�U�`6�`I��YN<C&��iM�7��<��ᎎ� 	��JHRS�e�qe����$�����Bi�o0����������s�s�s��]\���9�L9���W	���Ur�s��e���p9W9�s�ck��9�V���s�SmTr�b7Z��qa-��'Z3C����)��l���ZmT�:l�(5%�-R��6��I�;Xݥ�FĄ6t�J� eZ�#R�YGWk[�mՎ��.�)uڻ]4DQ�eд�2͊	+V�B�U�Y��i(a�V��ҭ5�u���[Iu��(9�6�)2ٝ�)m�h�,m3YZ��f[3Z[�U�R*5�rBقWi�j�ėka�F��Z�x��R)3/itUq]-�.Õ,��*�+B�[�Q�iL�/%!-.�Ֆ� V�j��v��ݫ2�٬�-��is�����A-�\�*T�:�M���7Q�c]���	�l��;�l@��)���#���4�
T�lXGj虺YM.
�\��%Q�&�vc*�5�f-Ep�f�-���T�.6�VZ������S]��\OLC�7Ke��|����:\<���Z�&#YSYA�rs�lK�;�iv�[�F�t�,�1k�M�gJ�f�J�:���+�L�ʘ���+-m�c\-Jԕ�A��l�/3`�˱fi���!1fc6�j\P���{@��;m�&�D%V[�6�+ĲaYf�u�7D�e�p�nk�2����V;�����jun�؍�n��;d�X�kY��I�Z�>����! }t)����Q>OP"�i1��q�Sj��|�{�`5v ��O���{�%" л �xH  h� ]�������	2��J�%����<�����eJ�[is�S!��-�D�t�%��qY����1$Tѷz�JT1�%�t*A��r��J|�Ij�j�5�m2RT麾���bU�Itc�_QKV�Ü�]"��yw���B��(Z�,Ъ���:��c� �W�<#��d^��'���r�r)���.0 �� �~���qd &�� 7=ÈG�4?�H�Pd %[�! >��ݶ�|������R"BBHII@����/�����9k�lծ�1�Q��*� �����6��j虻Z�M6�5P�J�Ң��.st`�.x�KCZ:�lYZ�kF:%��cK�fb/:	������b31�� j�l�$,s*��L]lK��8���\��R]�t��?�չ���Ǽ)dI�0"L�+��|v�������Q1y���anjL8�RUhcB���u���%� �_� o�Q��	{<_y��޺1sZ�
F˴v�Ԃ)��v�%���I-�.���8g� ��JT�v��O��TS�{w�DE)t��`�8�� �2�<4��۝��#�<5J�n
�H�l��~�F���'�o	 F�����O�."�x/)�\U���ۀ�RK#K�Eef��QZGx�|a|�!x��6�}� ��$�埛��Ɇ�M�f��A��Jmhl�_}����U_?{�;�IJ�ĺ��Дh4{����p���A�@d������ޤ���t]Ǝ�Mm��3Z׮ֺ�F2����Bʛ5nnA��u�I�f�ػ:�%��,E)m��[��9�Z2��!UWf�9[�LԤ԰�%��MQݐ�F�?�*�?��{�*���]�� �Ͻ� (�g��L�du�𵤵�y��^�ĩ!o�^/�%���F�7�{Na�з��p�w��0Nż$�\:�ޚu���:d��u�m���KrA�}E,�1-R+k����t�T�{�{	����W�"��$��g�^�_�rp�����j�բ͇j��L�)�13Y,�G���}<{�����uI-���������8��Ǵ�&
`4�T�lv��<�@��^L �s� 
9xs$6\�I,�1.�t�>Z!�ՒQ;ܓz��}���B�B�
$�+%��
�H��UBYRK-e���%��!�m�(�]�l���z����q!<b���;[*�b�;q�V��(y��۳:�pӖyeuT��~t?�����{�D��=tNd�,���FjZ�7&Z�Q��"�=�P2��Z7uά�r��n�%� i��JAFG�iݬ7��ua��r�����c�En����dTƛi��էP��t��y�Ӱ�}�;�^7�7��a )T�ä,���p$s�=�w|�l�-;�<o7ɨҘ�.%2��7�~ٹ'<�gۻ<F:q t�O=推>흅�\�xI
G��i�8�L��9'�Y'���d�p,���N;<k'�D�q�P9i�XM�%��Sˮ�d4qA�I%E"�H���n%3e��o\��w'����U�ğ�V#i�Grہet��g9�{��N���:���z����(}��7���U'B(�P>�Ն���-�t�P�~��|TK�XJګ�]5T�VI͞�d��bZ'���=�ج�ê�A�#N��TУ�>�N(�ι@�<��ѳd��v-,��j�c]���]P֬WPͰA����̫���fQ��v���4V5a[� �ܫ�u��5�Y��Yr�iR�ؒ�:5Վ���,]m�e��lR���r�[Hd�6�U����SJA���1���c�h6�T�%088+&����$�h*2�t�HL���ǛՂ$�`��ĩm�1e��A�̈́thq�H%���ݽr��ٝQ��K6eo��o(m�h����	�b��b�Z�Ϩ{�*sӪ�ӊ�o\����朂V;�u�ǎ��C-�VI�(l�'w\7���%����F%1�;Uy!2<�v������ ��p �J�VI��Z:q��6M:����G@��������<�� *{�d��K¸ѺBŃm��kݜP#1F���Y0b�����rJ�&Mkj�c9������BNJ.��Ah��-$������î�����e�Irhcm�S���k�LM
���Z��x-i�t�W,���`!0ت&�p�&s(ѻWfۨI�|�-�t�\�Y��	l*��&vƳt>��P}�P7sz���z��-;&J��T��Xj��@�c�TݜP=�P��:R�%��;�1�rV�g�%�T�O�?$wV�&4�dt�`P7ϹP>�Շ�fuA�Ǽ�xw5$$�R��c����oN�k��mV5p��cd���2��lֲ�骯ْ,$� �'�Ze�� �,������m�wt#�F���)4j�=��NA�$̭��D�������T|�|�v�4�Tm�0V�|��D �@"��!-�AH��PJ�j�,QaP� ��)_��}���ܓ����'r�+��0�x��7I��*VȻ'%C�D�����Õ[>$����d���Iв��(Ֆ�N�� Y�{�Dͨ}h���+'Án��a�W�E�-Hj�m��}�yPU6����f"Pk^u�u훀�Ĳ��xG�3�=�(�z�}h���we}`�A��&���Yn�iL�R$	D� T�ت]$�#�LʑY'�BOpu�61�G|�Kʊd�.۱t�:�͒s5�s� Q�y�l���|����/�~ȴ��0�e�%[�Y'~�]��s�u���E* t߾>�����P�w�X2~+r����C��5��D�@ǭ��'ÁM��d�6b߄Z���%@�^���/|� �F�5�S"��W4d"(6Ur�U�9���:I�T{��嚻n�v��#j�֭s�EL`�7�}�~�=tOv�VIܭ2�=����TJQ1+�+�(̠o�q�~ďk���9*x�$�k��SLU�KT�V��j�������Y'f��p��'���^�tf���K.�[��l�t|z]�ݓ�s���{��nLp�	���B �@���4-�湖�ح�i��r�mCD1s�j�g�*�k�ְ�l���G�]��Z�V9��Ԯ�3=RR٣]�%��t���\�q5sf`ڡ51��Դ01��a�0�u"ٵ�ƈ����j:�k�
�+v�"�(*m����9ۣ�t�����=�4��p�L&n���n�"�ٯ��.�����P���uk�����Y�u�-�kG4��翽?����{�,��S��rB�t�Wu| �`��M���#�R-֡�'���O)إ���'}_|����KD�jbxs���d�^�Y2���I�+���i�VI���~�p�p�����$��$��%���@�^1��T�5V���LŒ}����'��ˢ{�"�L�bZ8F!#�D�l��#m��h������|�����$�hl�>����+�_�*���D��E;��(%n��$��%�?���~cc5&a�������ݸ�2�Qn�a��@�_�� {�I��/�Y'%�Gt����aں�/������E��+$�I��	e���0��F���$�(�}��.�˛ې�;`a!6�6)$`E��f�MGB�!	! v����q��_�M5�q��l�4��zR�!�P�A4a�������<M!Ĕ+&�	�����.����ԯm�9��FB@dX�< ��$�3�n�h�9���Þp�C��@��/'56�!��������� �o�X�'�NͲ�5Q�Ƭ��ɚ-|4֔%H�'	g��u�$��,���3�g��&�,F$�	�:6�E0�lp�H!ZZJX������d�nv�Y5d�PgC����� ��I�����%� BD����ɛv3n��J��Y�����M�	xn�H]�"P=��JoT�L�ojhq,.�}LGL ze��L+\H{�u�'�r�mx�:d!,�#0ˇ�K`ىŕ�-����$��<��h>$�%���?.�
�*�b̬ԕ�ڂ��G
e[�*��V�%3c��2��%ʡ,�V�v�#�SE�wgAv	R�ld���]ķ���똪��k��.\I��C���;:ۋden�.ƃl�N�ͫ�;^�k6�uع�eu��n%��E�JИ6�uM�ݘg9�x�F��xD�Z2�s��2��l�5�P�,�XB�� �-�.-bX�emd,P��%�e�P���S&�ڪV�P�b�s �Z0��%t[���If����`X5cy����ԍ���Z�V�Xgg@�M��HMk*�vn�fcZ鵴�Z��*��xQ)��� YV��m�R�5 Z�,����t ͗M�ť&�0����vh��f:�#N�W�#�eYb��'�'I�E:�>T��:��x�(���瞞�V�i�-��j��qvYvY���e�[Y�(lE�Ͳ,/�{�K�1�An�Wī��[ab��� u&�mI��V���L�FgwF^��oy���Y��c�[
˙���BwO{���}���٩�h��ؽ�΢}��r����~jZ�+c�&F�כ�����$���]ܭ2��@�L'*�*cy`@�y�X}�;�����%���(��3��@��Rc�5Kh݉6�������$��]6��t|9����OFz�*��i�Վ������H���İl=�ӻNA�%���e�&�*�L�/P�v�
�MB�Z�ѩ�e�g�~�����}ı,O�h�ߨr&�X�'�h���"j%�?��_�<�O�O�~m�`��%v�qg�wh��ƞ���N��D�]��DȖ%��l�`r&D�,N����r%�`X�}���y"X���<uT�� :�G��]�#�@�,O{�w�CC��)`"B�qic#�	�c�0�6��HI�oi.�U(��p,O���v<������ϯp9 X�'��;���E������~����K�˒뚶��r"X6����Ӑuı>���
�`	`X�w�]����=���r@���ώ��5��.o�K�9���9ıT�<�]��DȖ%��tgݔ9Q,K���ND�,E,OsM{��x�~���F�O���y�36���%��~��"X6B�|�4%-�.��Q.��Cl�H��Wow���}�zw�F%�`}���hr�X�'}�;"X6�;��˩�ɭ���M�'&� kk�)�����'I�b�{>��D�l}�f��r�b{߻�9��,O>�f�Ȣ$A|������;�m9P,}���̳WVl�K�f��e�h�r%�`X�����,K��;ݏ j%�b}߻�6��`X�'�џv�"j������*�`���n�u��n�������� {g�m9ı,O=���09ơ�`T_P?ʉ"*A�D�$L����6k�A�%������D�l'�grgI-�Ȝֹrr��M�"X�E�����r&�X�'������Kı<�{��r%�`D ���wC�����^�v�q��V��@����������eB�W�٥�岎�eՍ����
X�M-��[��r{�������X6{��9 X�'��g{��`�{gm;{f�vr%͜�.�j�Mi3�f��n+2�h��|!����~�� �%���gyC�,��l�v�<�����~�f�:GHL~�6U��
�����tƮÑ,K���gݡ�*�%�b}�{����Kı=���r%�bX��Fw�9Q,z{�p�]��ț�9������aț�bX�{5�ݧ"X�%���>�ǐ5����9������`X�'����C�,�	�Ғ�S&�D޹�r�Yv<�Ȗ~F(����Z�`X�'��~��D�l�u�v� j%��7�fj�a�6�m���;jKRˮ�[��5T�M5�b4D�;9�M-�5e����*�b���@}c+�U��F�+��H�R\�!�5Σ�e٩L��иi�m)vpd��4���x�t�����,�SB��ۜ�uZ��1m,&��9�v��	�z�������r�c;>�u���{<9/|�>b��g�xr$�H��ъ��H�"8������e#T٠�+�4n6�g��p�qyݩrɣ��D��ߏ��9ı;٬��09ı,O>џv�"j%��}I��h]���Ϟ_��H�(�
a�d��պ3aȖ%�b_;�u��Kı;߶k;C�5ı=���m@șı=Ͽ~ͧ"X6�S���5�36r&��s9�d��"X6��y����
d�b}�Y�فȖ�bw�?~���X6}�z��ȟ�#���?~�\�Rl�K��˾l˒�9��,O{�;�� j%�`w߶wi�9ı/��]�D�l�~޳���%����s���[y���-��6<�`Y�QCQ>�fӐlĿv�����6��~�7�C�,K�{�ͧ"X�>�!�vMMh��D浛�h͙�.Ñ,K����]���D�ND���_2M�ˢ͡5u�	rѬ�l��cProEO=��wiȚ�`X�g~�m9İl���;C�2%��t�wn]l�Ng7�'Iu�V�-�k�cE\M�3-���)��3e�--@q�	�P��E�E[+�6�u,�(�˝CTl��a��&p-��¬��ku�t,��۔�c���>)�ı>���ݧ"X�%��~޻hr%�bX�g�;���
�������فȖ�����3Vf[�����9��4I����<��5���"���u��f"X6�߿o�����"ibz�:GDL�W�-�Vr'9��ָ]6�`�'}�z�����<�_N�9!����"��j'~ޯ�`r%�`X����Z��b#��/
��Վ������I����X�"�D�����r%�bX��w�7�C�,K��l�`r&D�?0"}����r%�c;�og�j]���kzќ���r%�`��4gݡ�:�cx��y����l����.x�������;����s����������߶wc���<�fw�9RD��}����������3�̷$bU�Ik0=�R�9{;�y5�y��,N���M� X���{;ݧ ��by��� r%�`X�w��{�9ı�}~���v�3�2Ys���9�,Kߵ���9� �"c �'�wz�Ȗ%�b{�џv�"j%�by����r'����ӢtN������m������{�iv��,K��������%�����r%���� j&�~�����K��>����C�u�ﻮ歹�Gc��v롴��n��G	����<��5���,Kߵ���9��?$Aȟ}���ǐ,Kg�O�]X��>=>O�"���X�'�k>�`r%�`Xo��n�Z�iJ��k+"ei��붹��/e�ֵ5����w���y"X6����"j�b{����r�a����sN�G�w[4��v��UBȀ��q�����8�''��v�"j%�`y�w�iȖ%�b}߻�p���DȖ%�����蜁��Ͼ��_��/g�%�"_6�����bX���xm9��5Pl����C�5ı?~�~��D�,K���͏ X�>���Ivr'9��z�����r&�X�'�����r&�X�'��;"X�T:�⟠ nD�~�����X6�h����: #�"$�W�UU��۷]��X)`��Aj�dOw�� dK��w�_�r@�,O~����,�ȟ}6gT�D�������4[��.m�2h�ֶ���%��~��P�K���=��|����D��6�#�к�-���n������ߦ~�S��`��h��m9q,K���ND�,|�}u�L3Y)��371.=��Ȏ��l�y�j�ӧ��y��M�"r%�by���9Q,K��ӆӑ,K��l�`r&D�,Os﮻�2%����I���9��5����WXl9��,O}�>�Ǔ�Q��MA�>��?P�@�,O����J�`�'���v<���T�L���C���捼�����]kZ-�r X�'~����,��>��jr�X6�h��NA���g�B���A�{�6t�t�+}��e޵�� j%����׻NDȖ%��~��"X�%�ﳻ5���,��`��I!# B��$dH2A$�@�B!Р�Hs���@ ��~Z��mR��V�i.(˖�TfH�*����rr�s�f�i��4�>�yL�6��p�@��[aL�kv5!�L]j+�s�S�Ii�v��S]A�j�ێ	,i��Q�	��,ZJ��8��Yv�5�+ԕ.�U�..ɳ ��:C��>��~�3?L��C�5�ﾤ�u-���D����]ͧ"X�%��{3���ɎD�Hi��"gZE�"�k�ZhRkk�6�+-�r�V����f^��wı<���09��,Oj���y����U6Jwΐ�]���Ýr�-�E�1+��?�	��8L� ��b~����C�,����ǐ5��=Ͼ��?�yP,K��ߵ�"X6��~��̓Rl�K�����eͧ j%�`{���c��
07"X�����C�lK�����N@���٣;���T��&G��B������ީ.��ӑ,K��;���D�,Kߴg{S�5ı;���6��`X�'������ҝ��k�֢����}[�>L�"dK���O߿~ׄD�,K�N�����bX������2%�� dO��5?P�L�c��%5�u��3����f��ND�l�����Lr$�w�7��R����k+L�c��:A�'K`������;����bX�g����,��1�X�H�#�O?Xt�_:@���8:O���b H��#	$kQ�	X���F(J�#- �FB$P�!I �N!��������vf��I�sZ.KDGf�u�)SKH�kk�F�݋�kG	�cs�nڣ��.�V6����Rh�ړ	v���e�f-&���3/h9�M�'w��Z����&��6�bw�g�فȖ�b{��u؜��,��xm9��,O��޻hr%�a哿[��5�e�ș�rk���3FӐ7��;��;��?� ���D�>����iȖ%�b|wFP�MD�,N���s�� r&G��3�CWVjl�No������ӑ,K���3�����%���o]-D�,K�u�ݧ"X6�|�{�9�<��Q^F�
���o��޷��A�,�@b��V1]D��?y��C�,���ǐ2%�`w﷩���,�UH��A�O����فȖ��{/��h��͜���d��d޵��D�l���6��`Yғ�7�>F;P���h�y�l����5�,6��w�������D�l�џv� j%�`w��m9���zY>3��3g"s���5�R�cM�Ơ0f�='I���'�C[ܻ�Ժ�yı,K��?~�Ț�bX��{���bX�'~��iȖ%�b{��5���,}/�d�̺�ș�oYɽ��JfÑ2%�by����C��,B��B�ĆF���&B0&(��ˁ�HE��8��a	"֥�Dem�-�Fc`�V`�J��b�HH�0a0	HZeɂ��x QO�� 7P,O�4{�ǐ5��?}�����6�b{�ϻ�A�DBW �>SIPl�����U�ӧc� Y�`�����hr�bX����s�,�#�2%�럿T�D�l߾���:Gj�y0�tS����շѳy�����A�
A��X�D�{�_�rA�,����NDȖ��u�ݧ"X��L��������K����m��T�ɳ�.��K9���r�bX�����9 X�����u��uu��*���X4J\Y���k���$���t$B���~�C蚃`X�������Kı=�Y��"X�?{S�_��<9<�_9a�\�������	M�czw�Jt�Jt�}��v��ı;��5���,K�~�f��@�DY$@_"dK��{�O�9"X�������]����y���Z�A����g{����+ 
� X��w�lyİl����9 X�'�k;���Kö�	zffl�Nk|�˭I��<�bX6���v���%�|�;��r%�� ��<�2�!�E��'��N�T�S5���r��c�h|
�1y,�	rB�'���2���jS��})@�a�c����&ÀB ��K_�	�%��� Ąc đh�e���-�(T*D�K`� JQ�kY�bF�tJFD6B!$u��0�-X3ЌCT3C�4ϼI�_�w��`BT�	�!)+V�+|Z��.�߀�%7�FB���0���>�Jn�� � �ow  &�e
V�ʸB��b��<0-�/�g>+|x @����˭� � =��f6ԧ�!�I��Ȱ�a&���t��C��e����	}u�h�i%$_X��}�i��m���-��ֵ�k�]4�%��ai
܆s���ܭr�s��&�k�ZֻlխkZ��ΘF)5)��<5�ZCd��,�*�̛�l�-Lٛ�����@���M�6����l�l�@6B-@��u�k-�GE�bm���3m#�Ll�e�60b��
A��n�-�5�&Iusbf�SG�����ˢ �Yj����cn٥6nі�F�.e��m�e:1v6�RW1�rLXٶ��-�X.�S"��)kv�R��l��\Õг7uk��a���6���ң�:��mM��[�֤CkL[TЖ�j�b����v�\̒�������KLiLE�(d�sWl�LX��Rو�t��3�4T�$-��R��T�1T���0B:�Bg6e�;K5L��;L[bXm������󴭰�elZ�m��AЫŵ�Q��]�cE��.3nٴc��\�ɶjT%���� �KT�4W,T0T�ے�D-��F[A�65�R���&ll����um&v���vb�De��`�M����q�vP!0��1���ūU�)�#Ca�ٲ�\ʆWb�0��JEc��v��Q�j�a/SL��5n� ���\��z)�f��R%��f������6�F���f[��]-���� �4fX�:��9�����7\XX�k,���R��)i�s2��S����$���Q߈�DM�|B��������D�D��Q6�U?*�@P��>���o]�9İl��?m9 X���d��h�g"]kz��oR�SaȖ�T(dN����C�2%�b{�F~�C�5ı<�]��r%�`��a����� :x�G��>6���6:x*�f����l9�,K��ݧ"X�1&�^��ܶ�bԦa��#�d���o5԰Dn�K�}����g=$D�l�F}���%�|�;��r"N$�{��B��3��ɷz`��H���i�ņ����;�详��Z��İl������ı>���mD�l�ާk�G�*'�7��>����i�:�c?�B[a�,t�>���Vi;���@G��^�jr�`����v���,KϾ޻hr%�bX����m@T�,g����������z�*�[�'�'NDK��{��"X�%���o]�9ı,N����C�,K��߷ٴ�K9���7�U���n�_4΋��	(����@��3����%���g�فȖ�bw�ٱ��ꁽA=-�%Z�-+�L�^�K�f�cf�t�C�b��2�fś�F�rЌ&���f�n�#I��"�d�Bհs����L��u���t�k&�sf-�УV�2d�K�j�k.	r�6Rp)�`-1�a��Ц\�<v��B»vH��h�
�k���D�	� }��5���,|��;��4]l�Nf��k��&��`�'}����xH��8�y��]q�����#2�Ls5�"���L6
>wӽ�v�X�'s��u�Ȗ�b{�w�ڜ�`�{N���3$ԛ|${�?��\�R����MZ�u�Q��7����6�`w�z��9ı,N��w�D�,K��g{S�5ı<�G{��@���;�j�g"s�޴S97saȖ�b{�vk�9"X6���ͧ"X�%����@�,K����� �9�}�?��q�ݞ����K�{'�&��'���6��bX�'�}�v��KC�2&D�������%���7�P�K��IMv��Ȝ��g5�֤͏ n%�`y��hr�X�'�}��C�,���vwc���<���r@���񓺙5�9|�55��2�ԛD�l�����!1ȓ�w<O-�tB˨�e��H�M��t�����ldN���?��NA�����xP�K��;���mN@�,~�}�s�&�Y��9�3�XDO��� ���y5�fd�V���կ�����3mwWl  �j��0�)m�e3���x+s4�)]]++�Iyf\mp�nкh���'�I'��[A�4��W"�k5� ��oU��؛�bX�w���ND�,K�����"j%�by��k�<���%�����"X�?�e韲Ɏ�O/|5�èvOLr'"r~���AP�%��޻hr%�`X�wG{��D�l��;��'�@p20��t���5����p�sw5�aȖ�b~�w�lyİl}��v���%���f�(r%�`X�g�;ڜ���=/���h�ݼ�����.��� ��)b}���9��,O}��]��ı<���DȖ%��{�ͧ"X�=����%�Ȝ��kWR�sSaȜ�bX�Ϯw�9Q,bK��,���FhYv�a��R[�AfD�����������Kı>�w���bX6�џv� ��K��;���k6r'5u��a�S��:����#�]}'"X6���w�@�K����hr�X�'�}��Q�,ľ���ǐ2%���]��p�j��k|0�3��i�:�bX����mB���H@V �h��"&���<��5؜��lK���v�������ȟ�Q2C��]5��[9[�^���]�"X�%�����9Q,K���v���~XdL����ߨr&��'��w�D�K/�L�뚒m��nNa��Fӑ,K �D�)�>����	���5�	b'�}�@�R@����ͧ"X�>_g�^�fi͜����d�7�ɰ�Mı,O=���C�,K��y��38]6+R�:��]*hGL����nj\֥��pDw����X6���;ݏ j%�`{�}�A�����������_'�5���h��]�_�+����'�ғ�%:{�w�ǐ5��>��붇 �%����Q�K��<���N@Ȗ=���[�۷�9��'.jL6���%��~޻hr%�`X��}��N@Ȗ���fӑ,K���w�NAQ�,}���w��.�D�l�y��]j�9Q,K�u���r&�X�'s��6��cM(�2&D���hr&�X��M���<�#��:D�$�(���s&s��kRl9��QϾ�ݏ dK�����`r@�,O;���C�,Ľ��ݏ dK���2͚$ͼ�w��s{�3z͇ �%��~��d��Iđ&�wx3K�]�b�،�+a�X��k5X�S� _��ϻS��`�߯{��@�,O���u�Ȗ���N��Lѳ�5����Cz
����bifMj�ֵnӐ9��>���m9ı,O}�}�ND�,Kϴgݨ(����%��{�]�ș�{;�d�L�ș��ɗY�j�9ı,K����DȖ%��o]�9��,O{�w�D�l����@TMD���emm�<$��K|���<':H��O���u�Ȗ�by�wc��`�}��6��`X�'��7�C�,,�v���MY�����'58ͧ n%���DQL����?m9 X6���~�9��,K���� X�pX�B,�`,c��[���YW�r�M�d&і�Yk?��x��(�8��sH]�n#��(Be�����m�*	P���%��lU�H��k3K������%��74�cj��c��玺*�m��\�b�[�][)]�̚3SH���v�������f�UA���"{����@�,{NߧunI�6r%��g3D���ı;���'�&'D��u�q�V)n�\V�Zb �մ�<q�дĴ�j��۝��j%�`w;��ӑ,K���g��D�,~�!N���������;�(
��̻�����ɦ�Z�6�`X�'��z��ș��<�_v�9İl>џv��r&�X�'��f��2%��})ܛ�WZ5��.��9�3Yv��bX�'��}�@�,�޻hr�bX��Y�s�,ľ�~�ǐ?�"&�d���� �_:@�{e��[���8�,K��;�09��,O}�z��%�`{�vwi�9ı<�Y�s�DzT^�E�<�zӡK��|����`y߶wi�9ı/��]�D�,K�{�v��Kı=����<�#ȧ��/0[V:x.�����ND�,K��ϻC�5İ~|k�Qe�\^en2�x�Ti�- 3$؞����������dK����nӑ,��߷ٱ�ǽ��ɩtd��@��u|����q�-�ܺ�E��T�ir��2��BKh����r�l�Ҋݩ�vZ�p��n[�ѫ��-�nB�[]+1X2�YZ�άJ���A��ڛ �S9��?��9�������,����ǐ5��<�NA�%�|����r%�a>>3o䢓�����~M��/�|$�JN�����m9��,O}�w��Ȗ�b_}��jr�X6���ݧ d9�}��E^�K��'��y<9���߷���bX�'���N��L�bX�}��v��bX�'�hϻC�5�0 O��V:x;�m�Wl�����C"g���[ND�l�������=���mA�,��3"{�y�فȖ����?f��ֳg"g7n�f����D�l�����rIN���ϟ��69fR6l��m���T�*��]��I���k���,��߷�ڜ�bX6o�z�:G(��2y���RM�<wV,Ά>F2�hZ����s�fÑ,���g��N@�,���͏"X%�|����C�l��[�@t�"8���y:h�i���ww�����kWaȖ%�`y�}۴�<@:�Akj��E�v�L�b]�;��r%�bX��]��N@Ȗ%��l�`r&A�����통&�D���&jMhѴ�K��>����DȖ%��u�w09��!S"dO{���ND�,K��޿Z�bX�N�fve3M���s5�ssz�A�����xP�K��;߷ٱ���<���9P,��3ﳿ������ �<~�H�	V:x:��:�I��yQ,�~�ݧ �×\2�����˷	L�Ԧo�kR�%-51{Ͼ����~9q$N���v� dK���wi�:�c�=��Q^�M�|�y{�e��14��f˰{��K�3�>):�X�w�붇"X�%�|��{C�5ı<����Kı>�w���bX�a��M[.�D��9u��sWaȚ�bX��~���"�2%���v~�r&D�l~��~��9ı=�[�@t�"8���A"�����
�l�s3Z���D�l=џv� ��by�D��|+j0�,����)B--���UBZ���Җ�ĂFX�B"���	B�*�T�F@RQ$%���iF#,*��iKmv���W�D�D����6<�bX6}�����dy��,*�t�.��g3z�aȖ�b}��]�9İl>��v���%�}�>��9��,N���v"dK���/Lə�g"f��Y��f����ND�,O}�}�ND��:R7���5�0�JcK���#��R`Ԗ˭��zt��Ԃ/~�u?P�&D�,O�h�ߨr&�X�'�k�ݧ"X�>��3��l�M�|��6�Y�Ds�Yy�%����=��9q$z߿�<'1"%�緽�Ȗ�b}��b�~R��2%�`}�Fw�A����m�����\�#b���ȓ�"'}�f��2%�`y�vwi�9ı=��붇"X6����D�Q�2&G�����5��5��9�,�Nd.Ǒ5ı=��l��o]�9��,K�>�D�K��߻�iȖ%�oe�w-�j͜�w����%�aȖ%�ʃE�����៿�r�X�%�o��ӑ5��;����r%�`w�D�ߙ����Z��Uu�)�WTV%j҆��j������S6�ݠ�HKV��(��fk[+R��Mj.����6�ۂ�P:��1;l��+SY�,��s�v���P�%�a��@��K�3n�nc�q�J�l#B�S2�U��:v�O	ﻳ]�șǷ�I�t��6r'9�kE3�w6�bX�'}�xm9ı,?� �NN\%�d�0ԓZՅ�m��h�v0l��[��K��b �ޙ����5ı=�Fw�A���gxP�K�Ͼ,�`��#���}��>rX����n�3��Z�n۳�t�Iē��ϻ��`X�'��w�D�l����@�K���{ݧ ��{>���l��xry��<�����ȓ�#�~ٮ��US�5 �}ݟ����,K�߿k�D�lϴgݩ��c������W[y��e���V�9Q,K���ND�,K�����"j(!�b)�2'�k;�09ı,O߿~��K�y��wY5��g"]����ZkaȚ�g�@ȟk響P�@�,O�w?p�Ȗ�b{��;���b(�1�}���p��=��R��*��<}��FՅB��K��<��;���`�� �y�<�Y��]6L�l��xqX�F��S32��a8�����}P,K�{��C�,��=��jr�X�>��/]f�6��U~!"w]
�F*@�!HĄL��!S1�`Sa�t�HB P�f�T��V @$�:c	�c,$,@��)�2��"FF0��+K"�	ra���&T����2��Y�3.#��14Ё	���HH�_�����eU�Z� �Ե5TX�c�U5-r�hUl�k��[p��9&җ:P��֍�\)��2�E��׶��1�F�9�eK6�L��K�r99t��LX	�+z�,fZʎ�]�Z]�Zl�c�)� t#A�X�K�vck2��4�"��u��YH �q�m�r�Um�5�15��ՌL��KYl��fv�H���@Εݜ¶�����3�gm��U�ڀ���ҹ�k�`ݥu��de��p�,K5m�]��ic3���u�m��(ʹU��d&��Z�p�	U�k6�G0mk��R�G��tqƬ�˖��K)�7�0"l�Q��7"F�۔�73���f��5���l�ԪS73)�f�!�
mGgb���9h�Ex�(��bu�z"m x� v��|�g�s�],��R���pk��6�U���ws`[	3��QB�bR.�z��R�F�n*ۜEeA!fz\��Kmc ��3�#�e��ۢ�]f�]O �%��gxP�K��=�F}ڜ���%��{3��	�Eț�bX����ND�,~/��?��6r'5�&rs3s6���%��l�`r&D�,N����r%�bX�}ݚ�DȖ��}3��ȟ�$��������Ų\�Ȝ�37�y���aȖ�bw;?lyQ,ϴgݡ�:�bX��s�(r%�`Y��bz�:@g�O��*M�Wΐ-�W�5���Ӑu��R��GQ?��?�(r%�`X����S�5��=����&@�,N���A�,<���kkO�O��W�}���:��<Ϧw�9Q,7ɾXLɺCXY����c�"�v�ˣj�h�	���ޛND�,K��w���Kı<�F}ڜ���=�>��h�4�xrv����|/-FLnfs���DCZپ�M��l������r&�X6��ϻC�5ı;���9ı,O}�ݻ@�,g��e;a�&�D���Nj��6�Ȗ%��{�n@�4=:�m��dY"���S ��RDrA����ڡ�x��"���bw�7�m9��,Os���ǐ5��=���mA�,|�N�t���g"k���]��2�Ñ,���wc��`�w��mA�T,Kﵟw09��,Osٝ�N@�K��ta;�
�t��}l$�j�:GKv���qi�Շ{�����%ˣM�\�*sj��l�$1e�rbx�'�d,�KC��DM5��	U�p͞�$��=�d�b��8���_[�
:z\�e�f\��Rn�*�+$�a���p�'2�/s���.;�������"1R[Tm�%�� H��=tN�?$�͕d��PT��s
���ݽr��{ʟv��	O�H�H�V�"��2(�!�@*�U#W�U��T���s�������Q�J��b�%b��vO��ʆz�o�b�=��~� ,�}�4�vІ:����#T/o:,��Q�lV�eJ��n{6�0�O�RA4Uf`�(���I�k������l����$�y�ǖt��T�Y��hh-v�{���P��"�OV��ps��lc֎����.[,i�Q~T-�t�P<�oV�쿀�pp���y/���V�;e��]��:��J��uA�<ެ��õ�Tm7b���;'À ��ǭ�^>�N-���󃃝�}T�j�Ti��[r�%�i��5�0�ku��2Ԍi�4adru�Ŷ�얋M�ket�WbmV�T���2�*��X��i���U�Q�#]c[�"ʻ�QM�jB�-,ٗ:�i]msm]�SG\�v�F!hh��-�9`ׇs���~�}���E��̉�X���v����݊ԙ���H�`��H�P����i-�wg��ں�>����R�Ptn������ �
��Y[IY��I;g��G��C�]{6;$��%�{�6]N-�e�Uv�J�]��N�Ŀs���#�O�tM[�΁��C>�o�#�W]U5��X{zP;�3����`}�҆��~�5��[�+���O�99���}��^���;#�8��#���S����W*j8���r��j�Fcțȩ�9ʙ�䎪u�km-%J���"$�#�N�bZ=AR��h��81H, � "E"�BB,��`�!��>B�3d��WQ��k\L��%]\K����j̀�V[71H�mv�YknR	�MD����P5�vTٚ�K3(��e�Z��̙��R�V'�� � ! � B���<Ֆ�9��LM�aV	J���w���&f�-ܡ�� u��{�d�A3ğ#Uwt��V�j�8����9�4b��O�ޱd��i��B���m�iݪ�7���:���oW�������=��
�mh᰹?��H���e�vG�d�Zv]�8��z��j�N�#��ev��S��ٝPd�X��v�\�k��#.ZK�Yl͐�aS/�9�;���"sg�Y'�Ceџ���пy���Q�\�fM�F�DI�,��(/Շ�v����r�����"s�v�FF��'�����P6 DDڧPgӾ�d��ǭ�5KG9%�F�S��I�dY'�Ce�=�.�89ĳ���'�N���$qͩṳVcM+C{�� �[Շ���ý�r��xF�������<���[�ca-k���k��]�GFѺ&�&�T�U/s�sw���O�^>�Ov�ˣ��'֒�%�_���<v�Xbf.牉<�&(����VY������7�>��̈y0�����m�3e������։�y}h=��3�.c��xL��6�9������=��}7>�{d�3����E�@�@�B1 �QL]�9� �]>ۢ|������!5L��[WWJ�$œ�
T3�D���36X�}�s�,�'��^�J�*���)R�
�X��mr(ҒG�E�$�L&�:�f[�z@��嵨�������ę�'��ɬKG��
f�)�ݙ�[����K��*��&�����>����wz�˷�V�Ր¢BQ%n��T�RVI�V����> r��<��O��X�Ov�VNP;P 	��2��-ݙ�/o:~�A��:�Cﮉ���+&n���*e]���U�ui�tN�l�ܭ�ɾs���I'�ȃ�j��b����KP��a�P��R�4�Y�mq�#bWF�9e�Gg*�ٙ�u��\@��X�a�D/X(x�ͷ4v&m��f�B��%m�U�*T+e�Q�!c��b�k�2��p��r�z����6��QtZ	>�9���� �׭KGwBQ��b��d�8�@�_r�d�+ba{B��l�\(�ԋq5��:d�j��|8>��b&{�>�N��t8<��}�'K2��QcRc2O�<#M���B&��"���g-ޫ$�ӳ�9�β}���#'���m�U�n��a�Ud��[/Ã�|�@�?����$����d��Ĵw�(�uEںvRUO��o:��z��l���Άo�`e�Fʣb�M����A�}=ߍ�o?��T�[Ն����B[���b�ً�>���u�99^x�8x�勭ZL���
D�]�P+�DЪ|?� y��}����{�U�{�$�;���X7j��!��� S��ڴ5y�cl��k�fV���i��J�`�҄���5��gl��W�M��Jd5ю��"�qf-BN��e]m�KKH�ٴ�����@���@զ�a����}ʇ�# 4�mڷwH�4SVI��� ps���g߫���3��~�L�bZ2m@�4�s-QZ���y�*�gy��-�t;˹)?D;-���Ȩ{��pʒ��]v}�Nn�l����G7{�s	c�� ��3�o������d.��$��2��"@��{���k�TݜP�;GѬs�j��&cXJ�s+e��W���:C���)����������$�(ItI�����,ܹ�oZ�35���y�{>�UZ�x8I���3u�h��$���[�'⾢D�NQ�1�J����
���V�:{�>�<�w�\B�n���ps��?�~����?��95�d���({����R#,�6�������o��۫��<d@���,c�!bf%�{�x{gy��f����+-�u89����9��'��/�=�~6I�%�'�#�NMp�#5h��<�d��q������fuA�y%�9�"��¨I���e�j��*��S[�{�v~ݓ�g�]�.�@��D�R51H���`ē��]o!0":���DܰD�$RA49Pk�̡�L6�D�Ga��	X��"�P-"�k5�5#1�CC�A$IE6I�R�*R9A��$HD
FE���������-HKŅ1��p�d��0�FX��)��P���a3	LM@��d�R0�B��v�����c � P�5�LO0��k+� ��#�lְ�3.,q�13P��ap�l ��Ȧ��.�$����/I�%�K8�,���a&pƘ�ᤍIFYM2ã,�hk�Û�{BKЮ�й�[l�gƌ�������vsc��0��M�K�*@��o5L�s7�H����H�-_/�p�M�y�։	pb>v�{��̒�'LI�%$������r�r�b�]\���9΋l�3r�9b�k�k\���9��Cg39W*�9�\ck��9�--k��f3s63M6Kj���;V�XC0)j�v�mjɭnB�b�݆�զ�J7H�Fذ[�v��u{mĹՍZ��2�T�ͭ�.���H��[��`��+l�&
:�WX`�U׬���m�:ն�\<�������]qp�U^%Ycv���iEڎa�
⎛p�3r��֔�,tĽ�%%��H#Amq]���{���a�Dj�n��5�s	m%��W�v ����Flm[v�*��6�34ś��DЖ�diL2�
,�fՍ�^�.ah��Rͬ9�f��q�����iWZ��6��^�ih�t�jj.]3��0F�(M���R�LiUkmI��B�ŀ��j�,�ݜ�ks]l�.��hc`54�U�P��7f&e�님�Z�\��6;b��F��v�ֱ��R7ڽvtu���.���
�R�Իs�Ҭ������v2�/f�Ze�V[�*R�Ix�h.M6�]�ZYZ�:��ֺ�uьZMrR]�f.�l8-��16��;�n�y
R�xb�6��.�u�4����2J$)Mf5�E���W2�j�n���vi�c�#v��cvenn3̕�m���Wm��tD`��r��%�&��n�n2V�݈�	�0R�F�����gt��$���"|�/�A���"�$x"'|TT�P҃�OA(!�m@v��U�=Q�g u]�b�3hIt{�H�b�][	V��?'@�l�����l������;�����\EM����I��y��0t����!{Fԏ��$�G��٠o�P}�N��E�.fA+e���2GLe�S��l�z#��|����ݠ{�K�rl��D��a����.���`�m3vL�p�� >�'��͡���wz��;i8+#�*Ӓ��kL�NelV~K=Bz蓑{�GwJT��",mWc�5�v�(s��÷��x'Iӻ�>�e�%�a��M�(STʸƍU�gQ��Cd�wc�����5f�SU�i�l�<�7�����\A���ie�����Z��`a͎�2�7as���ݵkm����!��x�@��X-����;cZ.�����ȹ%�2�i`.�g������_K�Q�;�2���a�޹@�ԓk�����V�gEM���M��b��swa�D�W��2�VH�����sU�����L�[�[?
D(Gs��}�z��w�P>�P>���Ϗn��2Jӵ	���$͡��ƎJ��3g�Y'�P�Do�vA�v��26���}ʁ�=%��9��;��OLE-8�]�1I+�d���
�c�]'��d��6]�y�Y�i���;cW*�y2���r������m�К#f�[���L<�%�&��c������k�T���o'Ѧ���by��~�`3�`�H�hT�ry/�楁�����e�Z�X�&���&��.�VhԽ�-۶�:�ųΰ^�͘h�nwR�FG���8."�<-��wI�:w{罾�"怑�0��I&�\Ee��û��P>��y��ps�������W��)$ٻM]�4j���ެ7��({�����5ڿ��pȁ�e��G�J�����P���v�(v����Ho���)[p�����V�:��z��1v��(w�y�#y!�m
����zuA���/x��Zč42�ַGk��NB7&8����rk�T^���H�}��r�J~dN#Y1� LD��	�T��z��D�T3��9���l���~�&x/��j���ѹ��ѫ�{��=���E"0HDH�*"I���&�_�ݬ7ώ���NFDZ��"x�dR�;5�g����Y'v����(�����p���N�ջ΁��ެ7�8�}�P��5�8��$��������?��:2����[mci�����˩.fݠ<�q���{��L[��\6H��U(%������z%J�+-�4��UPm�I̡�蘰�tN��_ppu��Vf��	��*��n��(z8o�(g���^>�OelVOp�LP�%��i�Sݳ���(g�ߗ������uf�۝�)m������p,�yY&l~6I�F%�z�eY:h���A*�%M�nK�zuA���p��Y[�d� ң�DK�0mb�^��π���ݻ��?)�D֝[�NI��yc�5,�f��!��r��n7�>~?���=:��^�{�8��Աs"�DWlZp��w���a�=:�qd�~ %�*�j�`۪v�U:mX��?���*����|����)��ݓb��VO��9�-�~6I͌�윾��nN/U4�XF"���)���G6O<���a����W[]�2i]]:��M�^؛S.sֵʶ7i����j]�k�啫,F��Mne7,�ۂ�+6mX�1�Klr��e9�8n65q
��m���b�� ��hE2�hJjK#QBɮ�[�E
�0��R�kV����N�t��'���ՙ���#��َd�����|y���mK&��$#lbڢ�j�
�Si���x�'w����������a��["�V�orj`���ˣ��n�������P�G�s5��9���N{�z�@R�f��wT��Dd��d��9��l��}�NMp�s�CJI��)%B��{��Y'�n����Jei�����pjdIDݭ�eJBc�}�3������΁�l⇽�y���J����*v�(�����x�3�ŋ-�j�y�8q[��߽���7ϹP<���w���mH[l>� $�HI�h�4$)T��H��E^�Ȩ�C\��beуή�l�
b�L��5��ne.�#.�-�M�H�Y-��!�b�&5ö%��J����* XVn�i�3`�c�b�C��G�o�gT�u���:��i�Y�]�<�C��)r��E@��q@���X{��P;�qC7{��9�[o���%����@�=:�� [��Z'v?'7i%B�5WJ�U�+G��88����'��$�k��>^7�7<����(�Ț�wN<ٰ� �1R��;gkWm�6�A��q�|�i��J��6m�t^��{w1;\����(j���L`j�,l������P>���M����·�g-h�Dow6f��5�]�<�O~��R�T��(wN(y�ug��A�(O��-BrI(�WT���wg��uGټ��x�b�$+bv��ws�{�q@��X{�8����c���d��rH��M��?ʵR��9ab�X\L�^��a�-4��IXI��R�9�Ĵa݄��e��ϏC04�:�0�M��[r�_����@���P>ZwV.;�v�ꏵ-曐�))*i�I-{gI�KIŧe�8��~��>��L,�UG?4P7zg�A���nfL�0�@��D2X�1XEB���b�B,B#I�4��"�lD #���7$��>��{=��ȂU�J����ݳ������{ʁ��r��xY��2��
H8Z^;� 4����"����5�Y@f
Kr[h����fuA����.`� ��:Q\F"����e�4�u�pπ��������a��������I��Ls���T���?~H��V����;�8����>��V�U#J:�����޹@�v��>\wVf�����ܭ0Q;����a�|uA��r��c�6��5AvܫIy�3(�ܒ�biFX�����4JT�!e�15Yn��+3�kK��i*���a-�5#6Y��aƓ���-���s)���R�(�4΅�6%�!�jV\�ڸ ����ݝ]K�R�Ƃ�$��������y�>�I,���Ln��l�$C��=�4��]���M��a�F�j�h*�n����ݨe�{$�C=���smp��$��&(�'��Lq���1�+�Շ�g/Շ����9	vw���%`52���a�㺰�l��=�C�a��Mڬ�'2����P>�T.;��P�����v���cJ���z�����w���ugݭ�m�k�u	*��{ʁ�,|��%%���,��g--�d����TK$�O74�D�Ib�=SeY;�E\t�MU۳�0Ը8�� ^�L�h%�	�50��� � �IP��0%e+��d�c��oS	Hp�\'�+���%�W8&h��a!�@�T+	�ʅi�%apj!H$�X��Z@�0���A&M!�Z�M��l6q�"U��P�
�
&I�BcF$��L
Uu��m4��Rd!�]�@�#$(Da$���4P�#�Z������uIZ"a�I>�B��BTÁ10 ��l��$�M'N�~���mAUU�a
�-���Uظs]UUBګ����MYZ���p5�i��l��j�Yn�!�k�K��� �d�U�K��jDx�(��0���aau�-�ٖ6��qR�˩�����en��A.P�͛A����/H��Z�j��[v��� �-�J��PaR�
d9t�4��ku�\��[v���J�m���v�kV����t��ج�`�mV���]��%��6��,��n
�Wi�F��R�P�-[�6�k��:��׬���K��Ai��]tq�Vc�h�p�mn�&++U)�Jj�XU��kX��]7���B�m�B�-ڈm�ֻ��#�����i{K6�β���� ��Bb��{q�JJM�K��Z�M�̚�8|��)�P�@*�B�¾��od�>ifu/;V30�Έ*Ʊ6h��#�L�r�eu�������
�F�M V�����k+V��J�%M�u�6��֪oޝ�~t�i���	K��m($�k�:(*��'61-�$����ûz�ލ�HK]	[P�����Xo�gT��T^7����-�i'�ȍLu7,q��<����M��{g/o:��r���RC�\#u�v����*��ua�ٝQ��gq��!d�A(�Ղ;�E�^��2�J�ᴲ[01��
?�(G�wv|-�t�d�:DKL�Mj����ye��˩&�B�.4]�[ �����N�;.��%�u������h���}|���r��?Y�̝����$#��!%Ua��RDY$ �R�T�Xa
8 �y�{�ܓ�����>��i�c��hYlqԣ�:�Ն��(^�t/ՙ�Zس�8�$�529({g]����߳�ݙ�՟��g�y ���[�m����t��[���a�V��;�F�RҲ爸ylIf�~����r�s�ol��-䛐�)(��eq��7��2��l̏�y{y�;��({fuA���Cp���b�n�c�mLn���oV/o:ݳ:��ώ���9r �]r������y|�}�诌R#`V�$������;�{���5�b�k�xQ�ya���?/>���;�c։̡����O;&o�>�J��VJ
cQJ��<ެ �V".���r��\��av`WQ�?ăq"߻��>���-����}SG0�wY����]XX7[PưNdMH���r���.�>^�t�LꏃR��7(�R���J�=ݎ��s�$sяZ'6���8��d��������:����T���^�V}�^�zŒwiE�GNh1��"ܲ�%G1���uA������7ww{����iB�6�.5E��\˴?�J�� &k��̖�4i�Vm+���тtca����k�9e릠2�T���-P���][L����vM�f��b�iQTۃim1aj�ֹW56ĽY���顦�����u����5�b����h��9�����
�Քȫd�U�~ q�4;�8r#lM4Hky�&��jݬ>j�h+�R�@�����D�ղ�Y���|�ϧ����`���h�v��@k��q
(I��5�����}�r���ެ�{�%v'^V�jc%����㺰��ް;��P�y.�NV��xVLj�=�X}��(y����{�To�k�cb��H�R1,�}�7�ܻ������?g�V��"��[�����-�N�2_����l���:��eeԚ��mis �j�i�����ߺ��.�ý�r��oF��8��EV����K�	(V��X�2>��:��f�͝4a�Z䭰�2լI�[mYX�f�1l��9n��)�Vh1t,�8p�g[-��
h]�%�F�i����t����C9¤IdF#c"q�rz����z��y�Xyw���w�'�wn����Vn������z�~���[�	^�6�@��Ӫ�'�=b�}�j��ں��޹Csس����b�bV����V�P>^7�,��9.2b��p�"6�Tu{�hv�Izg���[��S@��l��,w�Ͽ~������]Q���3�	��j���	���b\�L�ЗQT_`���������V�P�kY�StP��j�h�'�Ce�<��s�
ݲ��lA E�`B5	d
$�\"��H8A*H��p��A$d B4L��zX�K��#�Хj�e<L0G	B��GZB@JB6�b.�C��kW�rO/{�@7�z�;�^5�����T�#��r��tN��Z� %==b�9+�VL;�,}��:�Y[�m��=�3�����<ެ7��P�y$���-�V�8I@��z�ɍJ�F(p��S&㫥qa	��N6�E6���n��{q�*��uFỜ��ݪ���-�1[3*U�1+6�:����j�X{�gTy�*��Ș,��U1�{�:����@��z��l��xZr1�v��
X�}�z��w\�ř�3�f��T� d���F1�k �Ơ���$*#�*�Y��s�T�ӥf�9�N~��bUM�N��8V�U�qC=tN͗F�>]��}���I��kR9
ý����om���J�-��nڻa������
�R���~���ߗua��C�9vv5�R~y^%�3��dͣ�t�mu6:߯���5�h���^�8 D��=tD����NZ��6�Ɗ�o;���㿣���P>�= x���1�vؐ�;�Z��@�^�}ώu��fuFwi�����Udy`��=�@���:��~�	9o{��R;AeZ������qu�;f�M5)L1��&s[
�Ҭ�+T�.�؎n6��F�0���Ͱ��6t����փz�sv�\��HB��s�Q�[TMjGf-��nu�g�;J�@��j�*b�kl���v,����LW^�I$��{�i��%�;9�v�X�:�Ǽ�ij�:f\�9�[�fvZ+���Cm1E���&���ޜ{g�����	D�NA6�26�)�&��L0#dlL��2P=�3�����=�@�ެ��K��&Gdu6хqA�΁�l�����`}�҆��&&�+NX�8�n��=:���stv����z�uq�~����fL���7��(y����:��<{z4�m̒�������~��OL�(�C�A��L�<0X�dM�ɑ�q�����}���=�����]��2�WF4��Z�]3tYlY�V�K-�Ip������5��Ya`m?���m<�]�
=���u8�ю��0�B�u�B�,Kb�E���i��#*�jTm�s�n1Lq�������{ʁ��Y@�ώ����G5���J,E}ӊۏ7��ޔ�g;سW)!�c�)@��rtv����z���yPӒ�t"��%�8Ҩ>^�����}ӊ��z�ݩ�������s"���l�2G��c���X2j��eC�1�6�n�N,v����=�3�7۬��6�<�x�6��ض�u&�x5�Lb�7`}缨��A�ȥ�{��Y#qJ�0��j톙b�y�{�����2HI�xi@,�E%�;��d��p��s�%��%G����v1�Ԡo�O⁺�z���7���
�o,������s$���zuA�{ʁ�hެ�oVn���q�����P>�P1~q�4��n�Ы\�[-J�#��a2��wtn�(�7�4���S@g[��$�f|��;�ql�ᨥTG3��`������~�P}�T�ܨ|g�s�9����E�}�z����P>�P����� ���Kt�Z�uf��J��L�{y'=�߷��)#�e!H� �BU��"D����C`AЎ��Ȅ @��e�$CF��]$dp$�� J�4��p!II7 B�(2�#Рm���I0�(m*�	���(�$��JȖ�����!�]��b:�vx�������v�H�X�A)��$��BB$&�	�-[_%4��܄���$�+%!f�R&�#I#`�DVk~�f`���H`�H��xB�,�
�.>i�DtlA�Pb�!,A!����#��d� P�}��U�j�m����[mkZֵ�L�=��
��;K��)�mkZ�f��[nPkZֳ�V��\����s�.T-�t5$q����=�����mH�Ԫ�R�1b��f,��\t�Q�ʊ���F]��s@��6��&W,
F�\����-��[�8��4�e��Z�jjmk�ڜM�x@eמ���ޖ� �mYn�U���4Ii��Zl�4l}������&J��kp@�b��5�-*-�-��Yj��uNY�6�S�fk[!��8Yk&fQ�La3W)n5���m!2n��v	�38�˜��^�)3�-��	���Xh�m�R#I����/kۍu���J�G�G�,v��A���-j��r�ñhCSfˬ�b;04[tb�S�B3L�]��n��8 ��g.&5D�%�k���t!H[�[�+����5�]�
&�(�fƱ�bmZX�42B���+vc�fU�m�*�U��0�kX�	Mی\��ҕcc]wF��,-x�5R]f-�4�Ƥ����E5͕զئu�3J�k��E��i��ܘ�����v5ٖ��-]�\���.p�iZ��`�n�j�lҕa��Tu���F�e���hGh.���LW��f�MEkm���-��������w-nV�Q�
�z鞵�]�%ftp[�[I\�4fJ2�K�e5����ɭg ꊇ��Q4	� Q:`��P�Q�D8�/ʃ�x
Qv��*DV*��ߛ�rO>�g�G��HأV[u��Xo�r�}�Ձ����ݳ� waߔr��:��= �����%��v�5"�b�[z�3srC��m��	��v�@>��X}�7�3}�$q2\�oz�ὰ�GA���!���<n1��k�?������*��]Q��& �#�ą�����l����}寬{�3�������jYXc�>כՆ��
��� �u�F�Ib��qc��4�Xs9u@}�z��l�dQ���Ku3����Tt�7&�����#5J�-nj��&�����d�u�P��.UPG�lMU�là�2W\/j�t�F��ĸ��&Ћ�]�����֪Lؕ��u:s����k�WbX!��ż&\�Bk��*����/���ӡߌ=�	D�pk�%�5h{ώ�?��;�=�>���3�X����a�*�TB��d��'�$�P�����Q�\�C�v*J'�#Ib/a�+/3������=����Ӫ��΁�ܺ�s�vD5!Z�VPt�#V��e��9�8���wk�����C��:Oѵ:��1ܒ:�}���}�P�����8��i8��U\��&�t^����ꃻz��^;�>��v(����^8�ʀ�ޔTd	&��ᑨ��j�X1�b���fV����{�7�pT{�>�ؗ'ɬ
�Mp��1�"Bz���r�y��i0.��L�Nc-\�[����b�b��Z��-IMf���iQf�-��]*����
�6�T�zt�wO��|>@,�|ˌ(%W�y]k�a����T�o:/rꃷfuF�-91��NĦP=�Շ�����ޔ���f���a\u7����� �˺��>:��3y��jk"LJ�#U�9�V�3���{wV^;�>�k��8Ү;\�G�k�T����-�^12��".D���C�c�ҋ�����3��]ՙ������2[%?\�X��ѹ�H�O��d�%�(Z�o:��&n�>���O����@�6�u&�zə�[�y|�}��'�(@ ,@G�u$����9�{ʁ�������w��9��ԴQ��A�����/Շ����=��Cp��R�N����-RaՓ� �/��9�^�Y'.�պ���
�U&	B�Z5\��}����dN�Y���S;j�1C�.����J�����w&����J�OT2]"j �S���&��{ulY�٪����KV�9�;$���d��Q9�:������<�3#i�c�5n�~���rT�L���D�#��8){�G���F���&8���_���a��k�P" X���\���:��(w$����E#����5��LZ}�wkL�}� �ݗ�v���q�RT��Ɗ���Pn崬-;�j:ҵ�MP���Y2W$Z�>���?���=�N(qۃ�JdT�g�|db�
�t�z�nե����?$���=�RW�� :�վ�Y<���e��wf��Lղs5�~����D�ǭՒU���#hU�VS��v����uAݽr�ݳ��霚C�Da�5hy{�О�}�n����vmH����޳v�mf��m�U�o1�.��U[�ڱ�W5������\�1n�H����V6��b�yK���Y�e֥�G!�7jٙ���q-�K-��\J���������m���������6䉗5��mƷ+���$Z�GF�l��G8G��d�ͣ'AյwUH\AP|�ެ!�nA�����䎵�l���ìɬ��U����y�v������r�Ȇ�+�����Ec��A�+c�Z�X�ƚ�wN(xy�Xy{��5{WT{��#����Y��"�=흅��P|�ެ>]��q���q&�,C�cM��^7����P>�<ެ�Pk��q���[1ǒP;�Ih���-��d���qg�c֎r�U����S�C�ڴ��Pm��F��Z�[�q�:�ʎ�E/�B�p��I��2x���.�ɲœ�os�2~v�ST���dfL�+�n�)�sę�i���a��Z�i��H:���q���Z�jb����.��)-�c�M�qq^�wwI�F�Y3M-A0�m��sP�EA�y��a���@��]Py{WTx�����ց�Vc�}��(/Ձ�wJݛ8����gd��Q��2@������N(�y�Xyx���|�4�J�`�dD�`y{WT罊��w\�|�ެ��7��F5(�L��+�7�P���L���#�&���v����,G�,q�xެ7�Pwt⇎�M�ψ���nx-b�6��DbJF6�C��ua�������zvT{��X'?7Z�*�H���������Rn}y>��O}>��`yxެ�3t|�(ң�527Pt�Œq�]| 	j��]���Åj\�b�$�ī��/j�>���r���uf����1��,��(^7��#bx��I�1H��GmQ�ķT,�6�i�{N���b�z�t䃱�7
���3�4]]�,��KZh��L�p�'7X��ź���60���X���Gm�Y���n�{=4�yx�<�oVi���G(������P=�M��W�����0�?�H
J 0�{���y��o!�oI��*��$��+����襢z����� qO	~6O��5����W���(^7�!bɏ cm�f��j�`�3`�ݵ���L �#$�i'�i�tN,2]wLFDf���ޱ�Q҃Y�.�����H&P=缨�WeA�w\�|�y��Չ�"�TeM�8���%�Nf�d�Xv]$p�=�3yo1�Ec�J����}�:��ٙ�n��Tם����-Θ8�Yc�(�6I�͕d��;.��5�d�s���A"��kI��/����n�L2�6�.6�U���p�슸 �Y�6�X3k[0q��&�����Mb"`�V��`�4��M\^�K��!K�R��[)z�:%L�ZY�FW.��R��GM���֌9����x4k���b8Z����t���s�o~��ۡ��oq�\��,N�M����D64"������A��� %���g�}���oV��?~��5��7��ca�R�5��"50��5���ߧhy��vP>^�t�]՝��n%)1̱��t�ޔ^7���f��Cڃ^>�9����%��ٝPy{y�>Zoea�w\���ĵ>M~-���[N�'�ItN��$�͎�� ���N���û���?;d�NE(��o���%����X�kc4B�[����f%mZ�X�<����?MbZ'l�'R��Ɖ��lNj\��T%R"���؄A�[�-eBVB,���� 
��`�����J�$�X��E���!�V��wL����8
l�*.(h�'���N�FwE��p�L+db]FI���W H� B6T�ŉ�4�7	m���9��ł� �`A�$�J X+ B%b�)XP,JA��&L�b]6̚A(�!�D�ƑX�d�+đ�aicl$d��H%�$!1lCuP��&1i�@�A��A) �1F$Ґ�F,�$!���,/�(}���T��[C*�\��XK��
�ML�j*ؖ�T-��S���Л1@�F��nv�nsuѺ�m�6D�c`��)�*6��.����]4؋�����1n�_�܈_j��g�q��S;"JQf�c*�nڶ��E[���F�M"]rĀ��:ً`ƶn�l7��3l�θ�m���j�1
Ʈ�I���17+l�2��{n.Z����mT2CS+h�.��]6��	Af��Q�;�$�ipm�
�[��cbˠ�#6���s2�� ��̱�j�.X3\���=[�vv��]0	�n��a�3�%bLL�B:(�<#O_M�䎹�c-��D�Tbc#B�Hfa(�N.ՖX�7.��0jWU�Z��ҏ:��&5��ms�ޝ!�	��
�`�TS�� �#�� D��C�>��)��pJˌи\��ݭ�Ţ�]�֌c�N�I�74��4�$@U���f#+h�T_��z�����.�L5�te�3E������P���5���!v�e�3���N����>�/w:��������.���r�$DT/Շv����q@�{����>S�VW]�l�<�oV/oc�}�3��������&QKdɍ�J���8��ެ<�����({˹���IR����m����~�����6e�0�i��V:ʼ���˳Yi�Km���ϾC�N�����o�ܐ���i��L_�cX0!���EP��vs[�C�����L��vp�� �$��^`�*�bţL:�$ɲű��r%�qfʲNdb_�9K+�z��wl�(��Xywc�}�3������wJgsxv<�j����ެ<�����({b:�t�BbR:����1P=����آ�9��iL�
*^4Q����j:4EP=�2���Y'&�-�B
Ib��A�U i]NZ�1����Ӎ�D���P7��/Շ�{ʆ�������xHL�}�h�D��*�9��d��2_� ����!��,n4�Ǌ���3����;�o�7�E @j��c��`A$H7�@�l!	
��A
�o'�k�ܓ�O���8��FGI@�w�>��T����Pyn�����s�&;S�^�3:���v��9%�;Y|�RS8�Wa�(�Z�*0�+�����wc�;�8�}�՚X���ټ���Q�G9�疖��pJ����ZoVy��a��r��g��$�;U�©--���z��ua�M��B�郒K�bv%
��u`x��{7�P5i�Y���)NapX�i�n�l��֌�N��- ��y�=��Ս�A�a6����4���.u�f�Ҕk)jb�ҁ����-T�lN�BC͝c�ɂ�@�d�)�Ene3�նj�(L;[si��3�*��%����q*t���,�&4#����݈���4�v���鿹}�aYh��S�������~Ѭ&�Mf��\��Q��V��Xex�b�bo�i�v��k���5P�o9���Y6Ad��2]p��fEe&�M��|3B&f�u�k�M��@��ެ=�7�����Q� ם�I�(��y`{w�P>��T����ݽr���#S�����.�b�]�p��d�جY���JJ��y�VvoH�F;SV�H�({wV�Ӫ����ꏎZ�>�$Wa@lJ�,v��q�F֣v�+��4#��g����nL"��������Wua��\��5�>�*�6�Je�qk.��%<��Y6e�ؠ�]��+1K�j���f��V��J5k�5(B��b�A�a��FX�ݻ^;d��zRZ��c].t �V�v�]�L��ݡ�虺ĴOpP��ppu���G��?�Lo$b���`���{������;�wяZ'�[�7eP�
����:�Xol\�[��k��÷fuG���q'�T��u�H�(��Z&f�I��*��88��y�
��Wq���w[��=C��ߞ���s��y��+m�[m\Pd֡]��X٫�6R��
�T�c7��҉�֢�N)��{��]0�U��0o��&�U�t��0�qY�����t��y��yoV��>8Y��[d�˙�nI��h�[���ʈ-@t��G�fuA�{ʀ}�Y�v��c��.�]�]�Y'�VIݡ���s�/l��P{q���x�gBbR:8�ڨ���޹@�v�v�Ε��fuG{ X���El�)�F� ��z�����@2�u�tn�\)��][i&a0[E6�z{�zI՛*�9�7�4��ߒr�c��K&,xډA�iE.í��C�y�_~z�-��}�r����C>��	%R�u��72V���}ʀ}��@�ެ��ht��FI\umL-k��y'�{���5H�Ad�C9�y��
�
ج�{�����a(��YR\�&H�.������{�gTy��f��$vt��[��P7��<󻻾^l��Uc���$��pQ��5b��_߽��!��Y'r1-�A(�
�A� ��<�V]U �	ke`��������t���]P}�:*�[�����%�JH��>������ҁ��Y@�{�T}˸���N�cn���P}�y�Xn��{�8����AS1i�([`�m ���Vt���㺱�V�o$��xԘGmUU��t�� �5��D�bC�[fYw-���[�ʘ�$q.v���]�.,t.������+i����-��CQ�ft�[L�o��Wl�s+P��q��4"�\j덉M�Q�݁׳�e47R�3��C&ԥy''����G��j��R!9Kec��T��uAG��Ue�\V����`1T�U'T�%>4
a���a�L��h��BK��Щě�~C�"��M+��$Eq�6]R���o��lΨ;Ϲ��fuG��#[Gf+c?[�c�h{zP7��:���]P}�8��goF�O���(��*��a�Xn��{�8�}�3�<ykc�Eu��1)@�l����XyoV��Gx�ǝ�$�lu�#����:n��s-����J��e��*[M-��5����O�' R]{�e���Q�i+W\� %��W���z�Ci��f���ݷ	�.�m�֕��m��\�ql�ՊeEa���U�d(q�w[��bl�r�3m�'O�I�wI%5���fg:٪�Gl�ښC+?@���?��\���l��uf��x��9ZbuD�����ں��v	h�Y%_� %���-�A�����L�Ҵr����޹@��gTyj�õ6��O%��"�(ZwVܻ�ݝ���]Q���t	�������_�}zJ��fr�ˢ7+i����+R�ԌSvZjW��D�ˢs$�d��I�m����cǈ�E��1�з���%\�����}�M(Y���|Dڡ�v�v�t��OVE-s��� �=�bZ'V�VI=�jZ=9b���('[P�>�u�ݳ:�;�WX�N(}� Y�,J+mL[uWg���%�O]$~�=ʆZ'��:�Ɔ�Ʊ�j���<v ��o�Aݽ�r���B�%*k�]�c�&w��,����߽����r��l�{V� I+�R�Ŀ1�b	X�M�֮Ö�ͼ����-;���Ն����>�E1���S�2"���Ψ5{WTݛҁ��z����]�#$�E%Ȳd��ٮ$�¶]@ #� �'�!x��iR/�O &��#	F4�$�X�B$�b�,���!��I0�`�ZH1"��r,1��1�t�T�$0&p��e�-CC2*fSI	bZB�aX��#�.h���g�K�&���֥07��b@�]ԥFVҗ�)�����'��@�W%�7�3Wo"<��Wa�,d�d�chR�FHV�$%#(��j�a�B'��F�+$/B0`h�36A�h!K3D�o, d�LҤI�M�dH�ԩM��Ա�B�AdFfC��S�2��+iJ�+BRVА�e��F�,��� BB�����/�ʹ���+���s��:9Y��[�qNTX͛]Z�kZֶ5�j�e\���;9ĳZ�9�]�6���s��q`�u�,�m-+�Q.�]7 ��V��l���4��,�5%��i���`ֲ�4L�΍-�PJЌ��l��)	a
0%#1��k��2�eiu��{8�+r8Sc�CiHȳl�հif�"�=���F�\�]� 6����v[��c�8�ˋ[�V�D�W#���\��a�1����ZKn�	��U�Cq%��^!uDE�P)[�vbA�R�d�6��mql��Y�CB4[h U]-f��Y� �5a�pCp�����4H����1s��@.4֛X�Kf����Y��Ye`61�j�h8�ҥ��ˍ[�̺�$�Rf٢���h-�ۀ��s��[M[�[X�o�����\�ݣ�B�9�D��\�ѮģMn��֮�3"�slv�Zk�q�fIYu�����ͬ$� $��7���#�-�L���M)Kh��&J�a�k �Kn�	�k4l�4�.\���[�v�R�M��K�&BV��!K�n��<c-�tr���[��W��F9�[�Ke�,%��
e�-	�c���0n�mԱ��q�V��M��Y��i�9l��s[\�e+�d]����̵�v�-�Y�B4���SB\Mu�]ml�#�E]��Xܰ&�أ�".�G�}_*�����g�qS�j��&�j D>.��ww$���ٹ<<�Gq#�\�+�(Z�3����8�}�3�^��`.��:��4X���dTE�M�#J"K3�K����ձ�k5��oo�g��f�5���"�8-/e)3��׌�-��4�$Ct[��-7�ݙ�P}�P��3�I���.:%Pj�.��;�����t�wt�C��2�#��(��a��ua�����f���N	9��Qɉ�ʃ�t��9����������0)����A���E��.ys0�Y����l�F�2�X����i+Zh�V�X���u"�*6�y�+��*���eƑ5��.�uf�&�m�%{]f�k)e�mm�����R0�8�f�՛5n�6X0��0��|�w�iCKce3���3!5йQlc��N�;윀�URw���ܞyOs>%�i��[���i�{���o�������]-�	r��m���Jm�2��n�	'[.�Ňeт��L�O��:|����E5�b�
�l6U�I;��;��������:��Bz��#}�o�v�Uh&�7d����'�IVI�G�vk��H�m�",Y0TjE`yxެ7_r���@�ٝ��S�18�����<���� �˺�>�����·��Ȉ�U�+o$�olΨ�G�Ҍ�6�*�vE��.�\��
�
��$vI�Nˢfk��~�۴��;�m;�t��z��J���f�V��� ��H����P1�c�1c���m%ٔGV�1�+s�z�m�@���[k������J��m�d�Â�he���A��
��GH�J��ٝ�۳:���yP�oVw��qLn��8�J�>�t�}�8�olΨ���õ6��U�<i�F�����oJ�fvTv�ꏰ�nrp�宋&!��P�oV.�]P{�P>�N(o$qͩ�Ycu�7p*���@�Rȝ9�'c%uvZS0�:��	�luRH2���Q3c�'7c�p��",��{wS���n��79�('¨'HZ'�X�����d�ضxs��:��ǭ�x7f���f���9���oh)�D�, ���F @� �"��%@���ٝP�ޔ/՟w�79��q��ƕ��]�՛*�95�-{�K'���sj*i�}�br�ԛ��P>�ٝP|���{����w��$���El�2*����VG��mj˶��Pm��kX�Հ7�����w�<���n��jH����n�*V����+1�R4�9��>��T�oJݛ3�ՑKG����a�N�X,6Œvk�'�-�D�͕d��Ĵz1q#!m�ښ�cy`yn�:��:��3�I#�F$#BB,#BH0��!!$!$��33�_y��`owJ`.�M��v�V�n�'��]ݒŒvF%���q,S�FH�
��Wi�I�iU�fn�u��-	��E�amu�^`ټ���e�4�!;��oޡ����@�zgT}�vv)0qZ�D�O��jL��XbPRk[W��w��͙����a���P�oHD9�ꕶءm�͢OD[/���8ыg��oL�����<x��S	�e�G��$�c�=�.�=��{�-�9��~�Ԡ�#h�>�u��L��'>�߷��Q�dQ�#Y���bHqӟ|�.7�6Ն�cl�d�+]��Uv�0�
���uGX[.m��p���lnh(�����Km�����=-���KMh�Wm����l������J҉P�mq�e�	E�Ұ�-�6�LӖ:�J����6��X6�K�1��E�%њ���Qg���srs�������3,���>���1X�D��n�6	��WnTttn1�.�8�"ǿ{{��޹@�^oV{7�Q����ڒ��-�i��L"s�jP>�ٝPyoV{g�P���G2"�A֔����Xo��{_T^��C|r扎J�`�O����`v����͜PyoV{xgdB�4벥AI%G����z�l�d
z�Xd�'se�'���<;&UdhVE
��ڻ*	%u�����A�rV�fޤ�E"i1'0QG$Ϸ{��}�7��]՝��485	Z��3e&LN(�:�KfQ��5�5�w���\\�˦�X�E��,o�F IG-�m�m^�۩�HB�+D�tJ
.�r٢eޝ$����@�C6��`��a,j)�2HF�(^7����wN(n-��Ímw䫬*x�D��������ڻ*�����Ü&Ik����Pr�=ٳ������=:��#W7����m�d�s��/@����L��;�,Y'2��g�1o$��2�jtS2����P/�=s�<�l�\ŕ�`������ ژ���o��ywV����M>	����p�b����踒�GJh7�py��~�{���a�㺳��gtȓJ;]�{5�f��<�~��ATT6�[<�|�*������q��x��j��;$u��6q@���}�ՇwL��{��,�^���K�n��NrI�kO�tO�zŒs+b�N,������Jݗ��:����3?d��h;�l�%)�V�
�7=K��.��0�rEﲉ�ĴNel����x�K���Qt�;k��6��2bQb�S,��ۛҁ�㺰�l⇼�	w<vʲ؈بڷ�����P>�P�wV{�14�k�QG�A���@�Y���@�E��*?
��.�33���@;szP�jOc��jee�%�����{ʀ}�{+������	�qZݳ�n�]Մ����R�l�i��k��
�����B�A�]
A:�n���$�@��7�;��c�����&��.�+�eڥ�w�?>��(�wV�P=缨x�1(W"��NE����r����}�z��f����ics�V�'dHt��z��޹@�{�t����n%�v�Z�fY�	�}缨�[�X}��f�=4]y��`c$I�	V	A��!]��,�"HHhp����Hf���p��_�{���M��(0(�kΘm�s]��f�9ND!evL�f�!����WZ[&H���Bm�I���@3Mj-�#j��ɚm�\P�x��Zѫ�Uі,Nբn�2���\7\Vk�2!����HX��ɂJ��d�uUv�m�JP=ٳ:���Ć�*6Dԙ?5pK�U��i�6���=��{�>םՆ���y#���$[]6�����RFT�9�#��t��������z�>��7�f���
��� P>�����31��{��;���z��ps��Z'�ӑ�]�T�P;���P>^�]P|����P�7�Ǉc�)l�GrH�p%�x;$��Or��G�� %������?���+Y�n��A��oVI?�9���K���,)*����N)-�{����������vzC�=f�k_�_�( *��_�� *�AU�qW��_�� *����,V
�V"� �E*@��H*��@B*�T`�D@��AF
�`�DX*D��A
�A`�DV�*T�� H��U �@
�`*@��*D��AB
�U��A*
�Q��@
�F� �D�`�A"�X*A��@P����D��D*R���"*
����@*"�
� �E�H* *Eb*@B
�T��EDX
�A��DE*PX
� �� *�
�TH
�
�A*b* `*T`*E"* * �@D��@D��D��D��AD��DD��EA��AE��D��A *U��DD��@H
�PE��@X��D@��A *P
�H��H
�
�T
�Ub*@ ��E *"*T * *`�� H��F�Q��EH
�@T�"�@
�QR�P�"�  * *Q`��T"* *D �E@A����aW��^� *�AU� ��������
��� *�� ��������
��
���(+$�k98�C@ym�0
 ��d��.��@	��*��È     (��m�  �(d   �   �      �             �  	�       �   <���ff���e�t�c�up��:7��m^����r��gJ�N�]9� �(���4�a����=zz���޼U�i�vt��ۣ��aΠk�=׽a����y�{���=8(  ��%���%ۮ�a�{����o��m֥��l;��{������;�t���{V]y�Oz+��v����v�]��(P �]޹��*��뻅]w��ޕwu��q�үwk޶ہ�{��M�������=�ׯ<t�]�uV�w�xPR���y�Zj�/6٢���l҃<�ۣJQf�΂�Jh�n�픠i��٠wwkg@���)C-٠R�ܚh  AIPH��[kf���-��즂�.�4�4+[`+��Sr��ݻf��݄Ŕ�C-٢���l�::q���Ғր �AR����@d�Х:��T��N�pܠٮ����x=��]t��+�@�j�kO!��n < ER@yݨ�үC/oT�5[��z0���{�B��A�ni���sO^����{���O �)"�ͪx��5�Gx�T5v���uw	ۧTʍ��]�&��
���Jʏ  �ʀR�Q��נ��G��{�:����jh�����k�5���맧����Pq��ҧ�{@L$2���  *��
�J�� OѪH�RR10"{JQ��`�	�?�%6�RR�  &�ԕM  '���5F�}�?���4��c����ᬘ�Y�'�	!$��ޯ�����M�$ I!�`BHI'��BHI'�@���D	!I�z0�����?��������c��@�P�	�w9Ї{]�e?�Y��&�|0�yg�' 	p����f��R��dl�Xe�Dɣ[�h��hf�����IX���CBh�hVIC$�@�5}����^��_v�j����r醧�0O��Y���A
!�Pbn��kW~�l.]�硫��+i��&o3��Y����	A�ـ��EB­)!���f�ߥ��z�9��5g��3#e���4��-�l�|x�p�/�2R�؊S%��u���ħ8%�Q�0�����ħ�s�s{�).P����m�%�����]����n��"áw�,��hIv�����;qg��gr�\�ș��I�b�m�U�Hsï�� #H`���8"�w�>y���|��a�s�%'�Q��F:�G�˂F���%��<�_'�rf�<�a�8��d˔2d0Jd2H�L(Ж2�`��V�o<���xz������!��L8h��%0�o�e�ȌB�hg�d��ؔ��LՂ���: ��J���t����i��rc��GGc����Ӡ���ﳢ�mp���du��_<�MZj>g�������DK�Qf��Ŝ9���R%�Bᩰ��t�9��W�c�a��΁e7,BX�O��I^��_��׺ٹ������!����VR��z�LV�.\�����QS �Qi	xx�P �`���@o6sySVs�p��٭�͉�R�I�MA�r���(�(��sq�i����pv�`g��4�As��LK��Nf���R�hm)�$����[�g�������5
�������|ࢻ|�B�|T�\�����[��yI"nr`B`_8ϼ��fG~��-	��s�;���]�@�5�6��.�7���灃�D+ �$@�I�}���۸�E��y��hA� ��K��θ�;��|�	��{<
_�H�BtXR��=��$�zVow�����`�%̗�>�B'N���������`�#p���O&戂��cs_K��f�;�r>�c������f��k04noM�G4%�
 �(�A�1�X���rMc�Ħ�b0F1�i�GH&��j$�fF\2�	�S$lg���3F��u`%P4�Q.+��Np@�����ןh>��a���9���bza��"}���m<�z#��������&��QYL����Q��5cd��#Xm���(��l�9}�5�O'��x�k��d9��a���fH��1�xS�t���v���9�� �}��#��u��"�L�t>��{�����l0S��{�WΧ<}ۤ���_��9b[�o\�4z�^�}����O�n_;�u8w�q��܄:m�q߉;'��;|&g�dy7%NXp"P�:������:)��(B$�bhE-/��b��%c��h��ѥE�M:ь[1 ��yɣs�y��,)��b���Ɯօ�%6
`7�4Ĉ���LT�Q���G��Dy���2�rp����#$�$�*�)��.��sYL�K�%y�"]i�m05�|���23Pn9a��#$���8���Kb�M����0Ȗ`pT�H��3MKsZ��KA�a|�]p62�"D�d�*R%������B��K�K�	>$�K6�CQ)"$6�`�Y\�mIY�Ng7쾚62�62����A2\)���,FIc!DQ��=�3a���ǂSD��>T�r{��Po7��8H�����fo�\Fi�;̚����@��d�$NIsRSF��Z�j�@�4������[y�Y��Õ�3�K�Η�9I��w2���1���+�A}�8>a��/�D�"� �D�(��sApu����#q�c�����[ѸQ#xl�Ac���,������Q�0(N�xmq2ѳ_{����s�xP�lTI�rC ĉ��dH�H�搦 Q�VEA��SD��2�6�4d�mF�5����9��XjD��nON@���y"V_g	��A���P` Y��@B��S��jq��8�
��$RH������>Š����0��XpML�xBY�42��lL(���jr��4�q� � ),�D�p���Z��#b�M�%�R�f��y��;)�4��.��,��4���a�`3p�d���aR1���F��l�#�Ȗ7<���4�ӓ��kl�[;�l�03���V�OYy��5#�"d<�Cg�C�e��$�6s��=J	�4�"�  ,���0�{w�\��>�i9)�8y�2��)�Q�Г����MI4 �4zR�a��� �D�F�(FQ�89>��7���8�5<��sF�F��G��tyR��=�$pnFQ,j��R���n��y�	gp���,^�,ɲ������dޥ3����H�&��hri���4&�hK���0���+(h���6xj2� �Бf�$��6`�V����|�o<�E'9¯��ʮ���\W��P�Z�;���fg��,�g���@~=�]38a���<�H͑����E|�>ׇ�o����I(��P�K��,�2,Pade�LY�%
FP��`�`	L�L�L4	rh��!>�P�C[�K�s��)����D�����rhEM��p���H�EB�	r�5�j�Y���Mb%נc8|��Ɋ�H�#| �D��J����<�m7w���;����S�3[�n���ᱶavj4�5�Z�3Xh5���5<a�KFf��dIn�IY��T�J�
ʋ��VWC2Q�C����������ed2����k54�=��ens��NG9� ��,�`���X%����4�F�<�g<,<�5�6<��#tp�)�P�h.lЛ�Q��f5�[��EE�+uLb[�al��h�FsEձ<��ӗ,��ؗ7�L�8�/.�kO<���]�)f��6 Yv[������1��p߆`.3�5��S�ؓϹ�7���8
��8�QC�DGປ3SJ��`f[+]lnOwq1�D֓VM��r	�}!�<y1�r��{��Y�5����
��	��	��;���s02eۓ�y!_���&�=9��A��Ja����{ς�cL�ɫ�Z�9�0���2	d#P�()arL.��H�$eQ�Q#,�`X	H�f��C j&�&����ئd��n@J�h,b�[bDP2���U����#7�L�^�)�4� �If\���+�K߇��\7
f�������Y�����:<��0��=�y���B���LL�0MF�5�ѽ7� �D���8rT�e*��Zm��.����
j@f�
��c�y\��"��S��LU�JP9,c���'�=|��^��0�yvS"Q%-�b�˘6S*�`TÜ�r�,F�1(`��˂���0�U/��2��#M� ����}*opמ�k�����{p�M�Ñ��(z�k/�T!m� ;�a�rBrvN�z�H��n�����^e�й��F�]%�y�[N[����[8�<��y�7��g'�oDK�e���Mh�<�X���y�*�̉r	p�d�
y�嫢�';Ѕ�ۢ�:D"

�+�B҆��A-�D�ՙpM]�j@d�G�M��R8`���0Ѳ%#
j3F����`�h)2!A`�W�ٞ��+,�E`�`�,P�
]�m2u�j��	p�ߛ=���� �hM��D¥�6&���Ħ%���/�%�A��TUR�#�`�K��-o����>��pMԺѸkֈ��&\d��DDbȀ�Od�A� ��K��
j�^|y�ݔѼ�rn�4�x�7��ݎ�{�1���h�%�`zّFT��Od$�b�7B�{�x]�3Z��0�J�|��M�n2���%�i���@&�<��sA�l(d����'�VY�@�� �zz9��I����\����`)5�t�g��Ią��(0c��`��dK�R1��Ȃ�&F �B�l`0)Ɏ`1�����B����`s1��46�4n8�aVa�%#L���e��o�Б�OW��z%�l�ޤ�3B�4Df�.Yd0a�ڞ��Fȓ��%&<Lג9�d؋������F�ћ�t�4lt��ʕ#���*�*�� �Ys�nA�44�7[NA�B3�!U�I�7O|o���%��L4���.H18���ߺ9��;g�(��4��t��EAV'=�DO��vD}��}/����6�´�~n��	jM�.l;}�"*-�� �U� ���4�]��0��F�@�����PH��r�rm� c�mIRIs�{e��Hy�$
.�6�b܁AܐD�ht:�w��� �H�CRIi|�8��r���Z'k2 9&L{���2I�����{�w%<��4��Wʐd��=��μ�tX�C���GBL��t:�C���KRH:	-�wj������I%�x ���t:�C���t:�C���t:�C���t:��$�2�#|�a��t:�md�����t:�C���t:�C���t:�C���t:�C���t:�C�Ƞ3t� �%��$E�@�t:N��C���t:�C���t:���9�2$�x�(L}�}>���C���t:�C���t:�C���t:�d��$�����t:�C����	L���(��o>n�3��4't�H~�ۺb�[�`��Rw&��n�j��	H�IS��{coռ;ܧw3ߟg)�aW]�E�'�)��[Ͼ�R�'�����N�<�;;�s�\�õ�9wh��(�n���Q3[�!5 �v	�$����,��zO"�w#=ѽ�ͺ&��G�Io�`4,���Y8���'���Ʌ�	^�v�My���m��m��i�۝�^�
��Fd�vvC���g]]m��N}"k��޸�Jr[g/���m����v�Eo��դ·x�v��F��lWR�GOfl�c�"�F���۫ =y���1�ITm0H����� ����tX��^$����h�:EA`a���n����/��i\a��N<ã���L���BH0I%��E�Y�i�KB-Q�;2�$E��y�S]��O�d�-���S �Y���=�'cm1=�p���ӵ|��͸L�繣�.�)���W�=$�2@��C��R�x=˽��ى&����n�ۥt��Qht<�ޣw]���������d��s:{')�7�q�6�*zڍU�˥�B� wr�րܾ��-��X<��w6�`>�9�P*w�qIGS�W��4���2�Z����w0�zz��Y�6��y�)�k���H��q�u�>K�{˫cW�
���H�P|��Ǹ�Rz��	R�).f[���3(w�	'L�L6�cĥ$=�dD+yЂ��ř9$���|L�Ve]g$��\o�N�aN��U%��n�v���g.��2�T���6�-'��P;�$���'��� ��w�N�"�K����n��6w�o	+��| �hu�tt�Ý�l��^��C�!��N�Xܓ��͚$  ���n��J�ِ����l�H4÷:�@"���q���2�l�6I����1-P]T>n�;9���Z�}�|{;]�ˡA��C0,o�j�@�m��3�fv��:8�Yv�-s��f-�|���=E����w׻� �a��>��B҇&�@��� ~�M'��3�p�;���~KI489%͋KC�C����&xH�C���t:�C���t:�C���t;%�H��$�C���t:�C���t:�C���t:�C���t:�C���t:�C�[D�[D���t:���t:�C���t:�C���t:�C���t:�C���t:��$�@݂@�t:�C���t:�C���t:�C���t:Ht:�C���t:�C���t:  �C���t:4�e��ݭ/�� wIu���vs�J��;�#C[<kt55@`�<$�hu�`��v�}��EpG�6���q�b�t��>�҇�&ss��Cٓ�K�N˂�9.�`
�3^o��:��zڷ6(�Ԯ������h4���Q�t��-�k��^R�z�[�ٰ�j�r1_�����/|��O�{���6dY�v�;�\�����}�	c�� �fR��~>��9Bpy����>巴�[�ԕ㺺��.j��𢨻� �S�HRI~�u?�eݤ	�ϏK��q\�Y��Ev]+f
���Xj�k���B� 4L���v}�2-�V���uǕ|������ k�]��p���-�L�mޠ ;��p�@X�J&l�X^g^m�-���,ݞI*����<�n�.�t��G5l[M�1B���S$�wz���j��|���ܛ���d����2L��ۭ��/��H��]�\5"ض�r��
�u.@�_ p���V�<p.��O`�gYi�m�˙�T����gwL��tXu%���w ���sv����oO`�z��� �s�|{��c�W�J�ը��3{v��+(�;�-�b�, ��1�!�|�kg�ګ/u���kHA*ħ��{nh�B�^8u�z�]WP�u	�Շ��0�d����7����Rvtdy��@�u��\�<���i�/$^/Y�� ��Ã���E��I!}��a�3��u=%:ٞ	�vn<�݅mFr�#�k�US<i�1Ѿ���=�'?n�Mg{�y�{�y����}�ԭ��<$9�x%	�$����G�N�����s�kk���qz����%�W�������͘�ct�$1wK�z�I��ws�0t�yK�67K�Pf��ē�a��(2(��a����r2�Tnr����}�<�[XPm��'(j(�~�̡��� WC���b2�/J�lw��gDw�u��D�ԒIf6�(0��7u��R$�@�/u�X�y�Tb�M袦4�ѧ��ż1�a����Ԇ 9�@z��!$6�+Uu���V˅�?6�SW�m�'+ʄ/%X|���TĽОI=ۇ��:�h�J�L��/%���fs�y1=q�_�0c���e������L���aq.6���w^�Z.9���wͼA�����^��� �;��n�	o�q�9y-���Q���n�w��hm����,��|I2,B���f���*d�̇8y�r���y��L��[L�{k���w�0Mcק$:EiL�A>���8���{�D)  s�;7D�;8s�@��И�7������a����Tl%�6:�wb��wZCv��l��g�;}9����z��wr���P ���-TnQ=����3���q���fmm�<�VC���t�W�[Q�# �o��QT	�e;�I �ίM�wwL>�C�F�n�����O�&�lÜ�و�/x�N=��5�C�ы�);�di�s\YA���6��Z�A��  �v,z����������%��V����]���fM_�8 �v!]~U�B�ճ2�a����p�G�!�*dy����4�9{3.�zN��?j�oKo{F���V�*Ü�櫻� �$��y���i=ܝȭ@AAq'=�#$Nw77�H����ƭ��"�%>%���$KgX8�J����;����{w_���M<Nс��r.���C�P�Iv/t�ݒ�M��bp	��&	|`}��Pg��{�����9��m��zC������f����K�¾ٱ��r{�79Y��߇svQ���/����a�]��T�fg;��Hog�$���,M��1�CSP�=�.hyh�πĈZ�ks۴�)E�\ր5x�H�n�Mက��wtk��펉{��gI�-'
Im�ؒw`u��Ժ�
����-E�}$×i��`y�K;�w5��2��In�ǉ7I\4{��q5ܫ�u�1�����'5uZ���c�߷Bͺͤ�ͭ/N5g����t�7ٗw��&�����e)����z���hŪ77'Ä��ݧۤs�P:�_���ۆobO�o�Jw�7��	pM� ����lHb��"E��oza��?>�.�4oUn0Vx�+����~K:t�4��x6=�����|�蝓�7�%��'�oSt�ݽ0�X�·�;8��S���Œ}��.�u��pp�۾uKI�!iu�5fPm��S�{�?F��S��x�*�k�'Ob
�E��1����������X����3��Ǡ���
G4H�$�p�AA�{jx ��ɀT7ѭ�z�]Y��9I#˼��=u'|;���0 ��b ��V��[��j'�t�� �b���L�"���p����؈�CfK �n�t�	���U�{ջ���0^4��፸9����[����˸�npT����r�U��Ar=��ʻ�E�Vb��ٜU��g>�İ�7^w8Ne��ZwJ�2�Ӭfv�r�L��=T�$�.kJX�~�r+��K<j��9�3���>}�dg����B� �����[��s=��m���3x�F"��db8T��WH�}S�ɠE=�m;&��o������ pΓ3t���H��$�m�f�qg]i戠@N����]�]�)s0�&C�<��|�m�W�v��>l��͢�B���9�0���q��U�#v჈�7̿Zx����~���Q�#����_j�|E�s{ۀ��$	@��=ų�&��P{��#CKw�}LP�1��ִ��x�K�QS}��A����t�&l���S՟�>vtNVFc��ć��^�Ę�6���>~ؒ�o���7��
9�m�6�=�p h���3�og�z߹nݻ���I�E�蛂}�c�:21X�If�t�#�k@8�K����۾�9�,�K�v�h 
6y�<����^ˊ���{���&/#��wz��!��Cb�M��a,+�ͺ�u���rƴg?p���k.u. �D�B�9�k4"d�?m�IB{[J�9;�;��/Cy!K��J���PQ9^^���O5�Ԓ�i��.IѢqB��׻;=�������)��y&��wE�l�����v$��������x�1y�j1$���އ/�w�������ssC�n0F�a���$�(�:���>xsV�ʉC��N�/rӜf�y�U���Ԓ�2���twd��q�#l��h��.��C����oOw(:����\��jINT{��G���[a�I���n�R7�`p �j˺m���m�<O�D��}�8!I�����I}%��.��Iʭ��8���0T9w�r�$^�K�䚑�c��D�` ��6��p>���~O���M]��u!���s7�߸m >�$�ʕ��~�-���q?Ͼ3���E��q��D��n�W��tډ�Q�� ݶ�"�Y�Q�s�i2����{ŅZ���0ؿ3�4N���y���8�n�~:PZ+��&��x��r�`�;ӣ/'/�<�.�`5(>Z��9�<M�����_.�\�(������]n��n�W��M�u��[�O!�̤�|�J��\I>�M��Gݙ���<ǹk�<�r�ʎ�ε�y��\�D�	(۾'��$<�;�J"�z�_w��F�����:��C���/��\>�'���l�W���rwo�{<����A 憲��|L����2jy0<�"`Xk"@�p�K��	RI^Ĩ^B�R�a��Q>��$����o1���~ل�(�Y�d��  N�週 t�HX�e�$���7�Ⱥ�$�Wn�JQ��7����$Ǫ�wvl�����T��)�;@�K~��oj���r�`=��曈�9 9j�"Ă\2$+5I�4ת���}��p=_)����X������գ���t�M���ɘ8�7}`��e�ɻ�d�'vy<�6<IW�-afM;t��d}_��oN�[��30��!���C�F��K��s� [�\�&��:�ļ�w�gRG
�V�y� �é,>4[�2D��/)��ۇj����.��N��Ƿ�-��"wmZs��n��?�KZ� t^1J8٘�K�΅E��?9 ��$<��޽�|��x�؂�i�LͺNq�wb�;s9粿ǰB�.���9�8e
჆Խ��+C 6��X2�GI�;fwg$&��� _l�������`|i'wB���SZJǵ���]����nz�f����h~�&��섌��������W��<|��1k�[H�H���C�I�F��썗�n�Ԡ82i,�H�n쫻��x*Λ�Q�t���� �ZHww:���t:~i%C�T���<T炋jH�6��% �� D:�{��U�:<ޗr$�����rB���$�  :����w%�γD����[H7uZ��Ѻ�j��g�����w����Ā��Hd4 G����O��}��@��t�0�A�؃��I�C��{�k��a���q�����U��C������@:_�X�@(:�A)'{��4H���l��
���wi�j�@�t:�  }4�	$,zl#v���t^V��a��KRH:��N�x0�%B�܍�N~K�uS@������`�8�C���t:`�wI"n���^��3�.�A�O3{ݹ�� )Ā	�4�^��87��RC��]��Vb��ZH� (N@"D�vQh��t*(l$�c�0ސxA�{a����h��>�BM�ߝ��}��9�JRi�ے��'�]�n�j����I%$��X�M������u����]1�{�6g&V��D��V����;���'���˶GS��5Vy�z���R�2f�=���Dv=>g`���L��a��4��sg!�<� �%�Iw�@ ���ؒ� �n��N� �� �C�۪�cu���2��o���n>��nHi,��-'|���	��wF�u��g:�ܞ�r���h
�UP��	 ���N�r$��I�$;!	���H2I�	$ ����=�	��@��� 2{ j�X
F$R�H#�A���( A��$A�$`$������Q�	F$B2AX�DR�H�A@c� �bEA� 0���b��2��H@< ����@�p���H}H��#$�9 � ��D�� ȱa��"�K ,H����� ��|B�$�j�$0�	�@!�0!$�Hr$�!9$	�I>�&���� �I��!�H| �$�I$�����rHI�!�8H�I�����`A�=P�xAH�H�		�9&z"H�O��@��I 0$���@H�A�����$!$(PVF0� xI%$'�&�@6@,�Oa	DRF#��6Ij%��$`�HD� !�4����B����$�L�	$�C�BI��H` �'Đ�nI� ��C�$�Ԓ�BI;G���I� H$��}���\���Wl9 ��L��%
����l�+����k�^F���l�:�3��3��[Qc�*9����yЩA�ۊ�'��T��[UUmUUUJ��+k`�Uy{OX.S�����&6n�T[F W!Ř��3�b��<�Be�<iim��l�-���1g@펨M�i�0=%)�pm1ێZ✰ �{1�R�F�8�n��#h��;W:3f�g��=�v�ӈ�૮G���<(�t��Wқ��w`&%WD9u���Sb*0ut[ =�q���K��ݗ� ��⨸���ϓyv�(s�V��n��^˷�8yܼ��v` �2�㎘��p,F�6�V�
k�1�����d���\���<*iݭ��kW=$��$, z}� � B�Od�O!�n{�(nI}����k���*Mj��8��0ܷ0�]�%ƈ�<i|��Үn����nغ������d��۫sX�ˣK��I$�!��.�X��m���jɈ���a�t��{��W�/��)��T��=&I���@>��X}m��>�)����$�zn4F��=ze�����κ��t��ޣX�X,�㚘�&3@�z��e4/u���4=�ǂ�9�٩!I3@��˨3v&c[Jk��h�f��������J�j'5$�K�ut�e����=���a��M�^��!��n�Y1%���q�@��)�{���W�}�SC��!X���LodW	<�d�B�2�	��I�z�O���:�AE�lnfȣ�#P��>W�������_���g����$�i�OR�M�Jh^:��u�����K���f�LI�����	�mw��24��4�Aq-msb�ŏ���֥�߿g�P>�n��{�н^'RMdǦ��l�Dy��4��p��uY>�o�+u�.���)�yx���ԑ����6�6�z����Pz�V���.���*j1T�u��t>^��z�i�����31��[�*��tycrDV���f�iY;UUK��v���4z����.����H(9�wE�BH����P-Z���PQ��^E�����]s����?3}�ְ�ֽ�빡ꎭG2e�F���۰���v��i��7B��v�w4/��.���A(jS�b���.��>.���s@/��̾��ȏēM�;i+����I<�̷��	j�p���Oz��h`��rCi;!�.�<��=��>�2�>��ś5c�pqM
i�5��~��6�[� N�õq�Q�I��@�l��=��cWGE�2�%���kv��2��R�W
��t��b[�+�=�5\��۵7Np㋜L����0�i4b��A��V��I�o*�+��{��?�;h��o$L۷l��B�'�Y����ٞE�:=3\�ǋ �j%BdSL�i�X���9�d�3,Y�+u�*V�0ow=�mLS���d��$�K�D9�n�^����u���]a�t��ys�5&F�ݛ��cz�����w4.�u���ς�	&F��Ů,��y[�<����w4/�8�]f%�Q��Fk{�4�L����u���\��7z�խH�����{��2�㵕,��m7#�u�a��d���92L���s�yqn��;���	��9�D���BH�z�YM�(on��k�є�n���%.�p���C��9�Lڔ4�!�����HD���B�h8���se�{���z�ӎ6���爋$��#π���@>��X{�)�}��<rIuMk[�&Ѭ�{2��*�:�5�'�m�yܘl��ɬu�Mj���5�U㮰��4^���V�=�b�x'3R�m'�Lz��v������h]��}WYl����a�>���!�w�����0N-��K���Nd��m�o��p\u�����.B�n��<�H~!ƱH	�M�X�����V�{�e�{ט��;�m�zJj7�n�e��kZ�W��f� ��B��Ҷ�RT4�da@,�,
2IB$	Y8Hd �{}�>sl:�M ����S�ɻ!�ű(M�z���Z�����L����RH�5�G�����u�����z��-�u��!�����#4޶hhZP��
VW$kc2	�B9�F1eMD2/}㮰�n��ֽ��df��o���m+Ӟ��1[nn4�����.���U�}^[�=m���P�r�)6FDHM���e4/Z�
�k�����f,Z��6O͚/Z�/��߳�3�]�e��hq�������՛�$RMצ]A�ܮ���zץ4<\�ܓh�f^�G�{~{��+�\i�Ƶ�`����q<�v���1�Ez۟|�u޶hg�_���o���{^���8a�7D�x�rbz��yn��Ϫ�=ze�T8���[h��%"d�n!��zץ4�V�
�k�/[���Yn8��&M� �z5� �[4�L���yn���V���v�vjdLq;Gj�����D���d��%�!]Ǹ����g�CY�^��ū��Ps�Y;L�m>-ֹ北`�+��BƇ
�d�Ǯぽ�r��v�=��fG`��;F8�gn���S�s�c�l�+35�Ĵy�hL��1-c�Aw<n��`9�K���>���U
� }�[�χ�ǂ���l�s�/[��(j[?D���hQ�\�q�A�ݛ̊�]@u�h�2�<{��I��7v`��a�������7���I�O�^��@�t˨=�2�
�ס�^�"��$����h�����4��h�����sʈ��؞�r%0�/�e�s�u�yڴ^�u<1�ȋ�.�jZ?UUAk��d��f�$��f[;T(R]��d�&����lrn
I�G�^|]@�kk�k��E��c1,15nά�q3����H-��x�Jhy����m��j�Z󓜣����1�/g��zs�f�]�sE�^���ܺ��v���YX��X�)tv�4�ngU�!��F���K�3����m�=�+(r=�=���7����)�z�˨*�^��빡�rki	d֢KP�`���V��
 TGsvŒw�I�����"����#֘�a@��[�>�-��)�z�˨�.v,l����[����v�.�o�NbݶI�,�d�,Y>�K���4٦#�{��sZ]+ӽh��ɼG��m3��1������:���u����.��{{��h��b�xT�LDkヌq�4wL���;������9qn���c�<$���k��\'=�t*�B��Sg1��O�皃����J���2f�0�f%�`w�[�;�S@�t˨9e��^'R�8�կ"[fh��Xr�/u��/>.����A��Mou��s���@Y���f7�Ɔ�����j73gd%�ͪ]�h�Ͼ���=^[�/�SC�D�51�I&�~�lmT�:!�+�W	��9e�>���.-��[��=J�f%�v=Nd#�4Ϫ��wPw�-���T�X3aF'-݂.�r.��d�d����#LxS �4$��,��R�h7!��{�VѸ`_,t"Pɤ�DI"l�%�a�+%���+A��5��h0P-���[5�r�1��$3f�h�5Hf�%�슂���0H�����0����,2��ׂX#$HIc�� �r2B��¢#I&�0$�+Z%��.)�@�)R��R���J�Kx�J��6R�l�P|<bE�-��m��b�����,�B���AA��eU"0��A榟F��"(�[Z)�Qe0�Dp-�`��5�Q�$�D��# FL|��ֵp[n���1�6j�ڄ�8��X:��Wi�"!����؈���"" �Α�UםĽl��0����5(7k�4Jg����;���1����<+:�����ظ�źm����ndR�����Q͡��F�T]+��tТ�n�N���t��*DF�DDDDDDD\���h�Pܫ�ֳ�\N*��P��nZ`�r`��E����;���Mϣ�e4��m�i�f�1l�4Zl-���X�]L�wI�iMY��v������-��������g�M11���7m��:�+�q�����,�K�8�鬙�h��M�!E�^��\�W0�v��a)NW']�=����eS������,(�a�҄��=��y�n�Յ�#ٻ/��@����z��V����ݴqg�)�N�U��^3qY�2�5٪\ny��tl�pgֳk���WF�:�.���&�1���u�gr��l���Ͱ��⵴x��돡/���v%��㷵yJ�@��������0��tS;�l�vW�k��G&�o!j�Gf���=m�@=�r\j�◲g��:�é���6��sz
�vy|��OyI��֝�A��DGa=��c5�GhrYC���Ví#-R�M�:�p��������I�H!'�&��! � y ���B�=�;$�$�D@	��������í����krL&<���v�h�[�/t��{��ws�����2G�Cbz�ܒX}��ܺ~B��
[��@Fq�e����9��,�}�g_�}�e��)������ rk[��dƛ�֥���R��v�δ�{���OW��O1f}UU�N�M6N�	�()�٬5��<��wP����)�w�[��u��Ặj�G���>�u�ץ4+kХY�����TzB1�{�Jh��hy[�i�'��y�k�7�,�*�d4,o%�;��%�|�kFAi�b�s�Y_n�jx�Y��]=��;�ͶWV��I���הX������a����dI�������ͣ���[�c��Nx����8�i�<V�r��R��M�ܦ�� <�M��Ϸ^>�\��sw\KbsZy���Oڶ�0��l;LL�F�(��b%n(�ɄS"��{Ӎ�y�:~Bߴb�kޝPٺ��X��<b�7$�9"�Ъ���]u���/u�����DdrlZ��LZ��s���Қy����]G���rD���M�ap�>����u����١��M܏�bzjfG�^�M �V����wJhx
�������Xٰz�L���?~�9��'���ƕr��Dq2��Z�F������g�h|���d����G�)�(���s�(F�9<:L\�b��D��+�Վz�i&z�j��Y�$�ţpٕ�3���5pH�W�Ӳ�u���&e��
���#� 8kC�ѩL���!��M��m朧5[�֌El�]����޺��/t��w��u�O�lM"�v�V��_���{��;�mצ]E=�6ԍM{#kd#�/�Py{���l�>�SC�K��qc4���8ހ_[4����u�ڴ-T�j9կqi#�'�=}����@r�V�1�����s�����f8ݸ�n�Y:����@��Py{��{=�;�a$�z�C!��f�6��t�s��&YR=�e4�)��� �+u�Zb�H����O�$9Ȓ�y�߶� .�,���q��z#��Kݙ���Slb�q�j�6�N8�$��b�q���dԒ_^�}�I��Ѯ��恜�k��|�KE )��cm���/�����ORI_v���.�J�Ɍ�+{Z�s��������3�˥�C9ݍ���%����#40M0�>�K��]��%��ѯ����ZK{珞]m�e8�j	���@%2L�q}�^��ѡs��~I%ze�4�����_�ȐG6n�.�.	#�h��9��X�#��+=��$��,+)t�cl�Nq�q�j�^��m$���qr��*�
 .��*���H����_Ng9>�x�(�6ӱa�\j�[@A�fsO8�E��v�����-�@Sǖ��k�^�����A+�H��L�m$����N��ĨU�{^�&Ha2dP���F�}�W�i$���m%��O�Ig,�MQb�M���$4-�qn��E�uKV�=�~-��W��RI{�i��$,:��W�ۤO����_|b��|�\�"�i/vg9]ɖ�����s�(��S���e�[6-D�^�q$�}Z4�~-��W��R^=l��}��5/�Ndk�HX[wu%�]��$�]��G��Z�N�"lt��뢄��g&˻-ҽ�|�\C3��<%F�-��[���!%��p��vp��\��*���T�Wk���v�8q�7CW��ܛ&�7f����x��6�����b��4O%ƷK��1!���f���}�h8�d�lz��ⴒ]}��q��n��La�Mm�G�Q�K���7�1A@��^n���v���${��F�*]�+�r��� ��yEqeЌO��nb��W��RI{�i��I,:��B��i�$��Y��-&�675%_����)�B��+�̤W��_�?fވ_9c����H�uز�X�s/�EB�kuM6Z[��}���ѡI6L0�Y�-���f�4�/��Ic��_!Z��e�x�3dm ��.Z(�$s�$���|�o��.�^.w��M-�#��m��p��%��嫍8\����y���5$�~-��V�ƚx9�֨�/�T�P@��9((r�Z����#�|[���:Me�9�K����]��u<r.�-Zh�j��Y�����hdhM3f�����	�G�4m�.snc5���?�����~����$�]+�r$�ه6�w�%�f�i/{��U�����<T�|��~����U�f�s�$�c{m���s�Q��֢���f�ٌ�BZI-هyƒ^�[� �M����I"����b�q��s�|�Q�
|�Kh�oK��X�syȒ�A[k@o����^azA�r]�S)ڈ[�.<Ŝ�IpO9)&\QhI��J�n�0�(�!�=�?��߾�$�����i%�L�����d�� }��|�6,q%M�VQ�]�ߤ�m�<��>��Ұ���\���q���a�;"K�~�"CP��(�ɻ�ݨ���m%�{�焟ђBC$����死����Ic����4���Ŀ�4jI�N�P��s��,��"I}��m��p_«�U$+�K1%�﯐�x"��,�2K����_U� j�}xw�r�i��m��8/�/��_ *I�菱�	��!.s�|H�8!�_!H��bYH��!�i�]�_cp�k[:l��AI��e��U|����Ȥ_�3���wv�~IU�`D��#Bѳ�L��l4m�����������O�I.���ߠ�+2�~�������D��L[k���˂	�>s���c��i$��%���_��K��q���~�l����Ns�T>$8��T�V�R�嶒����$Ws��^�C� ����r����sV������z<IA��.Z_E�/�U}>����K3l}�4�]̒�_P�o��9����\�.$�1�1$����$���{<�t�Uh-�vĮ-i ��f���u�K������������I/�o��$�]�r�X�6�B���~~�5�s+�s�س~�ޡp��
��Ku�e$���|�Iy�̺�K�����.ˍ'`$=rh�mnE-$��g9�
�����p�I%��ӜI%���@�z#�79�rZ�9�H�n�i$�1{9ɴ(���F�Ik�k�]^�\0(\�p�lZ��n�� 7���K��i$��s9ȗ@&�b,��IahRH�F
d
��fc�n������ۓ���^F�t޹��b�LZ��Y���6�}-ٛ(ݛWD�(�[g���K��۝6��t�<<�4����|q���	%3a입}��Fk�v=7q����]IѺ�Qx���������&��������������l����n(��w��#j7�-����Z0a�]�WiT]l�#��Ҩ�����F�s����C�@�#7w��I�ߥ�O:�-�afR�[ӽN�WGl�l��cA\��9����$5�����{�6��}�����t}�O� 	$�)	�����kߺ����u����i.j�ھy�����!I#!"�����������~v�������2��$I3=����eu���ZKqf�E4���4s��
����0�<�H{"�"����b��?UU}F�(EP~�}l�-��d�� �G�U_ A�	�麾�w�O��l%�a.$E�}�L6I� �Ip�ap��֭!k�Jq������l�I�C�	�������[�;$���-��F�R5-�k�}ES� �$�i��$���ˉ�!����[%��#s��jk�o�\�嘜2�`�k5��&�E9�<�,]N]MJh��q1FRd�ӛ����{������*�#�����6��I�J�zڶ���NQ�49}�Pq�Qp� �I�|�G�)O������2 ��^F��(9MF�|h7{��(##[L��a�	�V����FbFDMLـĈ��x�C��H"(��6r ��D24��%�'���8y��0`�V�$n��IbCcY�����R#`�����`�Q_8q���� ��1���g#�m��lXYJx��m���*jZ#�02�Ĉ�Hȉ�j� ��QQ`��[h�c"0CQ`S)10+�PH��4��Ol��:�"1�<޵�ha60F0A�\js{J�(�*FH2FD��4�Ȣc���	�T"a�|�k@��)TMY\��P3B@�yɍ�d���w��a�g�-�H0㴰U�*X����[Y��6�q.���9ȵmҭ[%�yUX��7��X���E�+H���1]k�V�����U�
���{�V�UV��.�rҫg�M��Ɏho6]mq�@�9�m/K��)��1u�����{��tQ͞GI-f�T��K�K��b^h5�mnҶ���;�Ռ��v���1gm�U���k����5&�i�y6�"-�+f热����qط
����pB���%�c�jö��͋v�V�x�]�;�7V��qۧ�++B���1haК�ڔ�!��ɘ�F��)[Tj����0�y^"S)��b��2v^1�<oV�I��-�,)�t�j+�rI��97;	!�!�H����OB����ā$����y�
�ϵ��Tx����$X�cFg�V:�������X�ѭ�*hg��`�]��B�3�S�b�v{gu!K�7Ca+퓒bf�8l��͍�p�Z?�W�$W9}���>6I�}0�'�c3� ��>[����_"���v�ZlE��'�Y����l�}��$��ύ�w���U+x���֖�d�zs��]������/_�^�?�a��R�`�S77����u�'��6�'�Y�΀)o�x,���$�	��I�Š�n�DG�	d�C	���e�X�M�2qu.|�u� 9�͝$�=;h�^��DgFdDf�wz�Ni{:�$&�[�i�b�*�j��8I�dh�u�e�x�k�=�2�=��X�0�4pF���ֿy��7��4 �0D
@�(75#''�!4(�1�De�rnD�$�#���2��Bɭ�(*(,l�r���'I!�{�u�j��~��<]�w�UIw��=d�-�e[��퓫1m�O{�,�
	f�زOq��g��k���ڷ1�� ^���D�x��'��X�v��-��'�3`�(��ֳ`c�!�>^-�tՓ�o���c�劸��FJ�FFH�e�u\�����u�w+#����m`8�4acaʠj�d��@�6Z�p��cv�8�}���ra�
�(|*���Ňﭟf��q�q[r��Y'3�b�UUW�D �?j߭��ﭓ�{,Y<�>x�D �wi��4.}�<�O��b�T�@	]��	#$��I�H! �FBD� ��A�� �5���O������XP����Wj'�
 ~ UP���6���l����d��e�'�@�����$��џ�ߙl}6��C��J��>|����/�n��g/tǳj�"U���5Gӝ����F}�o�j����Pu�sC�*��I�f�2pW�l���eX�R��o��Fe�{ܘl��ә�UU�  #�O��������	��vͦ����Ny{/@�*#է6�9��,���z(U|h�"��h����r���6�߷�I�dk�B�	bûl�{f�'�<��ˎ;rʵq���W�
��@�������?~���$���[%Z
\d&Da7-�D�]�'��xX�[n�c���� 8��N��^�W3��[^�(��[r�"��Ze����X��`5&3ڸ�l��i�x�g\�e�B��Җ-�mʃ�-�v��m�x����4fv����w{��!:O� A�'>���7��%?~tb�Cv��dȈ�Oz�e�P��O���E�c(����Q����e֮�Ѫ���� 2A������}��,��dh�s
�!RղV��@XA������q+���0�'����<^>ͪ��U$�$d y������~��hn���Ĭ �H��x�s/hP |( �P��#$!�{��ٵ~�?~�U��s����A$�Ad�k=�Z|��PvUˉ��Y'�}>6I�̶Oz̺��ֽ뎱��)�ބ�oO@?0�`(�$���y�گ{��گ<�}�z�d	�{��җ���a&%6l��!#����{��>,q���)�z;v�[\F'6E�c_ܒO�s��������'s��O��e�Ο,E\�v�U
/(?\G����"d�x�C ��5B�������F�-4*��0�\R$���bH��Jf�R��<P����L�Z�m�39��y �,I9"�M��@wM�N���fX�P�U:�?n�,�j�L�wmn�p8�}�L7�>5@ @�����d��[��s��O��6���wv�2��1�l�� �_�(�P�F�M[��N/�߭�ﰵ� ��-&�EY:*��F�7����'ڷ�d�ޘl��ThT�/>��� Zp�n5�&�^빠f� �[L�1�+/2`#5�\�ٌ�
GVk�@Y'����a޳.���J!+�3��Y��+�0���musW:H~����frj����o�fX�I�{&�=d��}���(�e|"n[WjقF��޼�c�(
�*�d�r�9�Z'�Ɇ�UUU��F�"L����c05r�ʹ�;$����h�����U�(~�T��?~�N���œ�`9#DNkrjoL�h��@�Қ��e��P	wٲ�Ӹ�E�ZW
F�n�=��{A���h�&Y�cny���:�ws	�g�� ���ĝ݃�D�t�[#��2��}P�x��݂xm��Kx�Qh��h��������߾A���W��!�d�S�3`y����I�B�d�Mi���G�����G���v��."��Ǔu�58�SPy~�x��{�m� I��;O�d    �}��,�wu�h����´�6�n����C�@!��~��ڿ~y������f�{�]Gv���؞h���7C�ڴ�Y1=ҍ2$c�v�O�1��D��3P8�@�@�}��D���������>���̻g��{7l��E�CD�R��P |%��zI>�_։���^��>�κ�{�G16���P�҉Y'��2�U ?UU���c��d����O��e�C� ��F�����"���r1�6_���z�n�}y�A�^��YԐ�HlOpZ$�Z� �?e���'����<�L6K��&H�0A�A( (���D" ,	����8�ۆ�zt�:ٕS�uI�CSH�GD]+s[�j���ma1�+��#�F�l-�]HAn��!JX��H��[v���̝�룠���6Cs�9¸����rav'�l��Y��Z�s�v����ZBƏ�*���(
� �Ŷ?~�wۥG�)jÚ�X�K`w�˨֣�#��.ŕ!f,�k�b���G�3{�]aW���n懨rw"^�������AMs	�-�`��P�hvV8{	��W։�,Y'�c٢��ݲN�߭�|?�E�aB��6I��̿�P*#�76�9�l�}�콠*�
����m�Tݘ�V�{�����}���^WP{������6b��r�K2C%õB����߭���|l��әl�C�(=�w�ۨ��	�?=դb�#4�u�0&İ����ڜ��zX���:P�c�B~��u�^����u��>Ӭ�6�{��} �c$��$A�HFA@�@��$d^��-���ܥ�aGW(y�M�\mX���<�{b�'vn���nrL9 ֊W.�3)q%�eU��4хGh���Ѣ�,&.N2e"چJ�}F�|�'�Y9����y�X��X}�)��V��Nf�ȍ�p�R�O����UU}U�� 4;��~6I?|��l�/e��j��o�ߋRH�]ۆ�ŒO����q{�5����:]F[�԰�l�Fh�9p�C��@n���d��>�l���~ޟ��'�@�#k���v����`")�D�m�CX|��6@�\Wc6�&�u�ma,L���1ɉ�����> ���a�����AX�S[z��!#yP�F�kK��Z�у��� �$B@ܰ{�'u����{��l���e�~��u��Ddƴ�!�BFk�����F	4OJH�P�$�����"a
�I@a�!�b$p��$H�Bd�22D0F(A$(�c�Id!> �ä!�� )" 2DE

����d�Zw�d�}0��UP����0�00�� � H� 7��|�H����`�"*�9�O։�fX��T*���i�I�,�g�1<�$�N6��\��?UU�Q� A�@I�I B$��B��_�+$��7�d��Z?�Kۛ,<�O&'7vbz�a��)�~�w�̬(�T�LΌ̹�iu�2�F��ॺ�?$��d�Ȁ�$HF@��  @}���O���Z'�̱d��ĂH��w�hǙ���bl����[�I�W��=�2�<��Z*�����0a BFHD�bB���k��>��5���mٴ�K��}���d��F$`���# @�Eϖ��?fύ�O;�,�$��7ZL�2i&AHf�w[��_t��d)# dd���]���"�"�L�A�-�d%֡��L�ffB���H8%�5�6X`h�j$���(KL���1 F�i�a2D�!l ��(j�� �X"��@�堹�Ȅ�@bh���D�H�F�mie��"�,$,�!�!H�V�F (ĥ�����G�<��>Hܐ�.��WnUG6up�+eUV��l  vݒ"" �����؃v�y|u�r��'��Ű�������v�C�����ti���:��6tű��QMËT��W3Vkj�F^���Q��)D=�3k��4�M�8" �����""#4DD� cNg�.m�c;u�#5C���`br�-vA�i��c�hL�fon��V�;N�W8Y�g�.{<'T�rv+���"����M�;iR콽<��ض8S��=������m�v��Pw\nB�ƨ�S�3���z�>�k��^�:ⷪ����t�l	��&--Ѵ#-�Jl�!6�r��U����e�:8��,'m��Ǐg3W�szGzM�mͮ�si3k�q]e��2����:KЯ-�:�vۑ�Ǯx��q���J+,,k)\QMT4RR��Z¢��Sm0��FqKWva�t�+��8#%��/l���8'p��h�v"��#:@5�f��(�Z�J�R��[Z��v̐f�6��[�F�r��by�Ϯ�&یn\�+��-	�D^H�&��y8mvm�Tx�H���SM��r[��	'�0b�s\&Y]
�G��Z��gQK�cn�a��t��@���m��e ��n�`�y�+^n�%�o9N.6��s�i�{�{��hN�2@�II<K@d�!> 	$!���%!7$� !�	��Pd� h���=���'3DZ=��h�q;-[j,��( ��f�'36ŒOp�5��F,&w]{�x�;��kY��\��η�|�נ+�C��]ݰ;��i��(��j�'2,�
��sX{��h����`~�b�D��}΀��@u�u�70֋�@�A�\���W�_��������y���I'�HD�'�_�}�œ������-�-D�|�}���}0�$��>]�{T(�P4(�桿E��nܹ���w6��V�{�e�yڴ=�qGD����ޮ:5�m!��`@BG;���ھߎ�۫���k�� ��L�Pi"4��,4Dh�6�I�s�i�g7$����5�[[�A�[]���A�$�n@�K�l>�a��ga�+�L��Y���Ҍ4���B6n+9|�������d �ժ���%������
��.w�a�t��r�qS7��;Z��j�ֱ�30s2j� ��5�>����u���,׋�K`r�\z^��1��Q:�Ρ��B��H7�-�is�s������ �C������lZ$�ْ���CMJY�l��x�{;6����&�b9��BA$�$o5���_�����>�h�w4�y�E�]F�(-��%j&쓝��{@
UP4���[��ug��d��'��ț1@���`�NC-�sْ�<�2ցT>�	�߱���O�{�y�刄Ӕ�ڹ����wPr�^�}e4?�~����~����}�!#n�q8���)�6k���S�1�4�DP���mF)smeFe��߾� �����e�}U�&�3My�~?f$�{ a �H$	,����w�/��[K�����Q���+,��j2�36l<Q�:�mȠ�G���ݖɹs6
	)�е�4�݁۱Ѽ,S+�<{�I�	����v��[��?��s���|�	!ka;������fX�I�N<�P��c��B���P�6k�JIɠUn�*�Dq{t�$�ri�O=��P��tkԁi��"6�+$�p����X�[��h��hg��ԷSi4���/d�VI��lY$�e�|�se� �V	���i�5�}��.�����4�m:�B��6��e`�n�G`����s������πo��6I�X̶y�p���*�)S$(kMcWP���ʭ��{��z�wP}ϋ����>a��4=i�D��;m�l� m��ӘnUt E���A�	b���C��so�}͛WϽ���'f^��i�M�	�d�ZI�6I�1�l����
�	ffزI�b{h���L@��we���b�84P }TMߺ!$��l������O�>o�����ݎ]W�����I9��u���[�.�t��A!6�q(`��v7Y�w�$�������~����κ̽���bɻ�"���kb���T.jt�ϩ�y��-��õB���>�}���"u6�����L����빠}zS@�9�p���@|Cy����6�wZ��2쟱���>��*���	uw��A�>.��9:� ��ou��ihm
��~ϟ։Շ~6��fX�O;���;���j��F��rS@Ɍ�����$�����=Qba��F�sPo�'9?�9Hrn��'u���>��'�1<�Af[���F�O���A�/cQ¢�I矎Z'�Ɇ�'�ǛB���HB1�i{~~w��S���f�sY�8����h{��x���������]� ��@�#�$@�����qB��vV�df�;�>6I�|�Ő��P{�e�Z2��5��63Y�_�?H`H��I�w_?�6���O��y�e�%�R4MK. c�.)e�n+��2N��.��X��-]��2L�Bˋ�"k=���<��yǰ=n��E�3� 61vy��V��N�;�������x;;E˱1��;������-�%k ����S[m�ι]��6^+?�{��'EU l�x%����ջY2&��w�ށ�i7bT��d��r��7b�nl�D9���B@d�@�߾;���~�����ܮ��]F�Ŋf�4�$��GLja��L�ɝ[�>}g��y���9��'�
��F����'�}>6�ؠ�<ش�RB,��n���'-�<�d�����W�F��h~�K�BjK�n�n�Nn��Y'�x]A�t˨�l���,yF�jsL.D�r��
P j� ����>Ͼ���n��uE�u]R��3H�7�ȢI��:�MHz�	XG�@�^Z�X�x�����~_+wt}�Ng��I�̶{�)z�E���䜞wwbk�`t4��n��G��:7X��;-�
�v�u9�m�{e���Bx�sqF5����+��7<����hb�zsZ�d71���L`�(�kZ8J��޶h�k�)�����a�������� [qn4U�N'l�/b9l��j�/�U�wt˿��~�-��	,�R��F4���O����O{�e�O{�,����C��㰐SE���Hև���1�7�$���Y'�؎[?ʡ@
2n�'�����doZ��$Q�@��Pc�
�%(Gh�5�ҕ��ˁ�RrC$��~���o�I9���`}^u�{�+�"��7�M�q#�*3��ka6`�gp|�}��I�0�'�����Y'���d�w��В��˸�WP˄���,eP�(P �@P����oج���2�=��a��by���f�ȓ���]`w����B���M����s����>��x�(�n��q�F���f���E�ώZ?W�쿾VH�>�d.�Z�����>�)MdԓƖ���I8Њ����݆��OTb�����U�y�]`{��GÓm\Mn�lfcKV�K��`�Ɩ�rK���'�����ץ4�٠|�"�>���&��=�mC`_;V��9�A��}����<��VOH���i�iA�f�=�A��矲;7@S�$Pg�I'���7���v�w_�����㸙��n&ށ򼋬;�PU�@�t˨��;��%5�Z	�(���;V�ɬg�@�	�����l�Ƶ���t�����{��够��>�O1��G:��"Ik�~v��eɺ5۷!C���h��z٠|�e
��]d�?Z9��(Sve�M�i�&k�Jh�R����a�v��g9?�BI6�������{�a��n��?��5�����Қ|��Z\i����7u�V��֭��@�� �( �����n�����u_|��m~�$�w���8p���3�ճ����]bv�H9ۉ:��]�QǛh
.\����n�rcE��*�o+0�\{1rm�W�Q�Wv��USN���9p�0�J���5���ڙ��!��l�	h�6l2�jE�T̋0�>��1��F����Kd�b�O�T_8�k�ʑ�Xͪ#H��K�0�[��Z���!� FBw�ߏ��_�kp>��h|^����)��D�2̨�����Zހ{���p|������{��{�V��!ڹl�a�'�>�o����T>����w�����Y�Q�W�1EɪC�8×	�fX�Os����%��/��O����zWT���Z��6H����|���=�Y'���l�����>���4��1A{ڶ�J��@���{��9�M[o���]��s�6�I5\s�0�%��0��{�W��>�]��ҖH�<E6�ݴ*�>�"�LxJ�"P`�%��2FBa�����b�dԂ p�	��Bߛ�/�e�h4��kkv�Mu.R ������m!5s{tn9�S�/\/\D@*��`nNݻ[��Wq����8�<�x���&'ƹ�,8�J��.Z�UTU�]���ĴLF_�pN���V��c�:{S�c���̮�u�6����W��'3t`����-')���<xٴ�nw&�Z�k�7=k�+���WL·T"@S'<�$Nx�f5�����	��y��W`Ӥ����b\��5r@[dU���qa/.�wnN��n�x��Ԁ�Y������׏Y�;�Ḷ�%-l�rv1�Ɏʨ�p�l7 ���6�5ŀ�i�;"k�:GJ!v�-�*��`��Ziv �$�/(g^�e�����{�ǽ'���IA	Ѐ}$ tI,��C�@7�s�T�p֍�
����Mm��r[my4V�-��6��M*���0��aaj�����l�%fx�1=\I���;r�a:�f$�l���W���K�T�u�.�@�������|����-�PĦ�����}�-��3-���h�.�y  ������?�"�����,�;�������X|��u�s�>;.�27�H�"y�����{���N���I�̶Nu�f��u"D��İ�#@�V�3����g�7����q���ea��,X�d{֪�n�^]u�:�aBM&�ob@�Q��m0AI4Ah���t���ͱ�w�P�wPz�w4>�.�by19n�V"N���+�q�h MUDDA	H�b�( ��E�#"� 1����AQ����H}|�������o��/9�Z�n��&I��L[�� �������䭿ۚ�t��e��"-��Vc�Fnm#A�[84P�<�vk�8�0�*�G{�q&��+}���aXV>'�e��q�����<vc���A��G��<��%#;�(vh��PI�䉮��F���q�fHн��������
°�/�\�hq��V����h#]�#&��n�||p |�+3�2��6i�1�n��1��
��X_}����4¤�_}�k�q&!XV}��pBq�IP�<ͱ�+�h#^^:��MK���Ne�c��M!XV���ZO����=ϭ����aRT=ν��q&��+;��
IXT���-̺Վ�7g�ͷt8@�R4�Ni�a�%C��Ì+;$��Jlh��c�(d2L�P�d� ��P�>$�s�0��s��q�aXV߻��	1�N}�]?5�f���v���w$�W�$���~C�1%B���F~�C�4°�=����8°�hu�f��4��!��($��C\ָۜ���É4�aXy��]�8¼��ӽ���ś� M4��3s)�ї-L,�y����'ӅaXV�^��8�L*J��}�v����}��3"M���q�(Sw�7�ŭ�8̲�4K+��b���IP�;�v��8�0�*���ڇT+
�ϵ�w,8¤�V�F����F�M"����M]\�8��+=u��`q�IP�<Ϝ��CL*J�����IP�+�y���DR#�Zކ�f�|/������8Ì+
��޻hq�aXV�w70�+
���ϻC�4°�>���ڇV��g�q̭tl��{8k3Z�Ì+
��;��d�aRT>����I�V�����08�Rr���'7zR߁�[.es�`ٚ!�Tl�4�k�*�,�2���3�t=�xi�\���vn�wt�!@v�c�p�÷[�Y#n-;��5�:{7hJ-�lvz�]��ְ8�W���V�e����׏e�Nۋ�b�����Ut#�*'+y��vN!�A��iP�*]p��9ˊ��F���XV�g��T�
��-�G�XC����R1Z��P�-�l��w��C�h")7�o��ĕ
°�=��XaRT���l6۳g�&[���I�M���W)nu���es���ͮ��aRT;�߳��ĕ
°��]�aXV�~ѝ�0�
°���Ohq���sb+Z�DŎ	��5t8°�+3�>�0�
°�߻ͨq�aXV�}�naXV�{��+�h#Y�5 �ju��r]ڑ��É*�a}�;��q�IP�/�_��q0�*}��6�ĕ
°���H�Dwt�4Hɒ�;��ֲ�p�aRT=��;�q&!XV{��wXaRT+3�>��J¡��É*��>����C��7|�x훑#`p�F�4��il�%'��ͮ�6
�����ٓFY�NR�3K���;�߽�]�B��+�׽�8�HV����P4!�ոRH-Gc��|\�*y&��Ho~:k�ܾkIK��u�����v�i���F�%�7@�d1����ګ���Ƹ����l���׏P���GV�h�����R�����I�I<�<��M]LÖh���l�V�34k=XV%C����Ì+
°��}۲q
°�=����?���HVh{"/�4!����G�j%,p�|�x<�7p�
°�<����8°�+3﮺�b�a�w>�0�*���}�8�0��:9�3s�k5r�k9�C��M!XV�s���*J�a��]��8�e$@�wﻨm(@f��ؠH�3�`�A��k�����y��w$��a����*J�a��6���C�@�0�_�u�0��߿\��Kt�[8�|ְ��aXV�~�z�a�%9):�����JL�R؊]2���-ll�Vԩ�}��߿Xu��V��ﻭÌ+
°�߮��C�+
�;��D��nks�]�6^kq�H�	acu�q.ԗ1���!XVwY�s�*J�a߻��'�%C�u\��8�HV�����h")�9�l��8h79�ۆ%b��aRT=Ͼ��8������0�9�w_���%B���w��ÈV%C�����i
����MkE��B]�g�iFӰ8h")���s��V�a�z�ݡ�g��ÿ���p�
°�?w�����±���n^�l�k�˜���:�[0�
°��w�p�
°�<����8°�*��]u$�+
���t�aRT���v�.\���s+y�ջ'�)9I=�M��'��INJE;o���j{aD硸�mظ!�M��ch���r���l��Dhf���q
¤�{��wp�M!Y���Ǧfl�xr]��I9������ū6���E?�W.�n6W@񠈤@F��oO���%C�u_��q&��*{��s�*J�a��!��go�����nX��|S�]�j�p��hV}��7'�?ʆ��
��߷��C�*J�a�:���a�%B���[�h#^ڞĠp5c��|B�!P��q
°�=�\��8�HV��^��0�/���%��DbA�PB�
X$a
K0`�B5����Y � �(1�$>$��M͡����;�V%C����8�L+<���Q�^�L�7���S�xrt��!1��~��8¤�Vg{l�CT����tC�1
��a�~ׂE"=�|�"�,;4/�J�q���m�IP�v�{C�4�aSw[��caJE�eZ!���aX�!%Q8dm���*�r��O��EIP�=ι��CL*J�p���8��5��n&�r�q�&(��� ��v��6�!�w~ouIP�<�U��Èi�IP�����aXV{���aXV����]C��4�ihcz)����Ƹc&�0�
°������� caX^�s��a��a{����8�L+
��~��8¤����k�
:6q����39�d�aRT;�����M�XV}��ZaY�Fb�ߵ_߶N!�%C�h�ߨq&��{��r�]V�g\�f�u�*�8¤�V��]u��%C��MÉ1
°���\�
����@��q�s�*�4їP�:�Vq�qӢ�.�V�QM�S�fxr��gf� �nXMϮ������^ Nx�sB�qO��he�@��em�@�uڧ�ʻ�hd\��λ/F�[��v��ڙ¶�i��������}��9'>''��٦��F�=�P-��u��i���a��aｻ�q�aXT�?���7FX��E�p���d��ƪ۝�$���߿��D�aX{����a��a߻���S����柶GN�K�w���5�IW��ùy*��y���{�Ⱜ>�Fw�8�HV���7ևT�
����݇�$��aRT;�~��8E25���a��|��姬�0�*���׻'���l4��~���$��a��\��C�*J�a�z�ݰ�aY�ߛ{�T֮�8�4ow9u�7[�q
��߻��C�*J�a�{s��C�V�a��3���aXV{���IP�~�>��pևgozr�U�<.Ì4��X}���a�*J�����V�a���]�aXV���;�I�+>�u��.�gfr�V�1��sa���X{����8°�+�I
x<yR�xW+�Wx�s�9�4�	�p!<F.'�|gP�V���z{C�1�aXy�^�[�V���ow�]l�����6�el�j˙hs�ч����JܼF���Z�'π�ۉxI�v�6޸�\e�ҕ�<j�x�v!e��e��,��q���U�ֻF�f��h�^�xIӒ��y���m$�V���}�`q�IP�>�{zl�CT�=�y�$�k7DKa.�p�㻉I�*�ᢤ�V���l8��3l1%C�v���q&!XVg�����
��Xw���p�h��u�"�+��H>Dn��8��+3���8°�+}џv�i�aXy����a�+
���k�4��{^�BT2Xᠮ��u��ֲl8�V����ڇV�a����Ì*J�a~��vN!�%C�{w��8���^�K�m�l��e�͛�u��
��Xw={ݓ�h��<���;*[��ӏ6(j\���kv�b� �����Г�J�aXy�����*J�a��3��8@��5�9�l��\ 7�>&�%KhUttq�ݸ	F�{���+s�����
��X}��޶CL*J����7$�V����ˡ�A�������7g����0�
°�����'����{ ɶaXo5�sp�
°�;�����0�+��y�0�+~�r�gs\����c�5�Ì*J�a��;ݓ�i�IP�߷��8��+s�����
��X}�CL+<薵��p��wˎ�l+6�@G�*c�����q�IP�/߮w���
��ｻ�q%B��=�s���8uh:��c���Ӿ7nt8�aRT;���q�B���8���vi]gn�OQ�*�h$�dn�D���n���R #AwFw�8�I*����v��
³��=�~�F����w�՘9�uK��v[�f�]{���NJrS�ߺώ�V�a�ޞ�qaXV}��u0ĕ
����0�+:_j{��]�	�\k�X4��+s��u���aX}�۸q�aXV���jaXT�>���q&2S�ߧ���\/g�"��_�7d��RT+}�}vN!XT�s�>�$�RM���#PX)���L�)8nQ"1B.�
�B a&	A� � �KH(���$�E<������Ra.��1�I�(��ɔ��CF�0L���	�f��)%��$A&, �B�Ő��$�<޵!0<0@P�2�J6�I$���VT,B(�$���p���2F��B@�J�H(
��$� V`M�yn��B#!�$%�ߖ��p֠�
Z�!ۭ��7�X��dWi�PP҉ DDDD�Ԡ�T���.{s��ș�'�oM���\��/�,���N��Q+;r�ҕ�=�p�u��He3�{
&ܼ�N�q�m�6ZN�l6֣z�)zh<�'E�j�p���l�H]-�U" �����""""""&H�)w6���<мO�)uy�N{7l�Ѥu�=��h6 ��e��9�kY#��'�Y����]���.;<�v9Y8�N5kI@Ii]l�)���]4F
��p��)c)���h��b5��� [<t����ۧ��-Z�+n0�c��9�W��݁�O �m	u���j�K�];�ۈ	�#��pv��H���mԻ0t��j�XZi1�U	Qބ��؍��7��gR��69�x]�m!P6�W]���.*MF�y��(���и0n �k��&�Y��n�8 j�e�#ZbcB"Y��DVj�����(���G�g�dƷdr����d;n E1�^�wlX�=��U�W="��Č��n�ќ۠͹Ŝ�q'g�8���h�f.��3 )�5.K6��t�!�WY\f���"Hԅ���ܵdp^��Ŏ�tr�N�Y�����,pd�Lm�p=½0�]���h�j��'�Д��*��ِ Gn����#�ew��I�d��Og8OIȒC� rB`8B�$��`�$ `|I$��OV������
��Xw��ݓ�h#^ú�"�K������b�a~�w���
��X}���ÈV%C�����i
°����᠈�Ffv�%�c��._,�vmӫ��
°�<��f��c
³���y��T����b��܂j�&2bl���.����t4�F�°���]�8°�+s�>�0Ѡ�n�7���p�NZ@�8KF��kW��M���3�OJrV���gvN!�*J���κ�b�a~�w���
��X{����8�h#^��iM4D��K/����v�!XV�Y�s��f$�+�w���V%C�����q&!XV���E"�t�Z�%,p�N�E����+
���z��É4�aXw�g�s�+
°���Ohq�0�+s.j@p�F�5�p�%�b,pВ#v�qu�q�aXV�۽v��
°�=�\�hq��V�}�{w0�*Oy�s��yߗ|)Quauk���1�͎v䇖r���p�ִS;l8#N�J=)�ʶ�·n��e�p݆�X"s�6��s��˃��Bc`���,�)4Ysq���m+�4-#%�La\v\���sm$n;�W/.���4iu��Ia'6ÿw}6N #A�lgS���N+��q1aĚB��=�_k�C�*J�L�*�{�8r:�.�3�K�!%D��6$W^���h")�:�{C�4�aX}�㹁�%LǚQl��C���f�D(&`4ޱͰj�<���+�O	)�I�I��o��ĕ
°��w���
��Xy���ÈV%C����'i
Ϗޖ��Q�O;�{�*��O	�IHV���jaRT+:��]C�1�IP��}۸q�aXV��w�0�h���e���B���� �
°���8�I*������V%CϾ޻hq�aXV��{�0�+>�u��.�gf<yy�kNa�q
¿�1��l����aXVg�w�$��a�~�!�%B���lW�F��[q ]�����+���I�+
��u���8¤�RNNK�����S%6�(G:Ja��Z��+�\�U�_9�����g:��T����w$��a����%O���Z����s^C�`�+a
,���<�s=�e�Xi�R�⣝�#���(Q���B5t]��tl���m&P�e�P�+�D&*�9q�6T��(е�W�9'���'�c�ʐ
��`�]i�~��*J���{�q&Ь+�~���%B����l� 	�aXV�翷0�
�������p�w�%�F�B�p�F�4�܋�a�+
��{�]C�1�aX{���8°�+3�>�0�
��m��GL����M㯝]ǲxN$��'��;T�
�����'�*J���w�I�+
��^�xP�
���2��.�[���|�y�֮��8¤�w=~��ĚB��;�پ�8¤�V}���XqaRT=�_=�8�F�m�&%��!��J�᠒T+3�>��
§//%�kU���g�2��;��ڠ��d!h]g|^�@a�h#C���p�
°�<��붇V��{ۗ�׳Ñ�m�<�Q�,�$��uu�ƸS���va��a�w�p�
°�>Ϝ��8�L*J�}ѝퟤ�GěB��?}���T��Xu��͡c��9k���#1���T���f��$�(�$��I �C�!��������8¤�V����'�%C�����ĚB��=�v����c�ռ���a�%B��﷮�!XT���{�q�Ь+;�=�ĕ�B��{s���$��u����g,4��p�4,�DR o���+
°�o5ܡ��aX_~�5�CV���织b��|e����49s�pH̗C��4��kC�4°��Y��>6���k�L)���pYx3G�3U�%��;���懬+
°�߻�d��aXy<�h#Z���NCR�%�%�aEu�ƈB�a��`γE��a��aX_~���8¤�Vg�{�q0�*���ퟠ�&��+{۟�P�
��o�_��kZ����9���n����i�IP��|�q&!XVg~�uC�*J�a��3�CL*J���gw$�+<��sesWZ5��3\˼ռӉ��
��X_���l8��T�;ݽ��T�@La�/����8°�+�w�8�L+30mā2Ec��.rK����4�XV}��Ì+
°�{�k�q�0�+��κ�c
°�>`��F�hcz$e���vIg���\C�*J���z{C�1
¦��\��/���)���A4���G��%,�ds��k���須�@F����d�aRT<��ս��LB��M}�n�G��$���{�%�;+6�ٜ�R���m�O�%')%a�>s��!�%C�����b�a��\�
aRT+��>��
ǽ�j��n�8��m..rna��a�{�����aX{�|뻡�aXV{���0��a��w����Ѹu��
�8hI��8��.����a�w��a��a~�>��8¤�V�G{�q0�*{�����@F���f4c8h)��>[��l8¤�Vϯ��8��T�}�^�I�V���u�P�
��$�Nr�^O�(_�Tl��v�1��6
������K4�l��4��V�����]�20Y�GLFpEH�����<��5`���\p\80��۳̪rr�lA``�^<;�un�t��dt!�1���GOn͹"�KA���y��L�g$��rI�9>���>�C�h#]ǚSL'����G�'��kp�LB��=���(q%aP����:z��$��W(��v`�.F�j4�矾�����"NRs�׻�i�IP�}�u�q�aMxn��2�Z�Ċ�H;I
-���-6j��OJrS��>������a�~��q%B��/�\��~�>0�J�a߻�~C�0�F�o�|!E3��B��d�X0�+
�ߵ�u�'�+
��~ޞ��LB��=���q�0�+��w[�$����D�.���Ӻ�9�&�
A��v����/�P��T?0����d�¤�{�����ĕ��k�Av8hK�|6����
��X}��aRT<�{{�q&!XV}�����*J�a��ޞ�p��kh;	q��8冋\���M!XV�s���+
¦歷���	N�PY}���q�+]��x���
���ﵿ����NJp�}�k�q�0�+���p�
±���i�f�gf��yak$E����b�J"B�)D�	 �"A�0�4d(��I"�ɧ�Tf%�M�6���v3�5B�Ʀ �,s�m�j�Ɨe�;���Ob2hַZK+����PS]=�:(R�&�m�Ǉ�[,]v��\T~I���%9)���n��C�+
°�}�u�q�IP�>�G{�q0�*g���I�V>{~�B�^�M���oz�/d���$�>��;�qaRT=���m$�V�������
��Xy����Èi�5��)N]p�|�a0a�"����;��{�0�*���z{a�1��bLC����q%B��/���n4��n�ی6LK4��>K%K0�
�!"��}���a�+
�����f���aX}�w��8�V��}�v��
±��ֺ5��gkzN`�+��T�
�������4��:YZy�-t��;\K33u��iR,qs��<���CĘ�aX}�w]�0�*������4�Xq���Ⱥ���'�V�����x%�E�~��J�aXy����T�
�����Èi�IP�����Ę�aXy�}��08h")�K:��Վ|��-+d�3p�%aP���p�p'��`m��_��u�q�aXVg���`q�aXV{��u����^�E���|K��2�p�dh#C����a�*����]�8°�+>�}���
°�<�]��8�aY���MD�|��e�bX"�	���λ�a��
��{��V�a��o]�8°�*�n}�I�)�^��'!�Gc����\����X}��;�qaRWe���Q��e>��+k���l���2��[�b�@���F�w�@q�IP�=�뾻'�+>��=���h�焝��	债��lƺ[����e��r�p��4�܏u�8¤�V{���Èc
���z���8�hV���;T�<����攂X��9%�p�`p�F�4���>�0�
°�;ӹ�q�aXV{��u0��a��뮡����1�}��Q�+4/��x�2@��h#
����_�0�*J��hϻC�4��x�-�1	,?d`"B1�KBI6q�0�u���0DR #C7,}b�@f�5�ga��s�s{r�y�j�vI�+
��{��C�*J�a�~�]��V%B�����i
°�;����*J������a��a�k����5�8�0�*�~��8��*l��wY��uip�it��N� /�u;K�\����{���*J�a�~��m0�+
�ϴgݡ�aX��i�j��gfh�]��V ]	���8��E����Ì+
°���Ohq�0�+}ѝ�8�l+
��{��V�a�~�]��V���z8�N����r��Wy�6I�+
���w��8�� f$�+�ݟ�N!�*J���n�!Ę�aX{����T�<���שGN�Gxu����'����$�����q&��+=�}���
��Xy�w��CV}����ěB��s4��nu�7|���`p�F�4V���
aXV���>��
°�:���ĚB��o|�f��:֨L<GNe1iA�s[�X�mQy��q<L��y�V)�̜uʓ��i���{��a��-�a��B��Ŗ�����Y⠄I^=�����qocv'��,��Z<�e$ �Cͷ�֩�5 ����#u��;u����3قi��"��)��"�8hr_.����kNÌ6¤�{����8°�%#S�7�
*A��-k�dtZ� �\0�=����;9�
°�=�Fw�8�HV��h���i%Gߺ�4�r�8�z��p�&�d	�cM�����xB��+}ѝ�8�l+
��u��`q�aXV���
aRT+����CL+>�u)N�1�nq�9y�Y�ZvI�+
��~���%B��>��d�¤�{��u�8��+wu�E"7M;Dc�����to5�q0�*�G{�q&��+=�o�0�*�����q0��@�L�t8h#A���.;49ȭ��Yt�q�aXV�\��8�L+
�������aXV{�xnaX��y�i��4���h�Q�c�����m),P��h{w\� q�IP��pyvWW�EsU�h�9���S1ٮȕK5;�~��'�c
����3��ĚB��=�;Ҁ᠈�A��5
���%�	�d��� �d�Ja|5k�K
ȣ#�!��$���t7@$�*a�(���%�A5�2�h�b�^H��nI�$17E��\�b�,hS
@�"]A���m�ٻ��5
Z
[*�+Ft�pmY��I#���������(�HdBR$d%�$6�e�	I0,�(d��1�DAV!�I2Tx� �		h��`�+	�`�Ȑ��ɤc���U"��-�,VD4� ��221��BBNr~���[j�iMmBkN ��el�UUA]6ʍ
3�l����n��l$�h�A��˱�z�fބ�'���2!</-���܌�%�T/b���ڪ�W-��5�H�S �`콐��F]ղqg��S�Ҕ�,"�Җ8))Ar+��es�YN�LB<8Ӹ��c�`���]�m��Ys��8����r!�7n���I�6�G�����Z��n8IƱ��d�e��3e�� �79Ep
��I���g��\�g��Y��p��%�-���L5�C�����J�h�6��	ac�zD�Y���f�8z0G ��5�\W7 .�pi6�,������#2�ű����H��w6�]��U���>rI�<���|�O`h���|I !�s������
O,w�Jٚ�A��Uؑ���^�Q�@)ks���g�	�n@�%�s��N�mωg#�H���s���|�睝����Q��9X�.�B�UuNxIӒ��}����8��XVw��8¤�V�\��CL*J���h��f�Vh"2c�8h\���A��%B��}��XqaXVg���a�+
�����p�
°�>��5��F���%�	��'%�u����+}�}w0�+
�����hq��V��k>�`q%B��<�s�(q�IQ���k]�u��5�Zr�r�'�
���uϺ��M!XV{�w�0�*�����CL*J���׻�b��~�n=1ӳ�37��S�{�6aRT+���u�ǒ��P���얗Vk��a��]D6n�llQ��>��{���$�%C߻��C�*J�a�{s��C�V�>1�e�[��/4g�$����t��úoa�U�H���x��V���o�q%B��/�\��8�I*���>�g����T����p]�F������4-�\挻�X݇V�a�{��P�oD5 %�J �2�C�5$�)6C�+�|�mC�*J�a��]Ì+
�������i�g�t(��8hr��3vͳ,�F�4;���0�*�����CL*J��wz�ĕ
°��>��8¤��Ir;4ٲ��lW4P�߷��IP�+��w��%B��=��8�0�~A1�����𜤔������F�{<97|��u�a�%B��tgݰ�aRW{�x� mXnF�A3yZ�8�E��I�{������Ĕ�<���[�V�a�3���0����۳j����>yӭ�9����0��S��I�<9)�NJr^��u�q�aXVg\��0�
°�߷��aXV����w��%N���"��C�6�L�����P��y�$�V�}���P�
��Xw�>���4¤�{����I����vD�\�`H�ȃ�I�1�m|��m�K��C%ǿ}�m^޾�l��/l��n�Z0�'@��K�ݖI=ջl�x�,Y':����#MI�,�TX����]A���Qbn�������m'0�{��c(��I�����y�X{�w4:�\zf6�����;V$3v�1Y��H�m� �U;.��t��}�f�}ˮ����Z���!���q4�;��UT�ř��>�A���=�K'���&6Hj��M��!�u��˻� 
	unvI��i�z3�'�ơ��J-�9��>�@��L����4/$���Te%��1T�j�k�<͐[b�K�^y�J�\�3ÜN�]u�����=\��L�tl�c��:�C��%���UÞ�LO'S��}���a�k^ygA�	B@�:
���;�0��b�����v�r��Y�=-��@
UP����n��#I�V���ôm�z����
�G�y��)���jj\�(�8�X1L�L�9�����_޷s@/s��:��eɌ�I�i"��a$w,\<�1�v�s��ϯ�@>�Xu�@���]G�*Ȓ��	k��^��Y�P|�.����Z���ڊ'��7&I"q��wPr����Jh�]u���%���T�)#�>�&]A���a��z���cm��-P�-Y�v��F����﷠u����-+���6���H#��[U���S�~������<���:�\20Rl�g��$I �I�7[Gf+��R8f�vہ-9D��I��c�u���](��Blrn��z}t�*�G�m&��(�h&5B�e��NI;޵����+l"B�P�
�L�'����Y�}��.���n����!9�{��
=�f]A��Y���<�d�g��� )!�u$$,�n;l$�p�-��<�$��z��lХ+be�CE�j��{�-�W��>�e�/%�Yݗ�T��X�b�z���<K&k��u�5Ov.f���'��D�Y������sP_[��ϳ߷خ�sgh^�\��4y�LI�I���'�����m�@����=�����⫉���h�n&���ڼ�[��� �����4�IXtI�A@	DEu��(��f�J@H2�6K@���M��JE��Y ,E����H��@֩ �0���U���g���'=�d����E=S��6��I�68�����h�Y�� Gun�'��i�p�����M�qL�I�)z���h/%n����YԵ�MBHi�	���h�wPi�Q��ѵ,R8ŉ�\3L%s�jJ��T�C}�߷���.��u�"P�$ݍ~���؂�fTXG
�AY���S@��[�
^��e4-�k+��vD���=����X}�����y\�wp���jݘ�hٵ}��~�W�_~�l�HnH��XH$�$# � � 
Co�'Ɓ�<����2�x)��d��e�;@ ��zl���m��1�l�{��e�����^jm��z�.jt�ާ(P�l�5m-��ж樰����������ꮠ-V�/�9�ۃ͋EѰ�,1�9�2�ʰLf9��|�����y��O3&����'�V�s�n��	f�F\M��<������d�_�:f���d���#P�)�)&= ���a��e��h�[�ϯe�$���)f���Ul�9�3-����z*�/�L��rME ���e6�m�.�`��,�V֤�d�h�vBa�e�(��/8d�]���d��e�7l��[�������HhB��;B�&��!-��\�aA�!y��q���s.8�=��v�"�I��*��Nw��#$�o���>��ŋ�G��h�&lz��b����%
[˒�U.�6db�I�Ƥ��W�ˮ��ԙupp�"K�E�`�d$o"֡i���e�ס���?_߻��.��Ul�>�-�|z�#D�7d�5HԏP��@���X{��h]��u���Qɮj�8�$�^ɗPyzנUn�������TAɫun��I�@����t˨z٠r�nk/b\1L�)7�"��}�t3��TɉZ�$]R�L��k����n L��{~���.L�������G��%&��,Q���=���f����G?��-��}�R�՞�g=L�v�`E���rQ��k(0����S�S۶ܱ�Y����p�$�f3ü[+�Y�6Q�ƚM�cNMa��4�+f�kκ��t˨ϻP�)�n��{	�r�nkz��˺� �u�w*��P��#�m��ij��z��h�]��R�Y���;�-5�{1L{��P{��<��z��.��A�&F���M��&�-�4��7rZw��x$�u�Ԩ:�9�9&(�����������:}��p���{�4Q-��E�?&��b����:����@��.�>�YN�ZnF��M2f�\1����t}�BC��F���H) 2�@����=�j�Y�}�L��q��d�qn�D̈́���l�=�u��-}V����6�MZ�S��b��V�^�=��Pyw+���Y���wQ�f�Ϟ���?�9��[���A��X�Rb�u<�y<$��Y1���|���h�]�'��Cr6d�wmm
�b�`�'��1�u֦���¶x������/t˨y[�<��zNg�bɫ\K6a0��u��hz�.�>�̽UQe{�S�r@�v#J�>��ٵy|�3��Vy`4�i��$7���DD�,�d���
[,,!Z+TYGҒ��0H��"y�@Q�kL�jI� �D�	� a�XF� ��"3��� I�!&X�FCd!�	��X�����H� � ��%�i)l- �h7� �8	!��J%���P��"`5��x	"}H�����!�vcn�s»�Сt{mw +)�vH���}"D�$DD)�������n.������;%KP�Z�zR:+`�/�Xn��q�]k��[�G�L��v]9��CӸuclF���u���r�1H�]u�$����mu�(�Y��DDDD@�2D@`�	:�Y�t���������
<h�`c�x��Lq�ʬl��	*�ʹ-`玂Q-uutlFk�v 8	�J�)��8��	ؖ`|���ua�κ�[S����v'G;{s������.	�l���@٠��z��7G�ڷ'nĻ%7K5�6��B��'\{i�[���A�� ��	�-��6�st�i�kd�8MʣYRiR�M3p0��s6`��0Z(�V���i��n.��<H3�	�eʜg�`��.�P�;/<��)�^u��; &�ʏ4�}gS��1��r1�g=.cΎ��N���j�:G[P�0�S�:!���}��9D���Kd�p�k�t��&�����W9�n܋��g�v��'fBlh�f ����e%[��2�r��j�`�4]�*F,�	��3ю.��m싆L�Vpb�Y+l͔�2\��p�1[��&.3��P�Б�q���˸�]�����ٹ�r����.o�@��"@'�O�!�IRHnN�I����H@� �`nI%�A��a@��k�חj��>�x-�2d���V��7�/u��Y�P{�e��f��G7[P{���j���/��Fbn�n!T�f�p=��4�c�\'k���mM���0�۹�|�[����I�9}��)��nA�%:�A��7Ln)�^�M �]u�������SC�J��<�I[������ܥ4�V���g��,���z���f���j�y��
������}�I�1��r��Mצ]@S��7X�i!����#9�ˁ�l�,��:[Q�&�5Σs���ޖù��zE���^�����tY��5��xv9�6<!ظ\���[�q������=l��S1�1A�[^��e�s�V�)�A��v��2�hPFV���:�>�����x��M�q����O;��5-�Fe�!�����gH��qc������:�_5u�K�����8�M�Q��&B�r����WE]M��V�/Ma�t����Q֕5#R[�f[NB�2�=�)���H�aݶ����������:���#����7�����wW��Xyx�k/bS��'���Q��]@x����)�|��Y���8�Rk�n]���=}:���ueq�mG�0`MKs�\.�7E��3'��5y���wW���-Q1(�����2j�`(�0QE���9/8����2��v-1-�ϱ2%ƶ�-�m�#�Цp+66��!pݥ�区
����.l��F�X�"�upr�v2M�G�6�Nr}����烦ڠ�)6� Z�89:.:���YM�ҚO[��U�<�qf��I=dĵˋu��+u��e4�U����LoĖ��$���*�+��f���SX}�2�)؎˓#kuĔZ�C@/����t�>]k���Y�v\I܃sb؛5̃�z���hf�q�&�6ғq��m�M��7���x�d��}���U�����z֓�)_���"�mꃜ��0�	Lm�6n���.��t��_+�~�����C�i��O߆��������zϯ�n�D$H��$Y! � 0` 0!@��$5����'�Ŗ,���r�
��=� mC��ũ���:��yw+5���.��t���q؛DQkز'�I	����� ��d�z�u�$��2�=�A��z��T��=[k6D�@�ź��a��~��➹�R��n�#��rCs1���w+P�Y�r�Vk=�Y��
V���M��#Ǌ!�$ǂ�A��M ������#�(�OVn�'k�^��-˒"L�#v��r�� SG��4�'W��q{�/hP�����`��jݛn4ӲN,͒�<̃-R��x]��I�P��e�G7[Pz�c�cؤ�ݝ �7]�OsvY'��2�ڪ �j���ui!h��N$T�#p�d��>�{C���1K+�6в�Hت���&���b��}��{��˺ɠ}�2�>˕�Y"�90f5��#R�,�cw�-ˎ�9��d���9l�����q�{����#a�`Wn�َe�y�Pe誡A��ٮ�:�wm�{�<�{�,,06��sHG0�@��˨=ze���@�܋����L�nǢM�nj�h���n�<���kÂ�	 �<���C��η�9���b��Yb�ك�9��h�V��gT��Ü��ę&b�,Zv9�f��J\���\��[�Է��s�g���vf��Bn�(g;�̼��ʶf���0
�ܜ���a���	�rYB�4k\:��sB)�e��h��q� @��u���ʫ���4Z,���l���ن-���cv����	&\�9℟�N>���@�f]A��{�}��{L��7[��q�1��Ɂ?9�McR�E�U�E����l�>�e�~�;��h��R��m��*��@��]a��.��wY4/�%i�<�k��y�Ǩ=�2���h�2�y�uԲLo�6Gt����O3 �D�qA�����d�B���ۮ��F,�,�Z'���W�9�����ZaCWU��V��x��¨`��g�P�f]@_[4;�lL�qf��H�ۉ���<<��.�������v�ڋS���/H��t��^Qi%Z(����l�YТ�%zLE#9z�c�޽������\n�����O��!5ɂ�<�����u��h�S.��91�wZ&M�$j=aW�z�u˹Y�>�м�ȹ26�\�ި�M@_+u���,�<������(w&B9�h���3@���u^-�zנwt˨μ�*�)#׬���5�wJh&�x,����Mm�rl����ő�
d:�e�yu��e���)�H�ɫ@	L����\풴Ң���߻��<�d�O{����^;�φ�zҊA-ko5����W�}���5 IBC��%���l��צ]G�q��C^ő=�HM�_u&���WW����#�{h��ݖO:�̊8��cQ$ݸ��J�[�*��@��P|�[6�5���ճXn#@��.�ų5�-���9�z07<J�ηc7���&������&���WQ}����l�^㦵`n&c���
#�A�G���@�Z�4�[��
�P<�h&H)��-�4��/���-�Қ�V�/�9ٍ��V�ȵ�"���W��wSH" �P#D�8Iaڪv}��d�{1زy�	��q TՍ8������)�|�[6߳3?+�/������BE4q)����w���Ӷ���ei�˂P�̵2��L���F��~|��w��h���e�a�&�-{5��|�۟�RL��� �;i�|�׫����Xr��a�Қ�*��H�l{ ��u���hy[����}�*��dKvh(%�$���-y�ykj�R^��b�>ׇmʫl�ɢ�a�R���S@�ο}�_��_�^�H�2�AV B��Ns�'���6�ʼ�X[m�v�efk���<�v4*��3&�`P嘠ln���ƙ��h�kՀ/������a�n';]�����q��l\<q�ٺD
ެMw�aj��}�gn
����kav����*#}��}���:O�On�2c��h�E�XU㩬 �f�<��-s�N��B�ܼDZ����$D��nP���*�WQ���QA�ך� �0A�$Ł� Ȥm��;�PU�]a��S@���;ߒ�����S1)�����S@/����]Ma�u�ж�&7��&��ŋMXk
�U���4�����Y��" 9�l�@��<�Y��=����dh��۲��Z�OQn1n�Q'l�M�{�e΁�{ݥՕjX7t�<ئ��J"��]���=���O�e�}��œ��L�"���
B��@�� �d%���UU�Hea,@ѭi�V!�]fk1E�7r��Ub+xց"2,�o�aI��#FڒV@0�NBCD'��F �d&���� `�( T`�ń�#dH� 	 � H!r� (ȋKh�`�Y6V*,�$Adb(�����21�7n�!PuMa5��[�3@KT��iac((�BCr0}_/��l,Ήe�ٕ���R����-媠���FZ�7CE[)Ί��'���.�m�q%��+&آ3 �q��o ��M���(���n��T�PR�O��V�uK�+y���%zk�[6����E��E[M+p�cVXj�� 3�ˍm�q���zÞ{p�q��%�q/-���n#�݈�&FM�	F\F�n��̋"V4�La���dW�� ŝt�n��n�[�^�9�˜�Ɂ�5m��3rFŗV��J�ٖ�U�f`¡��Дf��K��n@��
��E�m�n_-�(;�,�pp3RV�4�2�Y�l h0�!h��t�`#��X>���<�q����z�zYn}xv���}����	8B�!�$�@Bp$����aa ��@�=	4	}��a�Wk$͸O���HJ#G<`C�����/&��u��o�lRj2#�:�\Buã���9f��ۡ��-o9�7$��'9�NO<oO6�`f�d�bc`vJ�V��=������u�jנ_<���r,��s[؉����[4/Ma�t��{��
��!�A-[1�Xu��hW�h��X}�2�3�,Eq�֭X�@S@�y�X{��hz٠�SYJ[�$�[�7#$j-���w@���bmfQu�HҒ�V\j1�`й[�����}�û���>��h}��`�$��#y�5�ƛ��k�.��ķ	�r�Ozױ�':ǳ��O�6œ��6�� �^���֯@=�~�t�9�O{�4޶hx�߳2.�g��Q��5=�bRG�=]�Z^-�z̺��5k��_�a-��3`F���e�$�w2Y$�W��:��6N�n��&�Ť�-�����&b�!���m˺�q�/bi�ܺ��v����|����.���]z�1��6й��(��H�oP}�u���u������4>�9ى��n�5f�!	�}ze����zנwr������w���#��l��W	չ��<��>��$d��B,BU������� 2@`�$!Y
B2I�$�/�_<�/���;=q�k$SG7d�bMǠ�wP|�h��L�����̾��C�M��-�zw)M8["ĠT�l���
�7,��e*�5	?o�;�9[^���Q�Q�^ݫK�Y��]�FSF���aDI �zנ{���w;�:���/�:�L�n͂lkCP��`w��w)M ���̷��7Y4Z�kԄ�[2���n��ֽ�����d�Lz܏E2,�_\Z�̺��V�'����o'����VPw]7�h�XwMIN����lm�$3Ӱ̻M�ĚVĔ�k��tz�-�@�cvq��uJE4m���JX9b;���5�T%�k�3�7�#�`;KV�(a*�	Y�5�b��J]�j8�6�[Q-Xmy�Ns�$U
��o%���0dHG,�Q6R��Z�+u�p��i�A"$�dH��YKk4np���mO|���z̺��4[���%i�bɻ�&�U,Ж1��]�r˶t[w4ם�_\Zצ]Gu�F�`湨ŋtK�/���Ws@=�n�8�v�P�L�&���	�O:��['�����PKۛb�'ُu�[�mCf�����X}��h�����a���h{�M��D�6H�Z����uks�Q�����C�u<u�$����t	����4�G]aW�u��b�)>�n_���{W��n�lȆ��h�ϱ[rE��g=���pG0�r�һ��ΦZ6-��貍�!���^e�ocW]�{�׮�j�m������m�[:�I��q�}ׇ�y��T8�;�l�>�@����Ijُ���w4�]u���=l��ؑ\DrkZ�1l��B��^��w;�>����8���q�Oq=J0� �V�ܺ�'���N��K�[�ϵ,	�R9vɖݷ	�'���f���\(]�C�ۑl�i�}΅������526�܋��9S���t����u��w=�k�2���ʡ�c�����	$[����>���ם���e�أ�䚵�l���hެ˰*����W!=9yp���$�掺���V��n�Flް�t�d�ެ�z ��u��h�{vœ����l�׸�$4�n���S@=�n�>�n���X�H��j��m��y�}����ݰ�gn�$��u��*Xb�"�&tf�f+��k�u�[4=D��Y	�bP� �IVQue�Ki���ܟ���]�˺� �����4>�A�n��i=q�= �����f]A�k��*�n���i=5�5�n'h���K$���
 @B��fI% �g�}��W���f���,1$9���1����^R��[4�V�[2�/�x�1�1j�kF݁z�����HFy`OX�+/2h3Y��VƆ4\/&.��� ;�f��㩬�h`�^�{���zu����p��[lM��������Xz���$�۲��u��EjZ��iGvO^��ծ�@��u���.��Y!���7�X�Zˎ���빠y^�@/+u����bY�j����UUR^��I��{��M�-;gv��Fupˁ��� �t��n���j�<�fI�1lmN�<����S��(�f�Y���s�=�1�*�+̚�J��W�X���.h6�F���+.�T��1kx0Ei��y�+���@�[g�B@�A#��@�$��]��	bx�p�.�6[��{����=�	G�޺Th��d�fF��YTA�#b�#0���*��=z�hx�\�D'4�W���R^?9�m��GI�퀲�LI|�����X_r��z٠[f�w. I�\��8���|��+k�;�e����}ʶ7����n�#&A���u�r���٠{�Jh{=q���KT�nl������h��WPUֽ�"������"P�Xk��H��ǝ�۠(��ҭ��MHj$H��h��2�.�u��FWB�C����y~7��Z@zs��C�m���.����6��J5a4mXJML-���k�m�b�jRŕ1�����y�D��21[�rrBI�����hiQ�g&��Ә�/����yu��٠z����������HŲt*�^�צ]@{��a�>���$s�JdrjN#d`���]@u�h�R��+u�勱܄�n��<K@�빠}Ϛ������u���N屺u���|�}/@�g[��C;���	,�+���f�H$q�C޽���f]@[lпm���tomo}�m^��2FqD�L��B&� �V 7��w�dy���w�q��-��`��$�ޘmP J �6O:�-��1�5��f]Gw�x,�=��P�&�-�h��{��a��T�ǋ$0�f;i;i�d���km�qm�}����Q*�bo!5'�,ofp|����3@��4Ʊ���t�fLe��Xn-GVe�>}��{�ǭ��WsB�PN�H����퐰�	�LǁWE�m�r������s@��j�
���{.p��4o[��["z�����<�����=ze�e�X$�^�&F����y��f�|�����pd����2F	Q��`"E��VXF4ȤB��R��Rf��H���4D]m3cs�M!!�8o���cM����c#1�fI�a���J����&r�������"!j1r���`�@XP�$%���&�`��(Ł� a�� pd#��� �"&��d�&��$��(�b �2! �d0��DA�,Hj�ed(�1c��AE�QEAhW���$Ԕ`�2E@I��D"#���da
��Bd42M����E!�.�,�
�f�f9�Ad��� GvT�t2��`(%�#�@�0!���oT��Yè���D����7a�cg=��U�""< �vH��D@;BOm1� ��z����xý���ŕr��=�a]�8��8625�uR��۝�:wc��6���x�T�k{W=m$��@�����NQL6-�uՓ7Xմ�TD@ DDDDtDDQD[��˯#pKy�cc��+�DM	����q����ç���`pa���J����R�[&Q�層���;B�c��k�`�s����;�]�QK��l-�ve�"�]4�/j�X�>1@�A��E֥x�/9qZ�ʰ�O�{���%0���J۸	1����-TJ��+��Nn��
�]w4IR�f
�����W��ޙ5��x6S�5+����u���[�C<�qa�����ىdF��sd3��6�Υ�nP,���ۢ�4\�]$H�L��HN����U�,[Y�1.A�d����U���hä"����	��ܙ������q���4,�3+�L�hv$ɶ{NMs������qq��YH��n�gq��ng<�vN��Ϟ�!p�͗3��	tMt�.��f��.;p���Y2�(��##�{&��L]�0z�k&7M�b�^���֛���5sZu�HB|�����$'�'�C�l��'${ �(X(�� 
�����'ٓ���&1�-RkBhok
���W�����y�SYx
�2"5��k�(#@��Pf��1�#X 8θ��f;XX�
���=��g[`u�w4�]u�^,M�B���t���h��Ќ�r��HI�t=z�hW�]AWr���uz/��Ǐu����c5��y�����=ze��۰�[Psu���4�@=��X|��Xz���>��z��'rd�ɻ�oH��r���'��h�u��f����(������ƪ�7u�:
E�Q�h���`�%m�q�z"�ٝ�m��Û��ɭ�F\Rƴ*h��5���mC$r��y.�ݥ�Ϩt�$��l=��v����om<[N6��Բ]8�uu\P ��
 M��������X�B�S��-�I,��8�4�lf3����5u��1�A$f}���z��Ku�����15^�~�����4�fm%� �uћbib˚T��?{��΁��Z'��Y�d�i�{�Slk,�qAz����}f]A��M���a��M��1��Ij���Q��Ku���4�w4
���}�g2�JM7bz∏X_t���y�X_Y�Pz���云�2$�2=Rcf��������--5�ā�!H��e�'�Ha1B<�&%����]d�=0�>=^E��ܵs���R�!��u�9:kjHjM��v��:��B�d�\[�u،���׹����,2�-���u�stG��6V �f1[Nrq��6���8CKu,^Y�������h}���h��������g�H�Ғ�9-'[C��)�_<�X|�+�����,\��G�X����k^��;��h������{�5\��ѹ�<؉&=�yn��Y�P{�S@�<�Yy.��<�Mص'��'�����x�툀���4�V�[�

!H��HE��}��I�d�`^빡���T��"���SE٬�&�c�Y�+�oϷ�D���l��<��*�������`ձ��N.��R(%�}ט��Pf�	UT
誡ACՑe�O��I���d���9�SH�[#O�{�4�l�j�%��v�>�A��`KȬ������@��]A��.����@�w+��PN�H����'s5����	�wP1��:�gP�n]�U�3��I�x9���M��h��C�s�px94�F�Ic�6�CB���F����H��{�2��j�/�˨;�e�e�X$�uȳc��O@�w+�z��>Vנ}l���x���0׳A6k� ��h]>�w^�(�� XUUw�v�Oq�+%�T�2!E�$�ckP^�P{�ج���,�tUPKُm;�blDQ��OI1��Jh� ֶ�mĔS����2p��v�v�a�9���wS@:�4^-�{;�\��n�d����
 �4�m���C���Z�ڴz̺��L����Zq���7vD��CX�wP|���/t��}e4=��N��1����9�r��@��S@�<�X_Y�Q�uuǑ(̚���A�y��<]�vI=��Z>�
�B�����K������/X΋p'3nޗ��?m=�,�.a�6�ȘO�[Q���T ���@n������g��K�2F��j�]�Tu��Lىb0bDm��4�ƻT-x����2�a&�2ݩx��i�d�L�Xj�;$���������ˢ�����B���4�Ա4l��x�ոx��o&p�=J~nL��V���mz޲��ʚ��oZ��vm���k,���xF�I8�G�w���{�]A�y�X|����{��:�jsX�ّk��u��/�S@>���\��JM5��DFށ�����݁޲��u�u ��)69��5����ؼ��zz��A򼮠�t���
�8���j1=�M �ˮ�Q-��6��Rs�=wn|5��Qa�S&�nc���W���<���S���w��z]y9'zKV�9Q�yJ�c٪n4��96RK���Q�No`{c��K֏d��$;=��y|\�a�ן�uuÜ�e��/���u����l��.X�1��I���L����ü�Z��u{��dS\z�Z(�`{�S@�t��}��Xr��B��uɎ9�Mƞi2H�,�v����L���˖���̉4ݙwi��Q��),�?�A����=�)�[�sC>�5��ɮE���k.-�7C�G翢�� V���)����~�9���b�{���@�-�����ǂ���;��U��%6�WX�M
I��/<�X}�:���hW��{��2%4�c[#O6�vo	!�Hh�Mis���������y廚�\�bo!58a�5�>�:��)�^yn���[�����'�ܹrDM��@��[h�̃m{��}��Y�Zc�<�M2!3TR�w2Œv��qY���2AF!X`��YbԄ�T����c]�/�����/���u��i䁽�����gY�Ff+V�!D�%���[�/�S@��WP{�e�_W��S�fjl�#4�s����]a����<�u�[�J��A5�˶ˁ�l��L6I��̷� �D!@B2A#	'�$� C�}��'���t���Z�6��8n�	�'��h�w�b�'���GE/<;�ϲ���"ǋu��Ǹ�Y�yx�6Hv��JP ��p2.Ѵ.�LJA(Ӊ�1�~���-�M��u�~�"Q9�� ը��#�ɏ,C�ƻK2
&�~}}:��נ{�e��w4=�uj<�dǮHٮ���n�����<����u�guuǎ6�Motǉ�#P^v��<�;�2�/uz{�&#	&��6D���빠u�@=U����2�#��S�a��-�J5��#�jF3,FJI�RJR.HhQ����h�HVH���Ӊ��p�}����H��y�#�u���k�n*�/	�u�3;�ȕ��)�� nf�����v�mrm]�m�@�V��p�J�W�Ґ%Ͳ��bk��KMV�E���Y���]��0\p��7'0ݽ+�Ѭ\�q����z�h_,����D��7�m��?���� ��`�\��`b���K�gf�?�^����Zˋu��b]���� ﹺ0Q����m�cY��-A��@�y�X_u����hw�ɫ1���Q�Ȉ������g�H���d��Y���fX� Ig��0���rG�LlZ�����;�2���4y�]g���*�"s[�Q��M��T�e�|���'�Ɇ�ڪ������r_��
"I6(�oRl�[w4��Hs�(����\`�IYL3����OP��'���x����L�fk������O�	!$���BHI'�@���J$����I��!$$�� BHI'�B@��O� c	  $!"���BE	 "@A���$��BI;BI?�$��tI	$�BHI' �I��!$$���BHI'�@���O��	!$��BI?��I��I���e5��z �5�!���������}�o�+(�\ �    8�0�8|�c���mu�p[�euҺ��<8M��")OY���H(D�@hɍˀ
 m�(�'+��'Vi����tM�ٷ3�G9�sm����V��#��DZ�9����.���� P      �?�UI��j�P        )�%J#�#@ ��#C)���U"4�        m#JU&�D402 2 14zD�))OD �4     I M2L����Oj�"z&h��FS�������D�_��G���E����^�h�� R*��������=�DQD��%i����ӟ���,Q�����Og���k9�~&�a�Q�^z�о!����l��"l�AQ+K���9���&�q�xj��&�B�R���A�����b�T�k�x. \�(�b^H�9ӏNu�����]����]]=/����}<u�;��z�]��ꮕW*�ꢪ�2�۷�m��nUW8���s��n�0�$�����[�����w����:=Z{r��|��wwww�����fcy٘��Fft_f�fvf����=�������Uʬm��]vvvEU�t����v�*�=UUUUUUUUU����wwv�wz<���������#�#ȍ�<�<���N[ڻ'�3��ww����4�c��~�aݯ��O�/���ۛs�V%$�Bɥ���DZ�
��f �s��IM�Cj����Z���ZkP�R���J�|���/�m<OzR�-ji� �E�V��z��#!y�Ĥ�S7<S%�i*�`��jĀQH5KZťZ�<HpB�B�%��x��Ԕe�
K0.�$)�Qy#D��¬1��ͪ%JaK�KB�q�ģDǙ�4��<<Cbi1Ո�V0�*�X#�"S�J,+!ld��!d`L`�VSDh��F�����H��4����fb̭G�S�T��Z���H66P�
Fd-n�*�c�[�u;G�m��ơboHVE��m��B�'��j�+e���vXQ4�RJ�	��h!�ʝ�,n7Z`\H1��V�Qb�ؕPV���U���̷��y��������
.�;��׫�����#����4^,X��}(�?bQ1��m��y�V�[r�������v.۫�׷j�hцhfU�o30Cm�u3z�I������T��r�u��e^��e`3%n�����Um=7�\�v�i�Ƨ	�YZ�w��Av�UP�-�r�u�j�m^���SG]�=��WL�Y�F���+*�kw2Cz�=*��$�'ZD:�dFm ����
��T�JV`wh�]�J�[YWvn�J����[��щՌޣ6�7W�{W�{W�z0�0�0�0�0�0�0�0�Tl6�0�0�0�0�0�0�0�0�0�0�0�Tm�F�0�0�0�0�0�0�0�0�0�0�0�Tm�F�0�0�0�0�0�0�0�0�0�����m�6j��a�a�a�a�a�a�a�a�a�a�m�6ڣa�a�a�a�a�a�a�a�a�a�a�m�6ڣa�a�a�a�a�a�a�a�a�a�a�m�6ڣa�a�a�a�a�a�a�a�a�a�a�j����ogp���a�a�a�a�a�a�a�a�a�a���j��a�a�a�a�a�a�a�a�a�a�a���j��a�a�a�a�a�a�a�a�a�a�m�6ڣa�a�a�a�a�a�a�a�a�a�a�m�6ڣa�a�a�a���pxs���a�a�a�a�a�a�ڣm�6a�:�]:v�]��������c_�E)o"�nI�UF��1QF�Dq�:�B�)!YQ-�5(�NpT��J�DrP�cS!�piY��W^;ej�G20��[�Z�eX6�T�ETQWlr!I�4�q��ln�&�D��!��P[����ߎ\�志>���������h�/�[ �8%=G|����q�ϛ������ ��$���BA�H*T�#UABC�0l@J�+"�"��Ͽ]������Ԍ��� ����l�1�,ݻ���Vo3k�q�m�덛m�+6�uěy�;u�x�n�ٶ�m�x�m�u�y��P�m�25���1���l�[E�Ul�v�b�[#�X�V�[�Ul�v�b�ZA����K����r�3� z��ȩ�IZ �Et��u�*:�M�f�EJ����K�A6�(Q��ȆPA�/p(��I>�04�a	$�������"����\�M
DB��pm��!��<Lh�M�+^�V�`72<6�m1AOI��^&������{�sx&����ww`w w w r��������� wx�^�=z{�Ww��qײ�
�)FJ0$�Ĺm��V���Q��u���J�+�
$�<������N���b�zid��I���(q@�㾋�"3!k�Ku��O�������J�wU� ����Q��o�y&���^�C3>6�uBy� :�(�\̈2�6j1IA��q�Pjs*�f<�2@A�3P�T��H#����ꄀb|����`��|�@5ͧ�{�OX��vF�H�w��a	F聛4*EQ�3#2��df|=�q� I!��J30�&](cSXIe���5qbE��]4 �qB��fB� �Jn�w��Rf��iH{���S��̦1F��  ��*X����$i%��!�55�U�E��ll��  �e$����QBYq���s*��D!n�� ���S3D�T faX��F�������'�y�l��3#2���7��Է�:�d��km�bObP,���d�)�4��Ҽw�� �侮5ĸ断�BZ[,���*$�M�H#\���޹ɻ��4��#�t�DE�0�I��z�k�Yx��A��4"�F����Y���ō  8��BHc ��/[�p֓�$z��̀ ���1�5�{�sý�?���y�&k�k.m�O�߼�K]d�Z��'�<�U�k���m��K�$�K�$�IT�I%RI$�I$�U$�IT�I%RI$�rI$��$�J���)@)JR�� ��d��]�,�5��}|G�,_K9S�wE�}�P����q�����s�3&f+loiN%���vrW{v�.|�5o~��%��[Ke��X3#2���>|=||o�������T��ffh(%�͙����ө<T3�sv+)F���8  ��~��L+���6d�ů^���+��;��߽ẗ��}c���vb�<�u8i�������� $�!S�fb��%��^��E�NN.�Í��ޟ��"#̼�>��,W�L̶ߧ����@3cY}�YQTVN�'�y�_�y
;	�k�Q��7ޟen�L�I��f�w��Y�j2M�ol��{�n�6�����#�܀fM	4(U�Fdf������zF���w���~ ��/>T��I��N�%)�a�4�I�Q���ާ�� ���yP�,��dfB�#2�^�g��LVV׾��lV��y�Yy�����f��ooU���C��3�0��s�腸V��{����mt.�À �������������ʫ�1�W��Qj�A}�>TWw�x��$fȦ�虘(M�\��Tw7NA���w��|n�y�N��ם<l�3#2��j[,/����d���;��� ,�^�^-4��c�R��5!�����cv��
5����(5�%��m3&�q|6L#b�E�{yZ^���&���$�\;��F���m�m�֣��G���}6�m�� 7�37���J��� !�C�)B�4$�BU._f-w����V�Y�.��^�9p\������ˀ;�>��z��;�;�y�u�Ι��o2�|)�4��L�{����
@�@ ����2�D<X����w��r"��`3kKjZ�R��e-�%���Y-F��`�����)��Kj�_x�e�ZO����`�Y<�I0���t�$��IJ�5DmIk��Kb�gi���E�k/>��kM�)#b�w��Fb�J"����)#��:R�ȳн��KkV/��<V�]!w}m���j8���(6<�Z�'�C��b�
¢!:�;U�"pqT\�����u^p�ZiA��t��Y�*��-��o���E�)��wV12Ȱ�sKgD��Rҝ&��H�n��(��Zܭ���X�&�[23L��3#23L��!F�*�eSk^k��u���m��xK���tmh(ډ���g!	�t��b�e��4���{Ն΋�� ���
�ưQ����g��	$�������N<]wuX��������'M�4��h�Iy��B�ߩhY֬���\�-V
q��
��sҫ8��W	-�r�}�;pΛ���%H&*��E�z�՞��>��Ց��{(���������'M;j��ܾ�,9�6鷹Z!J`�h���akuڡ`�`��
^�ɑEБ��o��F��-�i����ԫǿ6�o��t������ڒ�lQ������MV�.]�Aq��[x���ךzi��}|�:Q�-%���[,,���,���[<�?9��ׯ;�dm��g�f
�D򤀍bbB�{�[#6����J�r�����}��E�YC��Z��~m梅���t�������r�e-�%�%��e�b)�s�s� TEi��ܚ�X)!Q��J��"���t�"ȣ��j0�m�y�Hz�m�ӹ�)�$JE�r�T��
�,!�S��B���B���U�(�F!�(���-[[�@I ;qb�_i&f��Q����Ȉ�X��J%�#1Ċ��{Ԗ66|�� c i�|���|[y�,�̫�u>N+S*��XV䑻j)h�j��<I%RI$�I$�U$�IT�I%RI$�rI$��$�J��I*�I$�I$��$�J��U��z��}e�'�-��;ؽ�q�3�%�k�[T�[3�����QB�+W@�FUǝ�>�����\8�jB��V�S���X�T��4s�M�0�>;Ϲy���^[u��;#4̌��Ye-�YKb�5\n����uܹT.�m���a�2�l��I.0VYFs�E��,"�r���U��!�y� =-VY������֫%!--�%�%Q �q�*�yƅ�VG��m��أ���ٱp�'`�Mg9�{\[p����Z�:�m�P�����2��KbXl:���Zk��k��$��5��B��5��)ш��߻+B٢�z�*|��`ȇ�j����6����>�X��){ܨ�q�d��5b�5뙡`���x�ٱP�F�4嚔�[�2�{yj���p�rx�+����T��)b���
!Q%w��#�ąB٥ɕ�-����߾�d���,����)l���,����_y���/]�$�fz�ֵ(�r|'�V��|��/*�I�E��LL��Я]�J�F�"���U�l]|�m�fg]����F(Q�qS+k�X����y�ӎ�=z��)��\!a��
��)h�ٲ7���R��I�p�μ@E�Q�s+��6@f�6Ѵ���BU�ցi�M�c=0�zvl@���\�Z��S}��V(��v-w��[�m��޴�P��{tP��+�[(����VE�]6��s"�	{qM��E�ڇMP�B�zx�XF{tz[m�s[��O�%$�1�
�E����W�4-m�u8T+"дX���k��jE�|��zgUN�fFi��dfFi��Dj&jP��o����`��t/�UK�3�q:��"�F̬�=5��b��fд+����x`��.@=-m��q. � 0�o��	E�f�S!�3łB��T)I��x dA�4@�ۖ�%���0IV���۽x�S:6Uo/
������ˀ;�;�;�;�;���m��G$n�blS;�q��kU�$�/g���)�-h�D�
�$"�	D5��^4��ݺZٕ{ޭV������j����ٱ����ob�T�	a3>��,ß���*�X�VB�s��%bd�e0XGV�nfe��Voذ���3-˥�f�`�"�IO{TY�mN�������5�&a��W�*�ŒE�M99�v�Y�#co�,Ԧ-	k] ��X�X�Q�1R���b�8���h�ǲ$������X�fUϓJł�H��}���c����_'�@)8���GK`��f5��ɽFų��Jq�e�|~�lg����̌�23L�̏���&���n��[m�l�+!Χ��@2�Z�0��R�ku�S��XEcX��|���,�E�-o��.�b�A�i�����}�E�k�����ʈ����{w��hB�-b3�����9njqa.B����0XC"K����	I�!pV+"šM�n�ʌz���mt[:"�N����lY�+�v�Mh׽+-�qċ~�ꚳ��0Z4k~�F�fŲ6�����
�<R�}o]��%��s[0JLȅ2("(�6E�IFWg��(��$|IF�B�맄�5�JM#d-!Uw��
�%��m�A�6Z`���e	�+#\�-��bO�G��ȱY
E��u���o��}Ұ�u����)m!�̌�27ǭw�^��_�Wݶ���X+��6b����ńlO����4H)o�Ɩ	�*\�ŉиZ3��ud:u��g��U��ܢ|,Y���Z�e!--�R�BTV�@�ȈrP-I��-�$�%m���!6���Н5��J��*י1hT+!Ds˚~��� �4�j�����#uX��"��d�t��3�����0�-��Z��T�Ӆ@*�95-��{t�謋���wS����W�S�����	.���1�  9��}�9��gZI-����]�V4�+���lD��;μ�ۼ���wi$��$�J��I.�I.�I%RI$�I$�U$�IT�I%RI$�rI$�rI$��R��)@6i����pH��6M��Y�UO-���G��M\��mf1�c7H���%���̀�!CE4B�,]��R�S�&���J(�Q	D!D���(�+q�Ӧ��b��m4�����m��[����z�0媼j;֫O{+�o/Y��}�^_7�ٍ��fFam-�R�a}���_��r�4�q�� z���9F7uCo3W]���u:����@�-�k{���%|,Ձ,�����YI*hEj�K����}��M�E��|��Ӓo;��ހ	$��W6b��{�L��~���'!�{��۲�5B���m�fnf�*�D^�Riǵ�>�i�&�?�]���_������
m�-v�6��1et٤)��Of���>=^Ny�{�_]��n�d����e-�YKe����5��{^o�� ���R�f|FJ�j�w���:�+���p��t4��Ӡ�7��'�V[,�����YKS���-r���[��W5|^�ڳ$^�6͙�Ks�v�c  �G�꩚���n��:���<��+y����Xez��O��A '4b!�������U��<��>y��/�|�G�τ����K�vA$�=i��T���h1�t��|����ū����Ѓ�Ye-�R�[,����)l����bo�Z���}�I77�s0���Jm���u���U\�1e���m�m����	/�BI�0�@6   �;�ߞs�x����Di(��Bㆅ�1� Ɲ��m��x�J��������wy��;�۞h���. � � � � � ��9ppvׁ�m��wxw�����8�-��������m��,�|O�	Q�X�������=��_�{�w��@����AJT�7�Zd�q�gk{�'� �zwUm����/�����������j�
֋T=¢#�6o}� ���e�� t��g���5|[�e%$1�#�Kipu�&����YH#��%��b\����K8�1s�d��,ڄs� g�ɋ�nCHV��D-��$�6�8�7��,�� � �(6�E��n�����1/�N�g��)l���[,���YKe��Rٵ�k�1���f/����r�&n<BQ$%W����&��"�CH����~�.����o7m��	 s�LD^��kX1����_4LK6�#-��$�T��Y�Ibo#I~k6���-����YKi	A*��MZJ0��E	D���b'Ä9�6�9�7��m�����9�6�m����D��� m��c�g<1b ��bYƱ-<�k�XUV��,!H�B��!(�S�r�F�n�2=ҽFN�2=  1���S3�����%��u�^�y�\Y�o&�Ml ��u��om�ݯ;Sw�f��ikT^y٥���/|��}!��X��23!��k�ק��|�  �U$��&ff���[�BBD^�%*'t�]�2	$��5�=��G�i���-b3!wy�/���J��I���gsY��eF¶�y�ܻ�@IJf( P�A��s�<�ȵ�ōJ�Yz�4�@6]x!̰`���9�4h�斫�g�Cl&�6�y�z���)Q6 ��CS0�$hS.\�"���i�LQ�0m�;s�dH�v{��a�"�wm�]��nmx�.��&�Iw$�I*�I$�I$��$�J�'��^���$�K�$�K�$�IT�I%RI$�I!JR�R��)Jw�I,�ŉw����
�A3"}:n@  �(�'P3.L̽tg ����K����_��{>3�ِ���3#4̉e���� ��6�6ڏ5u8U�����D횠�[v  !H���o7���O=d-b�'��ԛhI0%5J"�{�a�?;�^����kK\"�� 5u�Cm�F���/f�<ſ1U�EB;��P��h.�@$� ׮��fb��Yub���L_�+�}��l` $�p�|��Ff.��Փ������w�p�u^�~Y�kf�F[l���,#23L��3|y���|�_0G�ih�7����ɧ[�9u5'��hni�b@@%o��BTUB�����<��,�������GCdFn�n`0���bt� 	ҚB<�������Ws���Ⱦ���ͽ;�n� kJ�9���Zf�CX�S_��}�W�wz��R zO-Zn����^�����/uD ���E�)be��3#4̌��3 �J;�t�@	݋*`Lȕ�Ni�#�Oz���虜��}q� 4�FO%{�� ��m�o5��7��c]��"0��W ��c�H�t�,DD�S)CƦ�r�-��i���p\�����ˀr�����뽛<:�D�)
�i��<"v�J�VBX�I,�3�$��p夤%�%�����-�uMl�5w�6�V_#tm�K
�k� #�E	�1M� N7Mp&bCqY��{c+0lsr���!!������j�4�{m�NM�EL ��ȏ1�s�ﮈ-AG�Mz� �T�P�fTL	غ����Q(�b�O�o����֒3#4̌�0�YKe�S���w� �+oM�h$����7�,.�l<�m�Tl�����}���3�3���������Ѣ�jҍƆ+���)�Ŕ���W��s�E�?:I <OT�zCp!ǼQ�k��o�p�H<�"�T�I!ʡQs0�Nh��!{�Zt���{�m����.x` q<(Ҙ�"gĤfeBXnT���s�������;����od���̌�23L����=8�����i_.�رn�����3x�/3��y��xRb  ������s�wյ�ZŬM�טx��S3$U
�C6:x"�嚫�]�ʋa���#� �`C�����K�+kt/ty瑍f��܊dU � p�%&tM+���&����m�iz��b�l/ܿy��TD!$BJ;�S�O��k�NV�P�YE�FU�qi$�I$�U$�IT�Iܴ�Iw$�I*�I$�I$���I%RI$�I$�U$�Iw%ؒJ�/ooo>7���琼��ꁭ�
�<��/�m�j���I =�rݦ�{e�޸UK	����'{���oO��t����3#22YKe��`�c�^kߘI$����12f>V����^w]�u����y^5���''6\��۠[HKKi	i	)��ř�,�M���/-H����>�����_�� ��lL,-�˫��ɵiD\%����2=:�/ug{���<�[�M6���tfwx����o��y���u��=��^N�  7l� @��R��jB��s�SZ��uuVV�Ė��S%����df���̍���=��qNe��1���jyw>�H����g��Ͻb�P�.`�����	��@y�8s|IIXJBZBZ[,����W�Mi��1s�#��Rr�s6\��ż�	$�7eRJf*b�I���ٯ���P��|s�}ޔ���5B�w@I%�i��F�[���=�W|��(�J1�7�gs@�x�y6�"e&R���_�yb>���������y����O5#2n�23V���Z�;�'5�/���鳻Ѷ�hUv�s�ֽ
�u�ٕ�1,�%	D��3�c<���~��%���Gܑ��c  	!��("�V�>�TD;���6 DB1O��E�T[�qW��m��;U�,����d"Q
�D(!Dj?t�X%��� ���E`� ň	�! ��RU�X#H$����5P� B�� S}EJ :KB�IF#����搼 
���PPT3ik-����(/Ie@�D� [:gR���c0�0△O༭@ z`�"$ ���±n3����r��+����E>��Q�D9������1��KB�S�q����g ��]�H)K�  GO���(�ݭ���!�DC{^�_b�l��AO�?�?s[��/� @�2w"!����6�B;̀�X!�g{rƜ�)�PnDB�����`�`�DӇ� i���(��⟴t٧�׮�ߌ�?���������E�� �(���d
����������v�\�|��ԅ���������<+��q3��D��"D�!"!�Р�$臓��\OD7��
=,���	���l[{�- m{��6I�uh��䑏��~�Ģ�y�C��h:c�L�^��)���������I綝*�Y�Qږ����n��=1�A͊��b�@HA�$HA �"Bб���BR
�!�)$K|T"�T`��E�"�X�� (��)�Z���#��0zq���Y�o7��_7�` z;O���(UbDT��	� i�����ݥt4u�`������/��<��t�szL����Fm���z�_�M{�9�מK�"�������� e��~#��Ͱw�_�ƥ��{w���x������#a����}���'��_C�O��ϵ�0���$��t>��������.yz�w�x���aQ:� DR����'w��Y>�Lh|�:���4xk,n���HgV;���h"�S�PE�h��������=���B�O���#FB o=�	�8P*(���G��b������N���豓�R�����d���m�4��wiut&h�v5��$a:"*EZ�!DA��;���r�p�m/�
Bڍ6��Nft
R�=p��>� ��U��A�׏Mw�{7 Y�?a�E��u�����܏�����Ϭ	@n5H�����՞�����@}�'x}3�� �yW�n:�O����a��)�|�����CL7ht�`�(���{|Sc�9?)ҮA	�,0���� z"�A�\2嗱���yG���̓���ըvr�{y�#�����tR>����|��(�j�HA��z���Q���WxV���}[����<-��_�����MDD��i�Ĝ�i!��0)x��H�ö�����k)ז��n7F Ȩ)�-!;��mn����r=�������:u��� �(�{��������J �3�|�_���8�@A:��w:Ǟ��܏��Km~��5��kTp>����b���P����@�>�NG���"�(HQ� 