BZh91AY&SY@�+�  �߀Py���������`^���� |4xx|u� �ݲ�PP�@ P   �q����@)@��(4��R�h�0�	��M�h5<�% ��@ &�h  SƪFD�mM      4 �Q@       )&Pz4J{T�FS�4�M�����5=j� @�<�i�蘚i#� т4@� E��V@
�TQ[Q�v��,+��Y���Ȃ��`T풷�$��L��$G�zX܁"��C�|��^�������ߗ����~&hZˢҐ�����DD�e����h��f̺�%����bR.�(gH����v3�Vi[��*�h�!hZS{L�h�Zl�JM""#Vhf�6��&�pͰ��ZC�9C�����,�-�VE�5rq�m�qƀ�QmA�`0��/~EUb4���W��T]���:��l5�e���{�2�U���;�;]S����wg""�B3M.]�/j&��bV����zq2��<�I�Q���ej[S5�ٚ����8�.�����phywx"�h��^�b��	�L�2{�p�5����fp�7�x$��I�K�T�f����c�X�SY#�t��/ub�gu�+Ȕ�,5PR�S�V���W2���i�t]�ff%�f-�c-�ե�XWQF�r����;�윻�\!���*�����k�q�������#m�F*9������N�*b\��n�
�5l�,Q�[*!~ޚ�_�wbF�y�8�\[�4�h�PC����M�p�߲��')G"5�h��㬵�~.<;n�F�D�ƈ�-������"�![U��A�du�G%�Jʀ�buZ��B����'U�X5$�b�,Ljҧ%d"�J�3u��{um϶���89'/�3ٷ` �<��T/��5�ڥə>�D�򹷧߾�S ��i�y�v-@ z�1�c�  `cm��m���� 5 �.��5V��3	�u =��Ѐ�����s,3�����
.M��d51oD��ч&($C@"�|�ԙݼ�(��n�r�%��ig�P�20�ŎZ�
�
�kZ3��Z2�x�����'��Q��Xy7T���b���Y��A@YAA`,�b�$��c�Z�u���YQP��_9�B��{�}o\���V�eP�UJ��b�#D��-Z��2ժ&�B�F�L���</�T��ۻ�fj�'�"ϟ��.�K6�����X�K%�lg��9�?2�P����J�a���_T�V>*�b��얳�n�����;Sz�$�s0.�����yvy-hH�3�D;9[*,>��t��v�/r���M9�b0ŵ���̨����
�/"�<�4���6m�T�b�I��ڛo}��vH��v�*��+�|>�=�m�d����<�6~\�����>��}��]_oϙ���0�����6A���qQ�5�������ǩ�ⷭ�Խ��p�dƬ����y���w0��X{]h��L�0�Qi/5���껼3��R���s��x>��:B6���΄��aPP&r�V<==��e0��M�y����*�
�f��+i��|%����>�^D�W|��[�Vnpͼ��n�svQn�����o��E�e���T>�>HI�C��lxzE0v��'���ʶ�bQ�t�g�6ޓܜR�xD������"^�e��pI!��	�(s��N8JK(��R�))R��hє�d�p��Tb"���aoe�fo^��_-��E�y�hf�QJ���X��M<n��#�*� 
���Ri	��4xhd�Qj���:�f���up�=f���c]x{�L<H�B{۸Cu0�o��⡤+��n��&.h���/\����u�!1�<]�i��)
C\jɃ��/44��w�M���.���y�$� l�6N.�*�x�9�f5 珃��i���:�":�������Ba~ �#�;U�*!�yB�pސ.!��#��/M$#U��`r�HvU��+5S��a�Mb�$��l�'�h�.E�6Z�~тZ�ar��������E�����ݺ�[l��!Tˢ��)5�*Td��R�����{>!���Ă[�W���Ƣ�8B�l՞ȼ��L����Ra�y��,*3���;o;Z����	>D�ȿx�&�{�ֹ�#}�/u��(KQaL��ڀ����� ��rf�^���w�\<�6I��r�rF]r�p*5���SG�6�gR�U�A�SS����S��t{գ8�B����ŗ��MJ��:W�bG_?�=��e�FC�K�8c�u���cY���u��Wq��j�	J�c&R�cɄM�ev+E+u�Qkw|Ǧ��Ǫ�f����e�&z��xzHcAY���]\�!m����w�M��sp��#��"S��u\{�#�.�ˠ��������CsvSʖ��I�o�8�=T:�vo���C��mя�gEU �ɽ��o(W�d`u�AS<��9L�
ٚ]���9otz�tD����3a��f35c�H�'���� *f�s�dP���"A��n�Ęfm������G�x?���U������$�M�j�?d����npp�L+�̨��l��J|�M?�����a3|�ӽ����f �Xw�c�{�E�*DQ�{n����w�`"���:$.���gJ*�5::ٺ���Gp�p8��-��.waD;��C�ضq��VE�,Hr"/b��S�ފ	���"B���ϴ�XƼ��%���-	D�ɱ��+b��JI3\�A:��'�����g��<��h�X��4w�R���*�抔�%uUP��tY� 3�t賠��.n�+��4�h����L�;E�[67�Χ�P���1���æ:�<���0�6��n�O��V���M�h���ds��8�E�0SI�=�b���f�a�d:^%�b�Ǚˤឲ�Ը�Xx�t�NDoh/R<Ǧr{q�g��b���j���g�e��oAt���8�9z�ܵV���ښ�^=�5�d6*�d<'rї8m[���L�e��>e�o4U�B�+J%X�he�%Ck�\�C�&�|��7������_�EK|�3�;��3J�#�(8�z�w{����8�L���<���h���1�f�3�<k>�#+�4(���J�Y��}���׮p�zl��v�-��2���v�zuW�9�T��Y!�xy�W�3[����BOj][҈@L�qx�.UQ���)�;���&*����L���d�س��ܭ��7�wx����.�Z��k��x���'d"ܗ���>���1��U�k6�/��x���t��5�ע�?��k�����|�]N�oυǽ#�(l&��`<�Z@�c2���,)k<�����_t!�Akw*Q�l@���̞mh�ďy� �kfc�H�7ny���{��|�����پk��U,�wk���d;�l�|�1�ѳ��B�7s3��0|��O%0�q(��k��͆�eJ��Z�(�.��=�� ����S�k�:&gdQs��n�y^W�A�-�i⯅���|��ړH?���Mõz�[���r1�U(��v�fj��&�V��?oh������b�T/�2e�lB!j�����w� �!�|A���$�Ib�,��_OP,wǢ$'��@PA]2+e
����$Z��[�WE�����!7P,a�L�b�����U
�Jp@iQETUEP_���*ґ[��aB�b�#DD��P������(���dFE����"1�EQA""#��,QQ���b"(�1E"��(�*�%R1EQb���4F�EQH
���X��Ң�*�X��)Q)
ŋ	L��"! P9���
`P��+%��[a�9b��p%��3`LY�L& L%	h���p�!����cKL\�����"�HE'(p�Yݦ��t��gQu���������uϮ�I�\�h�u��&�9,���93�ń����,����pT�����i)x��'Z{���x�^T���|��� ���_�Ȃ��<4L�{�&�P���2D�4{�{�����y��6(���)˻j .Ѥ��:zhA����L0JII<��!&��5l"�T.���.�fY�>o�g�r���@`���/��`":�ѡ9 �#����O:\{{S�_D�>2�̢�@V�dd��E
�(�"�`,��"""ER(��,DF*�(,�E1�"���#n�
��A@DUX1DEU���+@X�+����DF"�UQ`����Jd@��P�3��Dދ���]3�ړ�C������m4(4F�d)����(@�e��z>�|X��4;J���Ht&�c�ͤ�.$��~��4�N���c���f950(OB�
<�鿡���{�� �C��rt�/j~���KE8����l-K�ʛ���0�p�M�r|5���?\MC� .��{""45�?�`ϳqnFY~��;��M���B�$���Q��
��d<L��!���`;S�w#}X�B({#�Т8q#FX� ����Ex�Ϻ��!�۷0����4��Y�h����8(`�@A��6th��8�K̟V8����Ai0! ����'>C� /��QC��į*3�?�����'�?eX��� 0P�5��^<{���6`�ȣ���z:���.�b>`@�y|��v�D *d>b�Dl=��Z7k�p9>����� m=��"��H����PŒ̫mN��!��3���6g`3�=pp�;�&�����n�;LQrc�A�pq%ڪc���)B\��q'���˺/���F�/���*P�+���� p��7�bQ��ճ�q2(hF�ycc�B�Dq�iPFo.�g�dǄ�c��p�@��^�Hz5���mWO�]��BAh�p