BZh91AY&SY�c}$ �_�Px��g������P��#�b63	$ C��ڣ�z�'�4�@�3P4�b&"�     h 	����1l��C@  d�4d���`F�b0L�`�$�`�y��=L�I��� �2=Ae ��@@ ��O��P�� 2}���"E���8��E�&��X�2�����d@m��PW4L��,��#�<(��ެ�gɄ���UuȘ���-�S`����'�h3�y�`I��a}S%t5uY�_L.��^���c}�@�n�hf���#��-���Xr�O)�)���q)�uP(H��i�V��C:�eI��ČcPh��L#����J�)LP��F�!U!��yr&JJ���JX����Y�_D�K8T�uK�.!eV�����j*h&��(Hm�m��`8���y���հ����j�X���&z�0� i�1�TB"fI�Pu2�]B
a����#3Y2���ųu�K�l���C|���r�[�w�kw}���V1%$���@�ɴ�ˆ^�C���gձd6���x��V�p��@�v���oO�.�?�u����W�b�B��:��y��!�;�o%yZ�N�������7���];hT;�5����-hd~���c�����3Pѩ���
��y6��\3���v6�D�:E%��U�C�*	�ىIS��t�ྫ�O[���L��a����K�]n��>D�e|��vR�I~讋�~e}��2��,���6���	j����ߙ��25�"�0=�2��q[8`h��j
�i$Y�
�46�\�v�,����c�	���IAE�Υ�)���P��aJ��LêWT�f��p*6��uP����t� ��]ebN`<��>:Xn}��6�9�Wf��E�t�G��Q�y�X&ak����(=�WiM��o�Y�Bj�m�!3f�D!ְ�M�����;�.�]�s��J��:� )+nMƻU��2�6�U:OEL-��$	�5Z�����5<̆A�M���EP�-L��ZhA�H�FW�{��Kh���jeg�\6n�,��T����H�
�o��