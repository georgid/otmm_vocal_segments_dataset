BZh91AY&SY���� Z߀Px���������`=� �r�� @  �  6 O�����	����ԙ i� z�   d)HQ���#4��@ hhɉ�	���0 �`�0�&�DԠ � h  4�i2bz��2b�dA� �D0�A�4�=!��yLF����OS�z�PP��)�H*� ϯ̧���	$DS�DB@�?�M��?sHHI�HNXOq
 �$Lih�K���5��K����R�G%ʈ���w�ss�Xp�ËaØ�gÏ��Æ�f&�XF�ai8F#�'1�p�m�$�[Zt�m$�$�r'3��u3.�"L6�m����t�:i�Ø��f88��pm�D���Bqo���<C�>��I_ �G�2��7n�MV�����V�bzy�/I��T����b��Sb����Ш�ņ�+��&N:�N�|�(���g�D�%ѓ��)�[�p^g�;BuTw2 �uj�K�Vn�0y�*',0Q������N*_#K��U���T��%�g0�]q�pf�˶W.-�Mib*ܦ��۸������ۃ1.TknLԭ�73\ͣs&;ͻ�.������	8v���
!�v��w�c30+^����H�B����|xeL�/E�r�f���nd�Y��fff�[�K�خ9,wni�˻��-u\\ڦm�V��%���׷-�6�<��8�_jۊ	1v���13γ��b�kN.!l��6�m��    �c    9�0 � ��m�  c�      I$�  L֍��L����+"f�l�CwT>�ȃ6�0�t���qSH�T���
�}w���[�������'V#$h
�W��JԱk�:�?]f:�" �[��ڜ��?]��`

�n%�	c���T_})���Bq��:|��DJ׫T�;��������jE�r�����g�wy�.+�L�[�Pap�{,=����O����(�7��DIm�,'�.B.$��9�B3�=���f��%$!��rV�u�Zs��(�H�J3�?t�m�F
7*E��1�C�`���D ;50��/��4(��0�e|y�[|O�J$S7�-`���U��ߞwy�|zΗc���_@ ��f8��<�Ũ�;H:�P6J��l#�Y�F!����{���M�FHӞ��d��E��Q뉭�9�`[��"\�ިiiި��&Y͞��V��������.��зh�%���1�e�9�&$����C	!��.݆�#.� ��j@�"��ia�0��3;�M'�y��u�#'V�0��8�8���4A�52\n��/�ݜ���Gc���$8,�H#��J�çFBx�5�xeI�q�fl:�ԇ9K����Y�;%� �:�q��v.Í�Yg-z�ψ������'�~���B/��i���R�,&�����YgLM$���k�ǈ� ���o=�����tZ�DXAu���G��c��f�����S#���B��;���찧�w�͍s�G⛅����b;��k���ٛ���w���Bzf�v�v���9He�,f�ʟEl�A���{T@vv�B��o�%�۹�}v.�2��<�Z��Q؅��;�3���<與�,�ݙa�	�VD^��RTf�Pμla/��\���՗�D����ͽ-���d!9�=����zS�
^�|�5�00��C2%&�:JrR	<;�u��*������ƿJ��@j��>�GyX�\ &c���vt������_P�����<��٬��U�Ë37<���0	��y���4���Gz2 ˿P�X[|���oVO��~|��W����"��{��40?����`7$	%v��;����zK��?
��F���}$V�e��$�"��c�
S��-kս}���Fz܍�n�����!Zmd���=�����:�V]��M��eZ�x��Љ���W����oo]�T2A(:���tc�(�i;�{=��'�����`0�1p�T��+�a�N,��8�ܦc���f�k����t����1S6�o�s&)؜q���.���ު#����L\l,�D|j9co���FT������G��'��[[����i�K⛸��¦��]��;�F_��3���Չ�ͯ6���*ɣ.r�5q�b\�p�w�T��f �B����<�>�6��$]fɋ���j����)s��CL8�D�h}�Q���޴�l��mǉ;f#	��h]<��̑�>tN�ǭL��	�6���S���Sw���Z���1<μ,b�ӷكD�剼I����|=�[zLy=O����l��=��ɇ���3�H ��I8\�����ɹ���!� T ������k=�DB�RQo�uل��D��78���PS��@c�0N)��k�>y�5D/G5����?�����p=j�0���/�b��_^�7���,�rs�n�H�؄E�����6�ݓ��1,����z�î���B����&a�\%w�b24Eunvo;��Ժ
��[�NY�X��E)��RA�익��CLC�'�|}|c״�nȧ��_G�����َ�ԟή=劥�g�?z�)�y87--��=�+���lu]57y�uqo��~OvG��J~�z�Fp�X�$�d�$�I$X�!E�O�X�� ����p��a�;�<���<�ͦ�Ls�&r*��`������*(�h��R�"@� ��g�ɀ��k9�Y�������b���QQ��R��*�Q2�DETP�`��(,X�"*�̖I2@s��jH#$ �nqF�13� ��*��CYQTS)F�u���-**�e�QUr� Q)�KUT��t�UTDY�{ z�\p��D�
��}��v�AY�Fbb�b
�m�{Ek�����go�wo��{��������t�Gy,�u�=3:}86��ZF�%�.v�_��d7�nW����1����	�&�r�M>��}���B����A�4v�K�Ө��r�ؑ�iP���"�]}��C��;�3�*��J �d�4%*��<r� ��C}IjZ|"<��/]�%� H�����ǚ!�++�.��L2kS�Y�LE�%7=׹h�'����&?t�=����Um	�d��AA�#�EDQ�����"#QF"(�#�R"�*
�����h�b$V1R@Y	��D#�q��\��������`�1é'���q��F�@
r@A J����E #
! �|�̼:��4�g"��>`�t5s�e&Iq,9 ��20��$��qG��#���I�^5wWC!��y��'_cbs�/��X�/����|��I���\�Md�Y�=�+[�4u�16�D4�QE

���=E�de�wbA��gTE�آ!����03�by��^4`:C�@(_cI��Yp�
�F����F�X�X���<8��W�i�z��T�P��8 `Igi��l���^d�1�-d�?�Њ!F L��T#n��QɄ��m�d�q%�us�Q��h��JA�YI��O$�l����X�2�C̣�C��v�����H�80�#�a&3i��.Wk�l$�V#״qd`<8���(��%�V��{�ɉӯ�~�4�`3�=�8}��&��hh�u���UBO#[�5(K88��^����3s`���b��+��;sdg�!�`�"��m�3"<P�ppw:L�P�d䂅���?N�S�%�n9�=����C����܃5Zu��.�p�!{u��