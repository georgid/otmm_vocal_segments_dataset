BZh91AY&SY�0�� �_�Py���������`|� �<�     (  �)�iP��em@	"&���*mO'�~���3H�44i��i����P�Ѡ���  q�&LF& L�&@F ���Pz��   �  �	OSM��P6��4hh�@D�)��hi='�=��jC�4F�h�p�%�p��E@ EL�{�DЍ���Z��R 4 �A�~��Xcd^L�����	:qTˇYsc�Wlޣ���6�O*ݪ~
��t�Ӻ���N����t��CI;�iӧN��N�����HԴ�#H�4��}��ܭt����ݷ��iӧN��4���we�;���������7wkvƝդn�:B-����N���sPZ����n�'V�:F��Cu4�-���7wFg3fx9��ߝWϾ�N@�+��Ϸ�В�A��_i��F�E1��*dڄ*��ƥWSp�(X���]'�"��MK:�̅SO&؇�P�Yϋ�%� �;�L*~P�����+O:�VB}{ڥ��#1
��hlV��*a�V(J�=M\�,��URҤ�P|�E���J/�e��.k%A��5�oWr�Xdi��I4��0L�hkMl�T���%��UD�T�9c	[�B����2��v
I��6��[&Éw1��=E%C�_m��5�����eP$-�ZK���ܳ7e�<� �@9����GŒ��cv'�%bj
�(��,�c*��V��b��=d�}�yRB	#{�����  
ަ4RR(̰؍
��zhQP��L�v�����rOFE!�����8�7N�؏ϙ��0�{Kv��2�Akez7f���1�8�5&B���	:x%��Ͷ����Y��Z�)\�#"�G6˯�紗tm��b�0Y�6�rSO5��j��ޤ���LE9�w���oIι.m�oE�|�z$��?��n~��k�!��U7���׭�B�^T�<B�c���BAfn���݂4P3�=��I��	���	�q�E��rR}eKH���囡 �GdJ��������|�4H�q��%��B�n-�@E�]Hܑx���"\�$H�3���k@h�j벡ρ���aaK2���u0��'r���>Kx��>"�X�;aFNU�C�N5��7d;0��ZHӿq�#'^}��DyđD|G���ߘ�*�D>��F�,Ni��t�6na��	t��3aj3��E�k`�ә�+u{ɀg
�R�{۷!o����1��X��)���L�
AEܙr`�t(�*��ՂEd0p�Đ�(����ŋSeD��ޑv; G�bvr4����fi\X=��Dx�ZL�Cy��G���I!���!�]s���y�2	gp2 �,��%����+�~/��� 	G��K�A�/fN R�fo	���ld�lm(	Xsw�0�v,���aw,t�¡)G�瘞�߳�4r�~�;Qw�/ɮf����jHz�ǉ����F!��@�y|\����&�`9ώ�9$�;X���=Jd���8����m�A����N�!��8�6�]�z+F�u�1�T%ߵ�Sg��_J�.�t130�$?�<��}�H%�5@�R(�ȉ QP\<�;�/���`�CT2��F��]�9O^vD�8���i0v�a�b�;�6l܋���i�������&#���x�4�?���n��q�J��'���ZQ��G����['�/8%3y �y�H��2Ð0p]���!ŋ���w=t���ĉ����9讧�>}7S3�5ݹsʹJU�����}���Վqn���B��û���T���հ��zħ��$6ҡ��焻��rL�b�<l�RF7DY国]Oz�u9^�^,42��t^h��oY��Ȥ���/ٷSP�Jn��:��� �|�솿xE�]�(�����i��E"i�Ƹ�bYl[v��v��6��P��#�T�E����}7�u/!��謨.�t�����	��/�fj+�aZ�⡏h}a5�}��zG�6�.�pUm�#x��b�� ,�L� �#�"�\(�vfw%���[��.�Rx�06�g3�zٛZO��o\��]�)d�E�yPޥA�p���^w���G��z�*�y8:J�}�9��u����Ε��n���F�%zy@�,=a���D�M�4�a��L}��. ��;g�:�����X�.�
�1���wi�A%-e�B"�K��Ex9^�N�;cHQo�S!�>(U�ᯖq@���T��C�n�'R��
;ݵ��T֮�+l���@�����r��`�d`��YRr�^-��6*!ͫ0'��mO����Vp����_>!.~bK��)�����&�+��.�*�{�i�3���|f���
���=qF�8�7v�ְ^�^�U�$�N�Cמk]����N���x��Z��`���d,��+�������A��}�b�������0������6+�!��,��>W������&9Æζ�cwV�72SZV��W[�p� �bQ�ā(�S����eeI�	' �L��vT���v$b ��w�S}��r��Z��S{yY%+R�
#E,�hP.�PR�(BSF�4e#�S�q�N��Cy9�7၉���@�ңJ� 3"�ܶ6m϶�sS�|���E|�������r��Qm4�EF���v�*UlJ�Q7�gT5����|�κ�H@�ie�+�#��t�h�T>�9"��w�AؔFB��h������D���3��>`�q! �{�����X�� ���9k>-o~��V|7!�:V�Q���k��:�b����=~*|�t��n�l9�~\�
 t�P�c�[�X+�_7���0�M3�mB�Z�@���B��B���i32�$�c"T�Z��b��j��
�b"�Jf�@�}q��r�1��P�
�u�:��r�����Q9�P
�T���H�(R�(R RW�ba�����q6���G�!�h�du��� �`]�53�����u���c��(�L
���)�x_�>���؝��Ҏ g���[�|$�"��IA�L{�$�)�*j|�n��̎�L�@y�
ё����8�^[q1���{�b̃^�
���D�;�J0��y���h\9ô4*mLL��WYQ;R"�b�MrB��5�#���*
P�Pl6�t���9i�&Ә����t���g�s�.ӹ�ry3��J��DJ�3j�p�	6�;;;�+��}3���B��>��<}������zu^Sv�.WߖI����Q�C/YĮWd)��"C���1�q����e,z�8�]�g79h��8�=�I3*1����(Ԭ��FR�#u"`�������Fk�H�����L^a�GAp�%�|ؚ�M���)#���5(%uJ;x�8k��,�Q1b
�K���K��3����`Ȯ����|h�|�w9u�$W�D���c��uNp*[�>���2'9�ߌ1��4�C�OMU�x�����ܑN$0�*k 