BZh91AY&SY� &߀Px���������`�}n
>��{����D�(ҁ�l}�Ư�@�с�CA�zf�����6�F���D�T0 �0  b0�5T��0 4�0 12 ��SH%4m`�LF 4F�J)��F�a4є��244h���$!	��h�=OSjz��L#A�4CM��'!DJAAp
	�*� ���G�"H �������I%�\QWF��D	@Ճ(��uӷ�~�ݐ��kծ���(ʒ��YQ�BN	�B!B(�)8D"�D"�E:�Y�Y�:):,�D(p�D"qd"�N Y�HB(�E�"�E'D"���(�Y���C:�Io㩄uݖ�P��:�p�ꕤ�8N�j3"q����͊���UHNUBv�g�G�|(/r�+PqS/q5V]�j��vN"��d8�w6U�DޙxIf%���d�k��2�Sv�B�Z��^���S���K��6_r+�d��q�;^%�a<
9["U>�;9�iF�d�e�̔��;&Qб5dR�`��B:*��*U�d��B��5H��Yce,�t�@����pqڭ1Z1U �$v�^̙^F�M���KKڀ��`��x��T���Mf$$��=Sf������r�.�C˩�+n(��6,$B�*qۈ�E�exdE+�!��q���R�b�$e��������g��yq��ԒK�G���\�Dv��kq@�n��D��d���ާ\Pł�<)o�^.��n�P�w�7����jn�b�	��w7z�ʛ��{De�30ֶ��n/[�{��c"��#��G�H ��@�[��ܝ9J�V�Nj�<��	j�8�"@��z!	�j��e��.\s%��e
��W���)��[R@|vPآ���)���m�g\�x{FrF�&4�3{])��'0��#d��K�(�0t�yͼ�`:݃��;:���mlei͎~�n�w��˚���v��w��F��\�����GT/�f@�^5�}�@f��Z���p�dk��K� g4y.Ӱ &�� :D#��emt���.t�}�A벉���W�pnT��C��(�jG��P�N9j������׎���� Q�$�O���f(O�d��;�כpH����=2`h�0����"�^��v8R�L�b
8Ds��Ǻ�6�=�p��f�-���@��e�fj;��CU�m�����p4i�hH:o1.T����"b��ˍܗ9�V���\v�bN[P�m���/@���<�s���{� �³��ą@��G����ݘ8I�I6+)*.�"��Zs�C�tN��W�CLTq������"Hb@qN�t�"�#|��4/�<������I��t������p�@#�z��hi[V "�� �uk��r"� ����R�[+4�]ѕrrG,#A����q�Ss���&�mǅeu �[�n&��G��^B��nx��8c�=C	ʉfa��>�*��^x�Û��'�dL�w�Kc3��×����u^�H����'DV�+��/�7-�f �����OKet� �&��_��2%���&��XQrCM._�if,�\-1�� ^%̼9~�"��q���N�����$�vf�1nJ g\NƯWU���}cjf-l�4��0���¤���AA�y����@q�܇��6#O���H��3�%@��z�!�@U���My�N��y2	`=P�ܼ���幦'=��h�|���0ի��F�0 [SkK�P��i�+1Z��W7��G`|~�ϦՃә�c��TLM
9Ϳ J�@��ظx�b�}��DVp����2���Dׅ����S��Q�w��Am三��^� �A����kx��'9D]`G�c����n�b�R�2�A��X�(-@���zn2�*r��*@���;���)���n˷-Y�2�u@�soZLF��{��V�T�?>35�����:�kǮ����_ه\���cY������n#D�{�En��q_��u^U=��p�����K���&��g*�*!i����� �p��|�f 𮌩1���L]p�E�y��/?a�"]��ç�W>|n{��U��H�#���}���t��S?�E���|���B��������n��>2T���b��<&s9c�VϮ��!u���-��W*�ձp��&'�/���%��IE� � �Q���S5��&0�����D�.ͤQ�,��`p�٥K�(���m9V�J;@izt�fq�|�f3=0�Q���N֯���;ޭN���:!�����T��^��Ϸ���y`wL^�C�C$g�+f��(h�`��)d��u���Ċu����"��\��q^eQ�~��QG<"�;�N��������>��|��.4�fh���/B���g�.J0ek���.Ƭ(*����F�z�`�@y�_H�j�X��b���*�g��3�4��L3R��-���~$Z�����ͣ?P�)HFLrI$�E��(q*)�V���� �O�/m,b����2n�*��e�⋘m-�FE�fp�X�BP$A���� ���\KŊ�DT�H�Z X"-Ֆбh�\�����A@$,iHZ%�HK�l[
*�*��b�+�$����|�ظ��&2��;#ܛ������$$@��:+w�~�6�7#�y?W���������	�.��G���Ϩ���P�)��9����B�<��w� �A�����H���b<�*^@P�<$ ���tJ�||����:R4��
w������˲J���铯�DB�@5e)��B��OrF�Z{"= S��=��|p&D��-EGIYm����W����l��vꢙΌ����h�'m�//�:?4�<p�J#
� �V�@EZF��(Z�E(EB����D�DTQV�Q��ZAAE�AS� �����*�"��Т4)T*� ��UU+��4���q�g���5�:���jpʊl)�v)AB�P��Ȭ�Ȭ ��Ŧؘ֜��|�m�X<�����]
L��XsSߙ�/擝����q�`@Q
zJO��j�7#1�p���N�[��_'��ܾj�Q��:����\�˟ ÷d�ݦI{~�S	��! �*P(k����b��y��c�Ԑf�׍(*��Q�u��`ga��C�xс���K���dDxG|AR�¸��i%�0��v@ ����o8]\CL4�]������� 4��6�h���^f���-Y�~�b(��-pp�o(M�c�DC����o��,ª�`>^�N.}��dxκT��V4�FRg0��h��cV(s8����\E�dO:Fɨs��c[�����xw�7�zR���o�920<\Z(�E���|��Ǡ�����@�K�'@�~�;A��6m���<��QD�����b	b;��|��7v��TS����b�p+��|z2��C��D>5�9F���#�QO����|�ASz��J��;4e�wdJ��������ᬆ��5�(nW
����"�(H�K 