BZh91AY&SYֱ���߀pp����� ����ao�  ΌD�("�H
     
m� �('Xte
l�  K` 
]�                     h  P            4   �   ���}��5ݾں��[�sKqUv���W��`J��ӡ�A�����۽�<�uLl�> �*@��(8�Z�5*`;���H��]���WeJ�:�R�m�R��Sn�R�m�gJ�Y[R�[&ҕYwjT��g[T�]� ���Fl����v����F�^޺'�]�Ut�N꼺�٣=�ݽ5�w�/{V5Wo��^nu܀v�{mw�O   �,�����nf��c�����w��mn��[C7Pn֪�ۘcҽ�޷����a;N��n�u�9x��P���>�ݼol�,z��`;N�)����oz��R�n�I��.[�HfmL��݋����TJ�F;׵j^�n�6��+�Rv�����IFƝ���դV�����l�eXwuҚ�%�R(34��u���]�νڧuJ��էc\�v��,;�q��������uJ��S��x꧉R�(P�Ig=v�+�E�[J�{��m�!v먮��M�suv�-Қ�Uv�M�R��Ӫ�� �7�Ƞtk�B�)S����s����Үێ�궬�7\�7�J�:3ujV^��y��Ӕv��  � (�K<�����J���5|��zS�{�Z���x�h�k���N�ꋵ\Ք�w�9{��5� �       EO� ��R�M F  =C& ����J�Sj`      O�*��ʟ�       S�)�`F`�d�ѐ�L"�*J� �4 d   !H@��14M�I驦�S��Q�((����_���w���y��a�k�}׿�@U���%@W�!x�*� ���?����_���?����/�� ��P UX��UU�
 ��A�d��Ʉ� ��������<�@ʂ�)_�*+�`Q����PZA�d|�E��_ |��G�E$T|��T�G�_ |��G��T|��@�_!� �H� � /�����@� _$|�Q�G�Q�<�C�SR������������ w*�
��� �*y�*y�"Ԣ�P�J�N�Ez�U�AW� ^B"��"/���@��<��G�_%y �
��
>J�� 䪏����/� ��E��D�?����~G����ֺ�5��T��|n��w�⿸�~cQ����6�e��Y��!22�I&B<�{��NN�:G��Bo���3�j�g����R�b���<r�0�2�C�_������,ƴҤ�
�#���4�=q�����e�jx��p��83*T���MBy&�P��ۭ�$)��/q��{az�}sv��O��y�47i��to[7�5$t�4�����F�D&%|NTc�Ȁ���B3��y� 	�
U����VF�f<>H�H^@3�1�y�W��4��:����v��w�&�9	BP��n�JS���gR���g� �����-�#�X���7m���&�A�O6�)A���d�	BP��B��2R��JR%	BV�2�c��%	I������]��'�����ON�5��{z �V��Bj�C�;�&�3@a�x���,ۉ�����u��h�,XB��8��3b �+�`Ύ�j�C�����5C�m2\���rv�@fC��d��)mp�2�t��:ڴf�4:�#�d:��,�2���+l�n`��F�f��t"��BY��}��#��`Pam�υ��X7~��YLO��y���&����Y�/�g��Ha�fB�����<����	Jf`�du��''���g w�{���e������C�L��6H��u&F�PAD�0J����θ>��S;5|Hj�:aY����G�r���3��{�	I����!+�L�be2Kx��)ZbU�!,A�&y}�񖍣EV
�N�+Hdγ�RGOF>�D".�I�	L�X�~2����_*��}n��~�c%�����!4��,4���q�{u�Y�uxg�zh��a���r�ִh�-j�9:�\��R�л8���h��<��Z;KF���}y��Ѵ�A��ֺ�\�;^���p�Wo4n����;ف���
M�m�g��-��s\��3�o9Zx͚ܙ�čZ������\��P���z�|�G���/5���h[�:�h/�0�9�7�9���8s�c�4����GBNto;���#Ƃ�1�YI��	C%)F��X%)J�)��A���&��e J��R�f�(S���	��A���O��2P�0�$3S����5�f�Z5;�,���q<�k3��"�a��9�ym��4=AՔ�˜�c ���t�7��U.4DA���M�-���u8P��`�>��(��k����_-HP����D愰�5Z��@�N����'V�߆��p����c0�y��'���!����@��H���-{��F��rh��������NF!�b�F�9���Q�Z�����d'Y�IR��GT���p�Z�����j�$(J����̻�N>f�4d'��JjD͚ ђ8�@{�	ԇ���)HP��!Brd��/s�ڐ�� �
��(J��ma���I��h��a�u&��1�Z��P�%	����&A�n7h�z�N.@d�ٻR%)HP���bT�C	y�R%)HP��!Jk�SR&Jd�B\b	��rpy%����%	BP�%	BP�'wR	Jd%)��9q�=a5��V����Ý�]uW5^�GXh��2u&�8�	BP��R��)N��{	@x�a��x�n,�i�K�c����tՎ�P�8���i�V�;d��L��r�@G�����c
'��ے�a�����ݷ4&�&��M���M��;���s3�����:w�;h����N���4�q�ߙ�����;��a���q58�,T�Yr5��z�I��8BR��	JjCP�)�bG��M��u2���n����<�T�@�@w�*��r �fP��'(u�d���ӎ�a�O0;�d�y<���ac<�y��@�Ӥ��J r��C���@t�|�@����rz�*l�n����Vuk�c-R�LXN M�yL
���g\�]�]l�5a��[vOD�4T~��S�����F4�&7>f	�e��������@"(T�f�3-�3��1P"XXj$!SY��:-��ٙd�ُ�6�ٓO�"u�ƺ��w��4Ap�ւV��2�j��f��O�����(L�ԅ	�O$(N�)���z;����͙���|bY?}�?��a�G�LQ �`���*�S.υxX�,B]B`k.Xq��,�����0z�#i���G���*c68FX�=�bY)F�i�N��{�n�f��8NHw	BfA�SS�d�η���z��:��|��Prӽ��u���h���F��^'PabA��`����$�f��d0H�B�X		��.����!�i��!���``�"�x�+��N�h�c�c uCA��*�\Ô��G��V�DF��hѣ�Q���h�;�5Fsg7	F���I�3���Q�vf��q�@�@0�&�"<�� �Qo�D$�~e�iy&���Du	��b@q����a���-z�y&�٧P4!�nC$(JR��)i)���5d%/���%.�d �����.��h�� �@1J9Y��(^A܁�#;�7�G�{^Gz׶�ЗΦ5$:�(q*(2k$9�����z;�ރ5�N�Q��.baOv�����kX�b��$$яa�`i�Z�4�OmN�b�-.�K��e� ��yU�`���x�� 1v����� �D��v�Mu@eNM�``d�M3)!l�ʐ�#��S�HAC���}�!��6��̓ʱ%]_�c����P�b�X@C�b`��VC�����7� ,H�����=?�ﳏ}�����~W�#Q6=_J�1�﩯�������"jV�135�3.Ȃ���n����Ra�Bꀎ@ct��V��V��ozg�
d'`dE��C��_#'G�k��ٳ�ȋ�s��k�6dEc������&��r0j�L�	#PfHy!F`�h�Y���Ot8��d%/���!ʽZ 0�5A��̀oo|j��2�d!�ǈ?|&��1��D 6F iyP��f��������L���Gn���3J�#@_ �b�p���#����~c�!��Lwk�Fh�[h�(��?1��O�C��敖����^�M��r0��<c�"j�A��ǆ����=�PQ��U���c	a�c#�oų{�r��@/����@!�p/
�(�3 b�%�^�k�YÅ�9����<�è�o��p.Zv����DvV�1���u8f��B20(�W�a�ʙ �W�ȿ�`����rf�5�ə����t>��������X!aa4B�m߯32XG�L�P�[
��z��hu`t��.F���óxe��TWPdʗ�	iJIvr���
to7	HA�#�M	�`��&���-&�-�d�PoR�X;���B�
��X�QԹ&��N��PaQ��8s��h����<�5����Q�z���4a��|�bulx�:'Z������i�F�
�4w���%dd�!�fF�u��&;0)�0��]HP��!BR��>�<����u�ݏ�x��\�����(JR��=,͝/ptk�s�]�a{r�"c�ĳ5�cp8��lޢ���V����%,L��(<Nk0sV!GO���5�as���µ��H�f�HP��)ip���(J�3��2Mj=�׬
6JRfo2�<Ύ���Ld&������x�Y�,�E�S���%	BP�'r��!Jui�����Hw	J��62��x6>���/%���8vq#�/<��vZͽn�c�sĲ�@rCRj��f-ְx�������e�����V>Y�yz���a�	)	��&O�4� ���/��p�W��]�Q�b|���2M>��1��l�������`r�C��M�6�	������ꐃ�����m�jB�ԧ�%)���i�R��	JRg=�^�u��#}�k�wo^fxgy�˭ϙ�y�P���Q|�14#<���;$��ģ��n�Hl�:M���5�Pc�Plr�#��Ju�ӻ���}��μ��{=h��A���,�&�5�L�H��0�.*�&IBu;\� �B4�C �L�<a�C��R��Z�D�.5'A�17�dL�f�I1Σ�)JB��)�R��<�Ԧ��	��b�����,���P"���u����:L�tǶ��Y��)F.C�[�:wĴkaʋVư4��*��+�p{�F��{����������]�b�7g���<���1�ڵ������?��k�����������aG�}��������{�f�'���������H;%��tttttttttt����GGD޶ب��������A�-����������������w��ttttttcc��T�tw��61�����������������������������::::?ã������[I$������������������ww�������m�������������N�	��;�2��TB�]������׮vz�ӟ�rB7���]LT�����m����m$y���*�����GGGGG�����y.�Ŧ���� ��`�m������nfS^F���T����������:s�|2��e:��:v�$��Ih�7*��n ������������m������Q�(��$H���Ԑ��R�ꚢ��l�#i�GF��$��h2j��L�9�n�%�<�8
�wwIgyD�r��Аz�vBE�ﻉ~������o�W�8��l��'��
���'t�{���#�ttu��qG��s�.���U��K��uK�3~Iܻ�Β�ܔT��I5��߮�NǗ����Gd�p�[���s78xN^H�����}��w��/)1\Ǚ��{yGW�3�����f���π�gL��ttt���'��v�e����zj���c���~����R?�j7�I);��򙑭ٞs�If�7WM��٩j
	GG�Q�����������������������������������Т�RA����������������������:::;%��Ki ��������������zp���������������������(t$�	�������GGGGGGGGGGGGGGGGGGGGGGGGGGGGGd���m$�����������������������������LP�H:::::::::::::::::::;%���Ӥ�������������������:::?��GGI��:��� �::::::::::::::;%��Ki ���ۻ��������������������������[i�=K:�KGGGGGGGGGGGGd��Im$�tttttttttttS�t��룣����`�(�����y����������������n�[Id�����������������������(�:J:::::::::::::::::;%��s$����;m$��{/����'й4A���}eJf�E�����9[u�[��m}���i�Ɨ?V�_O�x��w>�N�����^��������W�vjל�
��n�{��Z��ݵ�H6���^��Аtt]�M�$!���v�����^������b�Xe�
Tռ�{�{�?6I ��O� %�=�o�:RA������ᱍ��v�l�՝�֝��xc�g����q�ǽ�O0���:���d#��5���y�ԏ�g� �����7g�Im�i5]PPpy1�T����ڟ�΄������lT�u���GGGGd��Im$/�{��5�ewq԰t�����$������m$��V�I!��+�db��w�����W����,�J��_�5�>��m⵾���?�����|��cI���}���*I��LGg}qg-ŷu9;$��Q�wj���������uZ�����5!�X-�yV��TP}����k~�ᙊ�go���� 8:::::::?��ދHHt(�^�� >�`AA�Ꝉ��Tjb����y�m�[��~�/߿�������~y�B��^�u������9�x�CX���(2γ� �n���f�_��*Ƣ���ww/ww7u�˙���3�>~���<��9�o����pg�,�*��Ywo�����wv�����;����Żݕ>�~�{�|�^�����8��G/��ZLR}�:,���ߡUm�.eޓ7�ϻ���}��o��y?|�A������7����k���1,���{ߒ䗼IR���l�}i5)��] =W{�����K1�b�2��%뗐��~�2�i�ޓ�߶�O-�����v��	7_�`sm_6��|vgT���K�6E����M��������̽��|���}1�+���w:vN��M��'ܣ_O����q�s���0�<���k������y �fM�L����]�KGl������ڷg�o���ד��ob]���J���}$�'�K辸��_Ko�ԸeW�$������tu���z���Qs����� ��l���G�E
@�/;�<��6N���Ke�%<�/���'wrjS���������D���6?��@����z��Y5�޻]z�Ԋ����Z::��mPs�kء<�5s�Τ���������ffc�=����~p��g�����)�%�O?����;w��4�Q՚{?�oM��p&=��o_&t�	GGGGN�wW�؄]]�+_���?z���$������{[o��HH:;3;�I�s�G�g�z7ux/A�)]:��{�2DT����\�)���j�}=���z����@|w���E�ٰ�"Iy�,�ُ~R � �����ԳtH��z)��oj��GG��>���=�x���=/�2}���4�o\��x~><�{̹���t��yQ�L~�z�����6̝� ��l�ǵ�Κ��{V�����\���.E�֤)>�Ϧ[ē��ie3���o����q�7�ׯV��I!��n�d;"G�wp|A;5��B&}���S�pOo{�x �J�d�]�v>���8�h�����o3��>*�d�EKGz?���s�e�o�E��Blc�[lp��vB{#�u����0��Ύ�������~��Z�{�{�]�/O,̽�d> ?S�)�դ:::;'�I$��#�$�37��z�L�73�O{_'�{���	٪�}����MM]PPy�����7w��M�ދܧBA���-�ʰÍݸw:|ײGw$T�u$�C�������::::jZ���|�\Q�p�mQ����������ې�uv��^{M���ը\����Z��D�i�3wuA�ԷVe�I)h���wu�t}�T����A�-��~3�kؾRk��y�m�����G���]���$�Q�wtC��������y+	��,YI��68:=ST�թKϷ[kCD*�j�$ϻ�6�%
 u��+�'�۹s��$97vl��ܶ�"A����61�-�����>lpttKHm�m�^���]��BAäPK��$tttttttttttttt/g��_m"����f+M޳�e���>��n��n�b*Ē.�]z�cc����$�����C��������[d��z_+7�r�E:�;�����kǻw˫l��{wX�6é!�!�a���㘕S��F�(�l3:N�H��ttt��y�ʭ�\�$��u���y�9��_R����=}�\�:�os�y/$�Vy���6ʳ����/6P��b�~}��G�=�����{���54����wgHY~����2�'��W�qb�}�|�;3W���wu-��Mo8��wv���"|�����ޖ�9�|�I��
�Ǚ��F{}�}="��=|��wh��]�6��g}��hIxհ����y�<�Ｓb/����{,�Fi��[a��b����=��+d��ko[�޵��H3�6��o3�̽��wxߤ��o���ޭ�Og�E��_i����zG}q[~�H�S����3{�w��\�1\Y��CX�뽩\�vF,�m�&=i���fq�I����n��9^��FogY�LK���Q^_j�|��>��#�N��ڝ�}��n�.�b����wr�Og�b�{��"��ow�W�L���q�~�q�QQ�w�wa�ovs��+̷7����v�}{K�/,�c���n��n��se ~��$X�d�F?>�t��-ŊK^��1����S�E�bz�l���3�Vzb}�>Ҿ���=��䶺�;^��K˻���ZG�b{V�����k�#X�ﮮx�G�F�GGGO�C�=�m��/��|�~�|�߅w��e�9���>$�Q���X����q�t��ϲkߖ������z�y�T�]�J͛U#�;���,L�>מ��>��w>���I����ߢ��7�m��:���s�����}�~J�*�/�č��R�+&$��:::;�9�) �������������u?~:E���:::w���GG^���6���}�_[I$��۷��Mw9^��}	��T>O{�H1�ԢI9IGGM��)V��og�}����M�d�󻧖�ݍ�C�	5�z�qК��(8::::;-ܾ�.�/��~�!���;�y�若�պ��[Cw��A�b�w�Z>��JH|��� ��󣣣���:2��Ko�aou=�L�j��Uݤ���^�T�wj��~�����������e�������ToϦܸ���I-��;_��V�F��WEϻ��s����}$�	x�������w�#�%>�w\�kɺ|N��-��I ���MPPpt�:���������������o�'N�����������wwQ���GGGGGGGGd�I ۤ� O�:RA��������{��W1+idl�o��ӧz-;�7x��:o�n���������������������N<�wt�c>lcc��k��l�'BA��-��[IGGGGGGGGGGGGGGGG}�/)��7��e�y�商�*�j��J�GGGdI$sx�ВKi$��A�Ē^�f*I!�N�Ա�g���w�$�QI����BB\�$��zA���߀������zKi$��A���������э�lttv t�����������ݰό�ʦ���GK��N�wp����lcc�����������������^�Yd�߉N�}�[���$/��,�n&ׄ����کem���������:+�������%oT���N�� �������$�����D�D���t����������M��{���w��>u$��Mo��(:::?z�c�����۟dOu�hvKi �������n���o1RQ�,Z�\�y����:=٢KwuI$$�I�zF�º$U�gk��N����� :N������[��[O��GOy�������^�.��m�tttttttttttttttttt�:rm�﷧��Q�������<�>��/k;8y����lt7�lZ��F�(u��wpޡ!��{�gt_z?}�㧼::I���������tcc�������������{/��8�4��OU%����m���H��˪ܞ���O�&��
lt��tttttu�,��[����7��31���.B���:|�����owwp�]���f+�'AK#wN��ؽg6 �V�E�L��R��CS�֮._t��FvgԔ�Θ��t�f�&j�ַ����ﻳ�^Թ ������<9�����ر{l�=%��N�Ē^#/�=�'��6�1/v��){�ܬ/oww;��4k��x�vU�������lw�{��=۽���2dI -�69�:e�y�>�~��P�����={ב���=of��!MZ�԰���P�R2d�_���@5�ǯ��9cJ�zw���vu���m��Z�]{���t�c������RD[���vww.�x�v��������{�S�n�::jZ���c_?�n�a���<M���߷��%����x�s9%>~�OcS�D�2�1|�Ϫ�:y3�rzz�].���N|�Q?sx�o�!���̓�Q잏�Ml�Ϗ���5$�x3�ˏ��|[��ڗGt��$�^3��GF�)u�׻����:u�b����`��UU�]ܺ���Q�u��� �ȾJ*�%w���,�C� ��� G��1���Z���Vi��#z��h��+�->�I�������曪s�n���Q�����Ø]��f.�5�u��T�Q�����э�l��������ƒ��K>(߻����+�][�S2Γ�H�b���߿~����~nk�)���d軗wwq ���gݝz���n��A���ڧM���z����|iޒ��{�e1��ԯI�ZK+���k�ܮ��g�K�6M[��G2��	F��K+k��L�3ãX�Y�n����Z31�K���6{���y�ww��11�ğn�?����9�+f������{RZ�ҁ��|�( 0S��u�̕��rW��zf-d��?�U�g��	���u���f�^�S�ȶ�������y��>��N%�뢓"H�tbթ
}���H�N�����t�'��Y������GGGGGG~��%Gd����4$�)�pR�A�ӟ=��680.:�L���lp���H::::::5���u�W�i�';ҍ���m��x����g+�v4�`���`���n��w���%���u�¯�g|��U~O��a ��H�<��!o���������'BN��! ��I.%T9����()��oeMAΒyyk�V����۲ZI%��w3O��?����51C� ���!=����Vt�hc�F޶�I$�}��m�IS-��ۧ��(5�|{e�l�e~�m���,;݇%s�D��<Y̰pt� th��'�L�T��T:wwu����P�����_����������s���t���� �ES�O�������� k_Њ���:����t ms�� D�T_ݠ�/���P{UMx�9ћ��|
=�蠞��UD�κ�Txq�Q����H�� Q�OAz������}��I(R �	CBR�4�1D��JB�!DBBE"���	CJR4��1)2J� &�v+�
=vo�SJ`!�7���1Q|4
���q{Pڮ����|v��5�u����<��!����ܦ��y���;Q�|��B
B)�� ���o�%O^��^s�݊ ��� b���qQ�|�6�'�$�2@@�JH� HT	)D�TID���(A
!�^�� ^��P8>v�v���֏=�^˷��{U3��z�C�n��h�]l��U�Q�vp΅�_OS�Z�;��̑�b��z #��߾�5�B"=����P<<��@6�� ����?�� ������������k����F������Y��@ �Z 	 g�1�ض` �(k	��V��N�h,�(��.�R(�@!�\�!H�?ǟˬ��y�6�k_�J�.��jPX,��Dn`�Ęn�>6�\ػ=tۅ�Lq�KMR�Um��­]U�/<�APUU�UM�U9^�\t:Ý[Y��mdzg�����jR�V����'*���������'�v�nӺ���cI���sv���C��'`���ڴ�ѓ�6�s�1����yvRí[:'�ai[a`E����*-��!�&<�ӈ�܄����� `�vM;����&�h"KU�Ě��]�B�{].�Z�����*�C��u��+��^:������[dܛ\�h����gk�G���Z�I`a�u��FwN��GQ�E�rK�n�؃�Ʉfb�ͳ��Mwp�sf؀ڦ�|g'u��(�����UM��@{�B=A�@�@]��=��'<�]j�v iN]�(.9s�a)@�\\� �eWb��5�*^������N�E{ϗO������#e�q�����'��pb}�'<��3�������B�Ta��1{���m W�����O�$�b}��I����dWd�4�'>cv�'��~��'+�0F���e(������z�7�\Xw��Wh��Z7��q5.]���f6,��ڶ�;������d�_�dxyn��Aw- �1h�'���d�K���`)�)�0F�ʤ�;��0�d��9�ϗ������l��z��9��%�Yn]˲o��lO(ti�)۬�\⦕�ힴ����D��F�ɧ������b n�6I'>cv�T+�~]��%������{��������~�Cʢ�dB�B�\�{k�1x���ċu��׷���iz�q�/�wh��F����$�\Y��v���kgF�O9Q�c�0&,6��~^�vI�%���5�c'V<ϷE��]��0�&�0���x��'}�m�q|w�[�ߗ�4�n��b�玡R6�j6�(ĂLԎ&���lY'�]�w�A����h������N9IX^;�C�;����鰕ӧu���0�@X�ݹr�E�h�_n�$���{���P� $SnŒqn�|~{�URVM\"WE��DBo���Kj����3�w���~=͂�#n۰e�V��~�o߽mҤ����ĕѺ�n&��,X s8�N���o�c�@j���j�<i�53y��֐�� -�*�5	�
A�_�n�$��m��6�8��vO�筦��m���q['�i���#ꓗ��5|}�\�{j:Ѿ�%qP��VI�qіI9�l���b�P��Ay{���\��w�5�$hr�ӶUUZ^� �-������CJ""?t�����~ޥ)Ie�X�0L8fVn�Zq��ɸ�ȝ�t��F�8C�8WgY��gm�]b�N՞�z2Y�j�:m�6Řnl���c�Egv�jMQq�����p�lA�s���A,�@��@�M;78;gp'8n�L]�Au�k������m�����mp���u�V��z�M�vĈ�D4\D�+���u݈=$��7h���� ��u�{v���ںHB�*;��;�lR��9].��c��>;����/o�>����n�����t�4j)Hr�vZf�N�����'ˎ��Tu�����A�OI�/fo%@��8o�����u�K�����m��~�n�\Am���5�K���p����u����l;C�)P���"�H���%����'� h�Xlp��r5;�l$��GD$�M�+;w��w�m�����>�tꊊ���
�@��[��3-��82sȤ�,/��p���vٺ�;tJtM��V����;��˸��i܄��#�MLT��oS!�F�������I�m�*�O���N�e�QSD�\I��h�Zwm����O�l�d�}�z 2\wV�,Z:wu� #}��>>=�3��v��{\MH�1�ۑ���{lo�����nV|��ϼVꌺJWhZ6>�^�Ͼ�������]�p�ԅ�l�
lVy�߿{�䴁gNe�.0��J��%���i`����}#����=#��$����p ��+"bЁ� �
6�sVݦ���yn|ۗ������9{�<ϥ��3�ooZ�[�S�~��:�C%�0V�)U�H�Q�F
�5UAi�"g۶>����w\m����߻=�{��m������2��Io|��Ѫ6#E�aA5���c�����������Դ)1�W,&�nX��zk�#�޴���]�ekJ�ЖXS 1P-�d�̉O�����!��߷�c>'F��%�ڀ"��$�(܄�
��*�C29���}� �}��0q�.8>����B���jǼ�n}c��rm��N^�z}6�i�fi������v^�W%����o��v��-�'X.(ݭ�x1���q��v��{���F��m� a�5��Ͻ���iuIJC-�7C�K�8�l�d��&KN���/���/j�|ꉢ��M�,BI(�$e71DK1@�V>�v��n�o�������֘��18Ab�����פY�����!���5�e�e�,����%Ϻ9z\�����)=t��M�q��${7vǏ������`��m�T��N�Z�r��Z��PIIt�X���t�'%��/5�N�ź�uz$��]b������N�/;Ga�ʫ��9�n��u�������m�����4��<�u�$V.��ԠUT�I��O+��.y�hۍL	6m(�P���n>�C)8ڳ���g������s����1eR裇Mv�/gہ�yD���c}��[庆o����BF@�$�($2XHq#)�R\i�����%��f�|�������}��m�=�vaڠ���7�1�G�۸�F�^����j�&3O���g�O�g�d�|�߯����>�=;����Ah��$��:� >u��o�c��s��������BP�3y��Ͻ�{֝��0S]T���g���B���
ڰzz�O�e��s~���}�q����ؽ��/$ͦ=qΖ�{NV�����e�m��{7Bh� �Fƌ�+�K	��lٖ�
�͡F���-j��W���[M��<\_�!�PBɰX�PD�	"6c�H�9^��C������Q;�n�ctn�R7M���9Dfn�����4mQ��w���Q���J�BE�ء\]BW��3}�l��mQ~��Y��=��i������[���o���7�0a��g��z�����dN�=�GQ�D`��@�	&�%;m��L���疳�￿?G�kk�{�u�%�@������F #��	�e�jmp��|������ʽ��`�k~�=�F�-˹LZh���f@}�ǻu�ݕ���c�߮��hg����r��r�Z�N��&�4�e��û����i�G7��r�����������|���7ۆi����ϟ{,�d�m�h�.�֕K�d�!( HI �Ң�%�K�����}�c�|��i�Cwm��D"T�-���n�^jmR�{ϟ>?}�W/}߯�j��?O��L����oۆH�ｶ?o������7�(,�����7w.;�����*�}���
��,
w�.�����{>(4v�����T4��ֶ��`1�N�4�hD�n�	���ۡ��<��, �{w9����ۼ�袔��Pi-&�A7�jK�^�N��D�,d�Q!�$�,,q��ִ!Щ�w[�kK�P)�L��L�,�a��#��$�0�H��i=6[D��4�Ki��Y��4X���
�4jѢC����I,X �9̳4Ef����0cD`@ִ�H�U�7�̌��<���V��Q�PH�2�Zf��[��D�1��cG8�c�1�1�2��e]��n�+yv�p��aM�J��i���ʛ��<\�ڣ&�l�.t�S�0�&0�	Ӧ1�ε�kZ�i�kZ�kZ��	h�c
�c��f�[)�A�1�cT�1�msěv��N��[��]�\$�؄MV���r;�,v��x����:+��U��Z�/mcu�.��pF8��VB�wZ,Gigvݷ�:B����@ܘ91K`�N&*`mVl�F�L�i��ZHE��1�`��N�mrճՒ��a9�lq���;m?qq�u�Z���ݸ-V�K�]s��z妫m��O/l�8.ڕ�ZvZ,�� �EC"�+*顢"˖tQ�v�tk�@	��s��ct��l��zM��B��wM��.�u��U�2��vN�S,�9�kZ�uF��!�e�4�C�ͮ�l=�r���Dv�v�N�:��kt�jڶ(b]uD�W����)^�ŗdQ�+:��݆����<u��6+�x��eֵ���[��v���Fv']�]b[�]��t�m
�!��/
vT�p�K���S���w�.gk�=����� CC
�V;Dq;+Q�(�E�%6�J댻��X��C!1XKvqb�D��tuqŭiqgZ���'W[C���.��h��J�l��Z���ݽu�V�H��_e�zE�ε��Sp �j m����(��K��e�3��[�!2ʇݻ�+P&�i���� K�7��&@}I������)N���g�):��{�PFJ^}���H7���.KhC�؉%]� ����;���qJ��n氳Ef�h�Q��{N��s盓�[p����������E!J^��~愥)3�cOEk�H��	� [�E�i���N�\��k�b���hJ����'R4'�}��`�A������T[�JSϵ���hJC����G�m9c	�����0�j��k�Й)I������R���w���	�����P&���v�pE�wm9J� Q"��zx��(n윕QG��h�S��}��;��/��G��tq�d2���a�_��\r�����k_}�	JRu�>��JR�ϵ��	�v��*W�xw��g��oJ]���mb�m����Z�J�l;�ntm�� �p�+U��b9E�up�6-M�5��b�6�����ٳ�=���ut�%Ò�F��.��Iv���}l��*�mѳ��tf�9Kp���8J(kb%�.����FhV7y�9Ϋ4>?��Ɔ(��8pH�eItM���oy�	@�w������9!͗�C��mڡ�
Uq�x�9���.2�H�*��+��*�g�Ɲ5T�}�=5@o�GI�i)��$±�v��ct���|�Lw���;��o��)<��{���JS�u���!�JN�=����)O�����c�(, ��7,%��ha�k�GR���{�8�)F������P#T��}�P�a o�{��AAc�e�Q�6� Q5Vl����5TH����Hy�5)�����J��˿�߰z���̽m|�� ֵa���<�$��5�؝@З����	�4v�40�@f��ϱ
����A��R�c�R�t0���O�Uj�#�Uwe�5�����E�Q�1(�\�������{�߷����~���	��S׾h����Mo��"���`�*����R�A1��
���Pw6�J`�{?7	XH*�0�?X��r�`��Q��������5�VE���(6i��cN��;�7s�N��d�<��<�'�P���
�d3����Fv?o{����~�چ�P$����U@�h}���� Q"�����h�+y(!Au���Z4fθ\�)O����X%)I�~�߱;���ou�}�u	I�~�Cۈ� Q#}���(�.�-ȕ����h:��{�'P4��f��4%?@a��b�5@�+�a�!A�~��8Dۂ� H��#v+P&�{��Td��$���t}R����ﳊR����Ӎ5@�?ykP��@%6g.f��SP��w��_�^��֠�,��m*V�����Z����i��)������ Q g��rP$5]�7�	�>�5���n���y{�e	�LZisDm��x܈�LLD�+�MP�X�)��M��r��
$P���*�(2�_Xj�5��tt(�ŀ��؁\F�(JN���A��w�����n���1Դ�C ����=MA�{��}�
�P������%�hd�d����%)�8��)>��߶=Hy���tk�`�����5��=JS߁��� � F�p�n�T	��ݺ>��JS����Й)I�~�����)ûx�!���42Fw�����MP����	���?�xʯ2y����+0���a8�"�7Y�{�VZ�͝�T	��N�:@�D�ѯ�d�.�I3���<�&�Ιv��mԘ��!$X(2�^򡆨 ���9��R���}��:��2~���T3�:���7c���=�z��/}�[�_�T�JR{�揯�:��<���R�ݒu�=��H�.<R��t��K2�r�5@����ߴ�@Н��︦�:���7�fm ����p:���
|��_(@i��%�+%�c\Mc-g�J�O�w�~p����7�'R4%��Bd'�5�}���:�&�/~!/�� ��Wj�,Ab�5@��cyP�( ��	*9% Pq��1�.1ݗnЀ����>��jC��=��߿hz��>�r�;��2˖0Йl+ ��˻-��0�#3,�Z,etޮP4��}��!�d�v��߰:��>�_[�S$*����I�����R $�6�ruA(�=��Ϥ�R���u�����5��=JTyoX�~w���V0��ɂ�\r] Q"����B� Q }���z��0�=��o�)Hr�:��~���Z8pAHr�a���Q���A�~}��R��w�1J����"����h
>D����%Gr��t��,���A�x6�e�f4�%��3KXY��x:������+�S��f���8�r���8�Nxm8۸	+ZH�c
��nVV�g0�8!��]�l�:�iݦ�
�Uԝy�ݰ��Yh6Ғ&�i�W��߻�(���t��%!�0л�c�Ǆ�h!�{��!A��H��v�$*8rLn���� -��֘�h�>�����ܥ)�����&��O~{�����D��t��f#����J���Yt�9D͕&	D
�.�vX�����~��)J}揾⚁�{�tj��T�gZ	�=��z����r�2D�CuXEj���9*�����5�؝@җ�f���%A�|�w�5@�>�ZH/��tm�8��)JN��G�bu	Jy�>�9��I��}s��JS�����#o�A���y�%!K6 �@�����P�@Ryߟl�N�)O��rB�5@�o��V(��;��ĒX ƥ��t�Y��x��r[$�O;Q�]II�\W]Nd�+n�M�f���=�~?�,�)=��}�R��K�swئ@u��y&�� S�	����L�H^lU�,�v5�妴�ǩ��qλ(j��to��А�v�]^:(�)Ske���m���MF��E�Ɩ�`�:ЊX!��P:�e����h�P&�$Q����
$P�0��M@�wߺ��N�)K�=���)J��v��V@���p�M� �� ������~4�5@�O�0��)=�=��0:��<�^��S$h{�P�#Qh[����Ӱ0ѸrS�>��L��2O<�`y�'R'�h��)�KXd���~�������F� I�r�Zp�F�R}�����	Jw��يP�����(a���"��'��h}��D��m�z��gW]k���u)Jw����(J����z݂���W[1��6�u�P������Ͽ�Ol�����>�	��:�<��R��������'P����V�D$E���Ē+	����cyP�����}�r�~��v}'P4��l���M�{��K��c�gƳ���JP7�{���.�R<�ΝJR~}��?0:����5�o�L���wz�a��n��'p����]�2[�KY� h;�=�~��R���kߵ�)�^�����k��)K�s_����8{�����42�G$��Mج Q"�=�\R����5�؝JR��k߹�	>:Y��iʆ@��ѯ�8`PX�9k�����r����I�.���"hF����J�k�����Ad)+���!A(���;�j�5C����h��y�᜽�^Cu�>v�^�P�J�%��\ 4\��^r['/���r7�I�{��JS�~���k�߾h���M|��HpN݀�bĳa��(O<�/~���	���}o�w�JN����I�	�ow�&Hxwx%ȫ%Iu��-c.�T0�i;ϵ��Д�'}���:��������<)K����:������)Ok���
.��Y��ĺ�MP&������)K�>�|R�����>��A W���"�4��s<�.X�AI��Z�pz��;�߸qJ��Gݜ�ִ=�,���U6�y��T5�.�[��\{'�����ćÜ�S��_}�	KAI�k�z���=��mG�ݛ$||����yQTX%X-�j��"�4;�b�O]@П{���`�������R���z�M" ^����60���
�9��ܥ	ߺ����]����GR��~���BR��;�>�~����ᣑ*@�� V�H;�+��S�����@Ӓ�~f������5�}0�a����.�@g��	rc��8x���T�=�(2(�y���z��<�_[�!1�� �Q(A�P�XbH"�dB�)�
����JP%�8��D6f�tVn�ZqӚMl��p�z��a1��A*1�ݶ�X�����8��9��r�qN��j����yܵ�^��6�5<S"Y��Y&�Kv�{=:�V`�����k�k��K3��a���v a��n�l�LX'rْ���P&�C5q�UXE@�i-<�yF7)la�;)��,kp�[��͎�������F�K'�y�������=��jC�+�t_n;�,���'>0��34��"��p ��R���C�T	�r��)I�����N�)K�3��)<�ǧ��4(�}䴐_Qr�|D�p9��5)NG}��Ϡ�R���~��)Bhf�r@�T	����(3@v��Kc�2�0�-d0ج5@��~�{�Q�J{�G��u	�d�}�}�BP��Cۯ�P��	�c��e�%�D��Z��T!	��y��CH���=�2����Iԥ��{�߷�	�9o"å,a��KC�,b��22�����J? D�WM�ȝg�J9�$=x֨���\���o+�s��P�(�����P&�|�F�P&��q�#e�`�
�����/ӠӼ%
�I�M:Q��6����-��� ��!V�(�P�ì�Z��u+�I1 E0I��̄�5'P`�a�
:mmd��b��gS��fRH���)`@IACEI1�Y᭸t@nDmٌb`�VQ�1j9����9���|n�)���!&q=ޞ�RE�6@ɨ����J!P�Z�#�]N�).s6�UfBA%�%��0D��7�2���w�9�������1�e�7�x��-�k���!���(b�)!��BgD�@aD,�C0RP�&��22��	7�Ǜ۠�jSR-��4d5��$�Zka8M��l�ac�v�d�j�:vDA�Kwa�ˑ��M#a�!y)=���0�8�V4��r�Pe�(�H�l*��G$��"�p�[�n錌7k��=k���WDh�����ׂ��G�2"F9��k��F9�p᷁+@u�s��
G7����&��{5�yxw����"�Tj8�T�;a-�^*�g�ڜݸ+ml�����l�=A��*�T�U�]TX��TcT�5��|:�S�<V'n`B'���T���aW�[t�*�2\�n�{��ñu'1su��(qf����#1��N�Y+��B�qx6�}�Sے �] ���t�qQ�k��J����헎dQ��h�6��)ڞwWq�m���ݼ]�� /;B�S�3�`l/���Emۅֽ���c<u@�.qκ�+ѽ���9��X2T�b���Z-��	[%A�P
��WXT��s��t-G��+�HT����k���SU� ͂;mT4)G	�,P�n2F��n��nss�-�Ѹ�4K�v�U�F{j0y��PN���{��?�"t������]������� ���~z�o�w���TՒI0I�r��ZJkl��&9nӗu�8�g�N�<_}���M���Z>�-��tn���4�P��&��Tq��]�`��&��6xw���_>�w��Y�v��a��f��5�X�n5�MP&���7�P&��}�&�)<��w��JS�ܾo�\�ԁ�\x��F�� )�j�v�e;�߷��������)Os�^���C=�yP��[�������JGuBTH���B��k�kM�L~����wt�k ��Oo�j���w�1ش�g'���d��=��,�:�3����f�i\"�Gh��wf�}���a�ۅ�ĆM	y�a+�Cc[hT�*T�|����s�̐�-��i&��ݺ��l�&�����VZ�RQ(�+0��n� {�Ǌ�yϱ�l��{��7*��ڑ�̌�'>ן}���c�B����ĳRRp�e0�"��
�&K#Ҥ	���h�k�y&$��_�	G���*�j�̥����T���������0�H�[��߽4�#�ѯ�" �"Ua4�j����䇵��i�ks�f$��ǾG��Ŏ8�x����%�$�����^�D��aRjĴa6ٱ�&�7Z�#sa	�'ߞ�� z�ws�䆒������J�^+c-�M�ۨ;����ٛ���c0�ռ���us����>-�ȺI�������V]�j��c���!��}�HA�?�����$���M*�]� ,��d�����I�[��o����8o�(�/<����Y_g�~k��yM�9���;	f�=�c��A��}��sôt�];C�C����^,ËN�4R���m�P����^C1���ݗ�LyWj7���MEHM#w��>o0�:�Izh�|�|;�m���I	jE�\AB(�j�EEUɀjӝ�g�s� ���L���!\p�9�I9{s/
UE`����j�r��s�3>��_�#���?E�+.����W>�z |���mp�}�:e.�!�o���cSR6���P%\JV��UD,���_�ĝ���X$�����1��p��h%�HZ��a�d%�K������N�s�W[`����\���M�������W#2��eti4�B�)c�v�n�J���6�/{��
=�`�:ca�4"�tF���E�\��;,�b�g��#I,�ሱ
 |��Uxa�ߗ�l�����
��7m��L��~��>���O;tO<m^����E Eԥ#E�ˈ�!w@?w��'��V{k���j\K�M\�?$��mQJR��2��������=�����h���s_�`Z�Sj����n��1<�0��[�A��?w< �����}���UT~Ѽ�e�#�݋i��,��5�w?З���`��>�w�Wt04f<qXP"���!B����}�HW;�����\�?�ﾏ�FF����Š[�Y'���|���?� \>�Fs�s�lٙiP Be�$�.�}��K$���{���l�ܗ-�˶��P ����0xz�,��,��3q�,L��@������ӝ'J��������l���M�>Ѥ+VN���l�)���u������5E��,�oa�����kf�
�!G��(a�4�m��[��S�Zo$=���;�������$�������0_�-�ё�'|���� Q?{�Ł��oF�:�n��J���k.���ӻ8I��ް�Ϸ{0����0
��?A���+5w���$�	�)��\y�G7k���da`Ͻ���몯�s��j��^B{�Z�	B<��.��
>	�,���D�,��K�[���,�J�mk`j�VR��R!"��D� !$�<���|��['=�y�<;Q�Sr�K��W��Zi�ku��7a���+�HD&w�%T�X���^ڎy!����4(W�B�4y.�S���;���P82�YN��*Fs	���/��#UB��Hz���YW�{����~�Ϯ�J�)� M����R �p�v�R1.;���d�q��U � 
���/��2{�~��w��Lpa�Ƙ�n̎E�H���l�ק�H{[��PD~��ݽo}"䆒��ASe]�%����3ϩ�DڱdLZ�G���]zW�S������p��
�@�{�/֏�~ޗ���m�ü�ħ	XMVNe�A�"��%B������
ER3�1��7w�`�n�~���EM�����L�P��!f�,�d�}齟�@
�T)����۽���uu���5�� �4�؃.�	�{o��O��[�� A� �GP���� ?�C���d������z��R��M����� ��UDO����������[�~���S>�F�}�ȑTT^f]��FEb0]�n ����U���6Mt[���Gg��ef�3f��a�� ~�U�o�??7��o�T}j}>�u���4%Ut��z��1ŀ]KT4Q+��rI���ߢ�������П?� �������~�7z�a���U�sjAM���>�^�s��)�� ��W�ߟ�!�@��M�-�<x�������D~" ��||�e����P�O���L$��w[���������N|O��
%�N�y��z�|�u�T�U&O}���*��?:꯳�﹫�t��*Vb��r&d�Y%��XJ[{����W��f�u�`�B�*I^�d�����р&�&�\@�5F�O��m��9�;L{v0��n0q�\3�S�q��<n��K���f�X��Z��p���+�]q��&�6����];����j���h���/99$�'�g�rs��?��.�%��W	U�QU*��{���9�)F#	�!$p�0I��V�*�Q���������>^�鄟���g�M�,�n�<:�n[(�cT�5ɘ6��99'����%95��U��r�b=�L���?|B�����T�SE�­R�*�7��?ģ���`v���A���~�������ELx�"� �s�['=��'СyՁ��y#��J�R��턐� jG,�+�[��ل�秿c����ߢ">#���g3�&f�ʹ3 �&a;탭�+	��[�vΕiM�< h�k�� �L)�����y3��g�����.�o7��o\�=�j�����]� ���J1d!b����,��A8#�0�9���H d�8!/$�����e�+�۰��][���;�����{�)�(��uf�shMR��5׽c���Y1�{1�N������=���ap�uǞ�7�!���W{�ð,�f@�6��h�ծ��9����b�bX�rd���v�w��� r��d����m���Zx-�w�������D�D~��(}�����@x�w��[@PZv����[6�7n���s�O��[
&�V>}p����ĸ
�.�1��	�~�B���?5Ȯ������U���e�TI �B�+*��� ������￑�"�M~���.d�
�^��#�M��ٽ�>�V�kMZ�*�K,b� d�KH�e��Ͽ��m�~���O�����w(����(��20���֜������=�rr�IU)i�!U!GF��H����K����y ַ?ё���b>���E��ʚ	�U0X�{�}�n����� ,�
�2kC
�C4�f� �5�a,@%�#D �h	Kj�0L���8@bNh�@�6�𸬨(�x�~� D ��`���$�`!�9�6{�+���>��Va���qW�U�HA��(Q��x�_�_�Ɩ%x�a��ϼ���]��uW9�?�DG����t����~��=$�6�ʒ�AfӁ7dЧ�@�(V�`B���}~u���|X��>y���C�q���]��!5Y�jQ������� ̹' ���Zq۪��M����a@��n��f��Y���T��H��=y����~z�/�_ZM�ȇ3Q2M��)D�q�q��	�a۶dX��;o�����W�(�����������ڏ�W�Ғ�)�Q1uB����~��������8�]��`o�wg��v�?�2�7�v�J;D��|����,Q5�'�D�u%�P?3'��Z�g!1#H���y���n}d��$�/"ӤJX �6�{Ƅ;�ՉIH'Sm�-2���o�9<�;�fXXs���h�،�&;M�m�{�S��ĕ104��tA�p�$�F����$�%3@/�؃�vY·�b��k1�����,���7}�4� �1��c�01� ։�Ҏ����%͹\�a�=�W#Qiˉ�؞n��u�XG<�D����Gf���1�� c�4rc��k:ִֵ�ֵh-k[e]k[kel�:Ӈ:ֵ�m��ֵ�=%=v�Pl���[h{���K�\�S��;iv�Y�X���
�jժӹX���ɴ��g��+Q��<�4���70mV�L�;���氒�-E�m�p�d˷d�N���h�bcVXA1�u��n��Is]۫ܘ�۰3v��,#�:4YOEm)>��;NgZ�&
��� 'Bݢ�9U�`�h�*�1f��o8V����^�Ocq)��C�ɘܺ�<sd�-;����<�t]b��a�	��v�%]��bP �oҁz�2����Upc�E&�q��uʰj�pR`�v�q���b�!<��x�s�=d�llU�f�vv�ۆx�δ�6ַ.&�lb��Vv�k\6�ε���m֭u����'/7>p��W;E��E�<@n�3@�q]�kbD��>�ϑ�;-׮��ȁn�,<e1@[���Y�wF�Um:�ۂ<�b9�sV�õ-�y��R�iNVɳ����Z
� �9q��":�mZm��!�e���1t��5��5&n�"�b2��e����D;Q�@�Ms}}�=��b����h����(�T�`�	^��t�����z����Ȳ���W8�&L� ����~��w�`=��`�L����ܛ�4��U	MYvw�n�۽�	7C%�[K�����M�׋�8�TU)��{�ɴyzg\�A��͆snUSu��M��w��gH����p��	��\DDJ��W��n�=������
�Y@T �oO��g����r�r��n���X�ɼ��|��됍���$�n��U�@�����?�e��YSSu�j��6���I9Ѽ�
�n��!��Qv�nZ�,��1Y4(�zwc'����>_j��i(m
"��?O=�n�\j:P���\-�fPv�hØ�V溝�gQ��&���t)�(����(����l86�v;V6�x���=���o(�Ս�t�Ȫ�V�GT[@A�p;Os;�.�R.B�щi.k3/ж��@� 74�,*�����������o�bv"��s0�庺�%Z��I$�`r	"j�t>��A����Gl)�ߣ�""<w�~��ﾛ�=���I��2��7C��ak+��r�#t&PL����ߣ��+Y\�����>�e����z������}%A0Md���TVft�w�?~�(���`]���ݯ���1Hҗv�L\h��	?{�}��/�~T ��hUS�__。{�~6Ov�5K��b�،��F��+$���v2wX��P��Q�hU ��߳s2|�*EE��T���� ��K�k�K;屗[�<�Q��XL�	H�,D�(8������܉߻���Ǻ��q���,�s�E :����8JA���WZ5��ޱZ�4�bgiu�φ��LKM\[s4�f{+�X7)I�v�/e=�=_+l5�kr�����T��N�U=��\��vͬ�&we��9�[�ײ�r���jkE�,�_��P5��u�k����ﾸ�7�M䇺a�����`|p�|��["�
�V�-�7��U@����#�\X_|��A��9���D~���U
�g��?*�F��W�h�����h3]1����w��y&�ȥJ����5lٽsR)�!D*�,���#�B���d �>��7z��Da���d������,y3�b�pf�����v,���ݤN!cu&���\���5/(w����r[dAA ��0*� *� ~��w�_�r澴��<C�7QD�c�s|��a0cmط;2j��뻻
��"��ms����r�yЋ�0��*�=�~g���ع�?�_���+x��y��w�Z�LW��Ъ%Y>SW}���j�D�����+���U ��Q��~f~�~��.)�Ӂ[%�����|���g�P�eoW�d�����R�T���MVNZ����:���4��Ph&E����[�?����C��)k���O���)&�qڴбd����$�@|/��ʚam��M<Nš�ۚ�Q*F��G��hP�����>����{�ۨg�L�J��Td�* �*���6�vԾyo�Y��[o���ss�g�ߡ|���ka�Q52���J�J��{-��,���`4.�7D�!����M!Fb��SFM�1�_ v�y�����}��vc?[$����3�Ἄp"�� Wq�V����oΟ�!��ŀc�� &w[?oj��P929y�\-XY����fӴ�����0k���4ĢJi�0����	��VP�����A;���G{y��7�SQ55UL���YL��ځ	,��#�1��d����&�Jnlk�j?~�{���}0��9�����M�Ln��Go;�W��Ӏ,�<����I�J%U���DԔ�	��~��܁��C�<���;��m7ć1;�yv�a4({vq�I�{z��~\{���� �޺�H$u�r�vGCWU[���3�0�cv��.�MXԴ�jǖ0�D���mg�M)N�<ֶ ��=8��G\vП�d�8>�R�B`u722�a-���.�p6|�6�&�:Iy����M����It*� (W������o(�.De�u�Q)X�� ���=���^G]�Œ���wetX����J�U!S���w|�"�m��^��Gڎ�0ʗ�<l`.�$�Tj'�D�T �@��Y��s�ϫ�H{vq��I9�޼'}��NB��l���"d��Y�m�`!��6k뇈����������8�.Xv�PFfa'���\4�)�����̩���������F"���7$l�(����N|���ݦ�A�����u7$�3Y*���w�8�$q��@�a�"�q�`�����o�/J��ߣ����:l�9+�o$f�&���^������rY!y����@�EU�˶�$�3�&�)�ﾗ���;x�}&46�H�:<X�pG\�sO:�]�v��7d�9�O���v�v�����C�V���U3P��A�m���� �������߈��_}��F��3�*�Q�N
-R���SyDE��f ���>��uք�%Y%BK=��3��kY���\�*�X]��J9w'k\L�]����wc,=h�EQ��y+&�T�W��A��`Q�!aF>�ֹ߯��d����?�~��(}�ό ���Ra*i�J�\�$�7���c��+��x�^�
��W>��[ޫ2�2޵� � ��
̣�����V�˚����N���$��4��z�,cʃSf��Ws8�UYU"�=�l�������`<�s���X%	l�������u���ߐ_�IIdF�,'t���޾9�P��J	 �"�*���_o��]��y%�u6�5���r
�*����<�yn��O�n�a�T{���@hP#�D�?���,	7�����FwB��$�)�Iu�j���CV��C�[��OĄHKw翟�����>?7oY��SL��B�'�c��(;�D�  �.uHXb&�,��X�UH"hY�ӞH4�v����{��	�u�������y�T%�#�Jժ���&��3��/?Z�_���Z���3ͼ�V�ܞq�q"�B�WX�̛T^ �����?G� ��}�Hk�����l�������B��UiLʙ����{��_���>�*\� �����C"@�Q�#RF �XXĔCQ��� ��'��ٌ����[?oj��P)X��E��P�0>]<}��ou}��=�L�C]���g{�H\�K1��N%$��9�u��L̼��"9��#h���HT��Ʀ��g$�}�N�n�[�[����%Q��0��c�y�[
IV;21Nܦ���s�7r�M�V��D~�D������U���U*���`7�9܆n�a�-n���~���,"k��p�����n���m1��BT�ܒ�����ͪ�EUYt��0F�
4 ���?~�N{�_ㄜ�N�d��*��*� ��K�l��2�C��Xxz�]d�]�8��M5af)hKH8�W�a��j��UW���^pݞ8F�[J�vr�p������I�Mx�7+A����6��cki�ڙ�
�mu��nJq�!5�XZC��`ْG	�@�!Ғm
�9ЯC&�듴���ED����g�b'�rxڛ�/�9&/�K<׌�R3X7�lBʖRr �2�D0�(�$y@{�Oڈ5�/�v��k��%5B��wIEȑ����x��GXBS��ꛠ�������z��Q���`���Y����`�V$30�.;ׄ��� 7[���p���5B���e�Œ~��r�u���{eP�}y�AIo����㳣�]������9�߿~��]3�A�w�f���H��n�!������աI+{�m���$����+	m�b̗�0X<�J��!��-�0O�߿����=�k i��\4�A4aS��+������{�[��>	�
�I��I��5��/���X�! �B��#�0�!EP��3��Ba#!���zC'#p�aRf�bF��B:�BA�T�Rd*�ytA!0��Ͽ�^�t����7�{�g�nｧ��-T�[`����\n�4�Z���:���K[���ՕZ�`
�U��
�uPVݺ��U��m�m���t�z�{a:�lQ(k�)�6e�۵��D��u��m�0I����n�۩��4&Yh�X�X�����pn3����g\�u���=c@���ݖ����Ζ���s�L� ���M��]��	�2<��6�&+��ױ����4�lh�
�X9�� UVؒ3yrC�j+�ɺ�4��!�`�(��9�{0�
\�Ξ�be#��ݛ�؀�V���O#R�gn:杫ت��:�V��l,dnE��*�����k�3�k�nt"��gct�j���3ַ�T�J:SP���9	$�9�Ns���� %�ס�t���}���,E{n�e!@�%
!MQB1RQT��(� {���^t�a���ݦ�[��Vʆ�2o��:ױ�GϽ�'��ˈM�M�mny9�޵�XF��V�������kp4�%�۰���}���z���'<֑��y���k}��>n�[��Hn�C�$3����CB�&�+��)]T܆�i�������䆾w�~���:���4��)NZ���U7�|��}h3]7�xGKu`G���$���Eڛ$�P�B�������r�<A�ua�s�_�Db��2$a>��	6�N�Gg��1ֺ�=D���UJT�QBJ��<׀i��	g;o$��>��`6����%��@	XYEIHA-+e�j�+$���{>��ֈo<�
NY���Z�SV�
�MdDF�k-�p��Uy��o��Q�!!�!,CD�&(XRLQ�c�
�yFF����_��L2RBJ�	�H# X�I3#(�E�2gJ
�A��%�ǈ��� ���
꧹!���<鵀����*&&�]\Ҫ�SV�;n�A˛�>�LO)����Q��7T��R���!7Df&���=�\<Z��7r����QJH��ݶ��N}ӹa'Kc"2��P�u����]=�I㤪�f�
I�����u�$�ӣw<�ڷ�-8
8�텏	e�#�$�Ȩ�a4�-�%� ��XD��o�s�YI{v��A�mRTQ5s6�̩���=���Gs����l�������j��' *LNe���	��Ǻٻ�=�G/�g�_ �B]��(��(�	4�.K��� 
�߮�N{��b;���"�Yw������?�����鿋 z�܆}���;��Xk��ʒ�˜��9U*�0�����K ET(U*eM�c?��P��G2���������rrڰ���A�D����QU0 �^�ݢ�<�y��su2�ݦ~�yw\I��C|Zv���Y������'�cz�^�;��~��>������B�vTT��o��������	p���&���A�ξ,�u
f�&o�+���n�9���$��8�?��*���I/�q�;eӻGt���
�W���[m��/b��]X��dՐ�����֞1$����7Z����N�h����'���N�Bv�fvE0��k�ra��wK�ͱ��x^&:�Vf:��9��M6�5��7�����_���}l��z�NF��v�W��$����o�%�=9���D���Z��nnMZ�A|����|����������M�L�FU����G���|}���ia��F4��w*�*�����%�,�]��y�y���L�&/�r�S,��C	IϜ>��^7�C;���F�HoN�r�Z�XVED�E����L�5�[��o��E+���0��xj6aj�Z. �H��<����w�0��?r��rkpp4TF
�)J���a�������̝m�ra+�:��(��R�T�R�\�f9���=��G�o$�bB��ʩ���Y�A�u�`2�
Ia^�i2i���ܒY4�99ke*ש͝p���a�I�B�F W�]�	�>}�t����6�hGL�D5�j1����@z�.q߿W�l��ư��C~�=��z����x��_ث���
������¶Y���6�9X�.�#�*�m�w}q`�=h=����b�w��˗�M`kn�I�'���q%��0ن�KZ�5ܛ��%Q*�Ŧ]�Q�N���"}�Zʮ�!uTu�7�n��k��Y6*��g�#��"m��?�C��#��������0��N_I��o)c'~c�l��x�-([KH5��\s;&����h8Xn{w�~��{=�Z#>^��[L����©%BJ��m�h�D��J�ē��։���$#������\�n�](�	�VY*�i;�s�����@P��\*�� 
�Ø�3��5�	^��u��T��D�x���3��h7��, =��p��}�����F��wm3bD���{��V�� ͝���i�a�sh�5I5��%<P��lh��XC
H�x��^��#V��f����**��0�]���07�����>��[st��W��[q$8��QJ)B �)���<���oS,��+$����;��<�tY�
x��͉Y��-������#����>�wb����&|�~����.��U)+��7qa'wvYO�}����B�
����f^b-v��wOs�Pb��ne�nxO� ���>��=�S�2��-��#�@�ُ���ӒDMZ���UIJ-��y�LھyC���ʹ��R4��V���)4�N�3����O��b�6��lëP=ć�4&lw0�VA�\,�-��Kf[��u��~|��^�v:�X-;��3�M䛼�AJ�B��v`��$�1����=�Zi~����N�����G�@��ƍᰯ�����[��v����a��򤦨����R���Vw�Sy!���c��>�+1�p�aNTL�TO[k�mK5@m�a�i��HL�X�g
��1�t8�v ׅ���]-�S���q[t�����8��]���e zIv��.�G�#c�͝���j��k,�nI`�ֹ61��[��Pz����pp>�&(��pEp(�80��{��"Da7�x���M�rr�%zh��Ԓ��Lʥ�*3wq�r�]h<�<��~����v�L]�q-F�LSLC	�"RC	�N|Ǻ�:��vHg�[��J}L�њ}/�U6J�����"�I�w��~���g��/7o���=%�*��LʸT�������o�T�k�^ޛnђ�-E"�'0/�y<Aޗ�������/����o��B�*HW*j����p
ݯ���;�Nŷ�h�%eKD#q	�&���U	 B>�0��`J��e�1��QR`�.ofU*�5�
`bgk�\R[�ޱ4�۞��hGaXm�F ���L�oQ�)�sl��.̹(h��o�{�%:��)�gPݐ��7j��
4+0Y2��L��f���D�L��2H�I���9��<�弝��:e�poM�Qj�D��n�V���<��~��wO�+���7k���}DL���+��B����9�w;��O.��;i��;��N�㸑m�uh�}Ӎ�~��m�{�\�I]��XG���.Ғk^fr��xq/�g$�"�H�Q�h�C�l!`۵mv�w����;f����ELi]xN��elei���1a{&�U�*f�3�������~�Kޭ�|��P+�EX]�8�I���Ь�  &�ͱd���M�~�M�u@ w�q��J[�I.{K��n�/O��P���0�z^#\�$SB9wx�)����vw�d���߱�5x�[-f�pY?�D���wW�s�m��������<K0��)T�$e�p
�l:�v*�Ƿ��@71��j���z�f��Gx)׷ �J��\�)O
��v����v��`�D�������I��˒�EX������v��v���<���5q�;�si*�W�j��nh��k�w$��a�@=T���A����mA�!T=D�"C$0d��$0�Q��FA��h#$
q""����B��+'�$M�`�<d+��!�i\�ֱB6�!L���u.�A���Rҕ�f8��-���3F:B�T�V��3����$$�T�M4���`-bD�F+�A����d�А��i`K"I�d(BGC2S�M{���Z�k�pZѦ�]kZְZ�m��r-�Z���F����um��&�n�t]�^�瑝'\���)U)s<���i�kJ��kF4rc�1�4rc��1�Zը7Z��Z�,k[mk��5�0��1�c c��ۊ�{d�Cf��SM��m��N��ݔ��-�ٴ��,iz�mٛ9E�@�,Yz�)��d�Wi�m�ll��xn�����\ڻe�����n5�6[sL������֢�rq�jaԏsX��"�e��7 '\SWv�;uq�[U*;��m�C;��h��:uC`��2[9��U�%bZ���S5����Q��m�y��bz	�K��a1@���tx�n-��<�����iU��`cf�r���A-�`^���i\%5%��T�*0c�+�u�6�[��F:�廞�ݙBw=R�Y^�!ֵ�iֵ�k��W3�3�lcD�\ �Ȗ̦��y,�i��@j�����04�e%U��IY���f�m�\�u�[rq����n�WP�z�&_���C��Tv6�kgg�Q��P��	gdu�n͸JN�6{]�������A����s�H�F';q�#w0 ɵ�FY��c1)5J��a���f�ƴ٬Ԯ��l,\��r�7�kyZ�o6o}���
�*/H#�������_v(�x�x.��QQ��߬��y̹���y���/��.ۊ�qG�Lﷳ�D����Cݽq`G�����6��%Ed������G�{��.B�D�\H��L�8���r����J�*'�ѽr��;[�����-H_q��'o���[X�AW<��R�����3Ρ���+������޶s|P�$�x��0'�	>�w��|��Cza�rهה��T���-ݔ��f�?o��	;��|�_t�����m{��82;���I�0>Nx\�oS,�����F�?~��힞���K*�-q.+2:¬��m���g��t��x���8+�ۓ��糲���-�|��!�;
�D����,x���f�tmm�(�����	�Cb-;�`���8��U�^�/@�t�zλ�ܵ. %
L������I��!fD���'�>�d�����@���@Z����%X���p��a �s�������$;y�Xg�-ʩ�7�;�'��7��k0�Za
5Ԫ����*��b[���<�9kN.{�\Xv�'��WJ�f&�*��5�sϢk���}r��+Wj��;�
�f�mM�R+�>���q`gL7s�Dt�]3C�����>b�2T��Ub�T�T�?�L�7��,׵�$��Ӝ��9�QR`�&�
�UxL}l��P��S.<-�a�T��H ����`��	�]4Ħk����KK������Ts�=�ޚ%T%Qsu��eB&bP�S  &����/L���E�9�v��c������=�˨��w^�gh@��������T�W���o�&�۷`tdOj]�jb9�;P��I'.��.�q6�QE6��!!���K3.,d�w��	5o'h���O7����	�$����%Z����ӝɋΝ�0ZW\���wc� ��Rc��­��`c�n�=�Ӯ{�<�9ksa�'�K�������-R���{�Ł�:�����(���d��ԣJ̻7aI"�K�}{�2r	�)2����B(�v�ŻǪ�WNKjݳws��V-7�O6�]⦲�k?;�uXE���-f홺�5ek!D�J=��s�l��@{v��?D~Ȉ�Z��ａﾏ��S�Y�X�ȪSq���6}���?*�!������A+�&��S�$#�����
D�g$̶#��:��޶O�ݾ�@ F���D��e��Q5*���u*f���o0�ѻ��mC��w�ÿn���A�m�̴�G�H�l�`�كB#c��톚���hh���&X���n
�(�ܰ�����'��_b;�ϓN$ٖS�H�%���<m��4;vv��5��\Y)omq`k������G�kg����ߘ��Pb���r5L�~缬P� ?us��L�K:�VA��[�RSiH��L��{�\�A��7|}��?@�x{2O��=�4�9���]BcR�Åf@� �x�K�Kݰ]�G�?j�;�M��AU5!WWu*l��Vk�VI��ǂ�L��`�MB���h�������;$�ޛ�����d��P�,$x���@P����?8��2cS��8�O�w���p��su�`C����۵ч.R��3V���TTZ�����L�
Y�ںH�������ѩ���2[ǎ`2C3	?yw['}�������VX&���H��L�rE�BW9J�=�P���'Z�����!9��9?w��~u̶յ���G�%�ι�N�tż�;g����g�3����ģʺCR&��v;V��*��8���U��;�ŕ��M�5��m��wlyi��t�fi�M�	���6��ej�mu�@�ePt*��w~�d��Ϲ��Z��2XP��~[�쒝��6 )A��\G�����{;�'������s�z�Ŕ�� �]�a���@'V_�g���Ԋ��G���_}�\��ݯ��?D~ɀ����GȘ�K*����J�0�L��l�w!�w���{�����-�@�Q
�D%A% O[��=��D���$��?/���=�,pQ0��$ˎI��sô�o0����\���P��J]�eۅ�d��ٽ��y��b(��Kn
�15�����#RF�^�N�2~��A>�M6O�=��J&�b�����$QC.z|{-AK+�gْ�.�i7 D�+4��{ܘ�Y��w�����ʘ��������l�ٻ)u�����cla�6j�]	WOp��>W��mJQ�����h}�M�k��}���v��ڇh3�N���0�7�\�TU+*�ԩ�Q`gL>�[�6���$<�n���n%Uʒb��z�zi\q��5�s��fR��r��Ň��U0MZ��a)�JKC���=����\X��O��9ܟ|ĜEMe�%VU(��<�n����J�H�RR�(CM��Z��h�h�[�������=�y'7��b���lT�/;5�ڥ�d��d3bn�=��,�ӭy��A���ãx���g�2 ǃ	�z��_��(Dy����zx�����_u�W�g�sUߏ�Y�wI&3j]�QXrH����$8�s�λ�j�Dw��iA	I�ܘ��;"��I�z��;��m��o{	�-k�p���	%wD+�l��
����ġW�%4[���X�[�˒���v�4�Kv�����;�;�9��U��g'�����
��0�i����Gr�~^=��ｷ؉���
�H��߬u��t/q0���Kyq�Y��{����{f��V����5P(�u7���H^����A�qd�mA���b�B�
�^��Xqx��&o���#�<:#�*�]�IqD\���������� ;[��	C�*R�y	Q�?,��g��m������R�x�`ː܂bQ"$�Q��T�2("%~����&7r�wr�OUL�w�D~�s����g�Ƈ�k�4q	TT� {�os�Ɛ{jx��w=�~[���-��0E!����t��B�#��~����:�;��ل����2�&�%J≹n�,^�uT���	>��Ni��j�Pc����0^�}��������;[�ϫ>۝���t�[�i�Bv9;@T�R����^�9���sWe`x�����B�u���nGa7nm�F'Wmz8��v�L�*=��s�Я �Ō/;��dt;:OLM�j�6��b��tY��-�Ʃ���<�����v՛a��HxS��߭��k%��.Ib�d�%�N����'�����I�qā��GT,ԃ,�Yr7&e�?�_��H'��� ���m��d�� ������j՛���uګ0/{�F ��� �y'��q��vlX�+$���u�}�A�����]<s�=�L?�M�Ue��"�9�ŀg��������\l���T.2
���vT2H���7���o:��W�O��\;F��}B*eW쩻E������}k2r�W�S�1���6؛b�I;q�(*j�]�wł��{��϶���r�d ����p
+ܸ�:��Asg�9u�j�ٹ|��5��֧k��f�M60/fg�7 �0��;�'p�$9�$^��	;�W|t�ucR���h[�|.�pW�T��(!��T��?<�yJ��(6�C�б߆���B`��9��í_�����"�Qb�u��� ^��3�ζ���ŝPý��֩��Q��t�d^,LT�Uڮ�,V�5ALTcUT��Sό���;a}�*K��;LS^���;m���i; ��]�2� �{i��@˱`Ì]*;�;[:͎�T7!�Iqmj����@�m5�u3`�3ia���N2c�����-:䆂hVb�ڶ��� �ې��mZ��P���p���L�:Ӷ��n���G�n1���o:^]���v�e���P�pd���g,3�@ m��+4*l��U���'=���6x�\hyIUb�`\ղx���8�J�]���1#��s��muۅN8�A�kT��dc��P}T�-��\na�=�����u�炂k����C^	��ٝ�2�����5U�Y��]�.X�v���K�t%�vw���0L�v��6����{���bԳ���?g��Ul'-��m�f�!l�X����O��=�w�X��޽��Ns���{kX����T�PL��*��)�������t��y!�F�N���T���U�pV`f�\<A������v�a��զ�m��i�l��wf}팳R}�h9{�n�	t�����xu(���w�BZ��ݨ�@{�Wb;�Dq@]�aX�Kl�$��$��������xmXǳ��-�І�&�Y���O}���i-�l�p�n&R��������O�		jE���
֍ј}��������]6�Z7���1l���y�B\�-�iXr;D�����E �(E���VC��������DDG�xڞj�����3�u�ގ�7ԂRbmK��a'����R>�m���m�$��7����
PKn�WtB�>Z����O����R�\Շ�x�\�eA��P
ԍG��~��m�{��q�$��i���s)!j$i�"�D�l�V}���&w���'�c�����aNڸ��P8�R�E-��B4q�"vI߶wc'��w!�-������7����H(�.�)AU���9�k닀��rJo[�Ç ꨘ�WV)�⠋ޘ�.y��}�G�ށ�"C�(��E@�@�J*9�	�J��uu���㾹9�Á�ªY1��^@}�G�<�|`�����<;G����'����ܴn̂Hn?w�v2o�'h��L&6��h�vK����5cĮ%��|����i~�=�����~[����*�Ҹ΂3uØ�]j�`�n�1h��{v���jZa�D}��
%a�;D��l_� �7Sw!��O�V�<��/|}/�U*�U�fEjC�O姿[?-�u��TP����+뒮|�>w'll���IUuwW�PUQ`}����X��uŇW���!?O����l$]0����6���^�&�Ѻ���魓8��u�H��#�@,ز�a�#q�;���v��#TG�i[	�iI��&�lekg���Y� *��n*kN�奫XK�d��n�u�^�v��iV���P�Xne�H
�_��Pf���-ǹ&�e���)Z�����q`LU���RR�H0�ج��;���ヷ*J3ކ�@��uȗy���j%R�q�����b�6�J��j@��D�tA�0��=�\Xϭ��p����~qRbUiM�5S��}.��߫�C{�/�=��'x�TMH����VM�UR���6� k��~K�c�{c�������cjV\�ǊY)��<;A����V~��?D/��d����d�"�nH�eȯ���ݲ\���[�u0���X���q
b�-�Q�C�%����N{��x�-{���z�5rB��x/�]w�Tk��T vayI��퓾�v��t}{�{���49�vݩ,V����oQ(�ʾm�V����3=�f򝗤�tV����5egBR��9lH�Be�*��0�I�0-�[-
�P�`�cK��ߟi����`�\<A��qa�~�<�0�]�څ3bE����A�t�:{��w����o��R��D�[ŗ��QD�	i�����OA	n�u�~����ʪ�	�f-\U��{{�,;z�۷؋���8�>�:5�f�3�'xI=�o��bDd� �pJ%΃���eɡ\^�
sl{��CS�6����ӷ�!TW�Uj߳��vR�9���ny*���@�[��c��G����3����t7ԂRcrcO-I3	��8�l�tF�%cA�A'��1Fk0�4�D��h��kF&�$:R�
`,�B3G!�0L� �����(KP�1i��Ւ�j,�$�#��Ȇ-,�+����I� ���C�W0d(o�B���9��Y$�˶�?o���~9�������	]�
���C۵i��[��c�ɚ���F
�*�U9xB[���}����L�^�*�V��#c�P��X�E��WA��o$?/��c���w-&��cqF;� 9Q���߿�?��~d޶O��h�Çs� �s�0n�0Z���l�%���:R��m����X�L���$>m�؎������j�M!TTg��X��6Gm7�J��N����.&�q^f�7�w�>�W�y�~�\5���������P�*����m���;��6N#����r�\jِI.�P>��O���l��1�l�+�k�~x%�"�c�S/0$������M��(�Q��V�O*p��mF˸�)��>Vn�u�{��IԹ
a:J>>#����2H�6��ֈaܕqS+ ��L�<�����~�ߢ#��o�Wņ�_?�\ԡTd�F^U�TfZ�ۄ��n�9w'h3���,�t��U\��\U��������j�%ӵŁ�uqaކ�5)!V<���3�u�,s܇/wM�|�G�2�H86�[��t�f@�ږI�6@�f4�݌��ȸ�-[`D�R[�lW�R�5p�V�)M�cqN٫r�h�9��wE�s�i�wH�YTc"��Z�x�Y�V��8��ln�S<m�9�ʆnҗ5�a� P@
�_n����w ѐ�qKHݓ�JΛ�	6.g�!(�Hrsʼ	�v�H ��xܪ����mv�<����V����8���I�<\L��yNU���&L�MT��$�Y`F�s���,y��g~>������ӱ$��Ď����k�;A�<Հ�zف�ᦩB���.�1W�`{��`n�2�{�:�)���������e�W2MR��oT7r�n��h��w�ـ4��Ѿ�ˣW$,Lw��c6�'W���cQܴit��5`���N�^���&R���b0ۆw�o~�N���dｽ������>����Ѕ-Vu2�G ��3��i7\�8�ƭ�P�?1pVu�t�H�k[�?�zKtɊ�B�{���SS�[.��ؠR�SS��ݦ�Β��`c.�p�'!HI�d �D�J	�& �:�C��Ł��f%�-�l��G(�r(�L+�0���v�3g�h5{zKBO���Q���$d�-�V$&8��w��I�}����}�vc1}��%������g�����U��7rw�`����ô|w�A
	JK1٠R��I�wc%��Ki��J�W6u�X�X&DAi�\�Å}���G��&���h��%&}%���A#jYQ2$B�
�����}��~��1�rj����Nh��QW���vNk��*��X5T ��[�`>�o{��65�T���ʩU8�0}P���y>I7L�=�7m���#�b@�.�I
�mo�����,	�뇈ų��a�p�ML���갊���{��

��� Q�P�ݛ]�#�v�.{M)"�3�k��3�\���y#��mG��t��ԍ�T���x��� *d�AUZl�+ԃ�W\�n��w;�`�	q5S�7�a5�Rf-��o�y�_��}�mW�g舏�hwC�	�2DYv$P�'�l��?y��H +���@r5�f�A@����|-�⩘�NY�AJb ���լ�k&k5.�֌Gp���pC\�ѥ�8kI���J�l������3�#�7 r��0F�$b�(c�NQ	HA9I�d#�y%�98�Y���c�^h�:8�� �Zt��;�~S���M��]s�]C�1���5%*�a%�����"m�q]-��ed�Wv՟������T⧙7l�A�؃p��kZֵ�րc�1���1����1�1�`c:0��0
�ֲ���qm�:��Zִcʦ1�c35"�5�XOm���v\q;]�(�n�a�vD�N�N������&��0 ����.Jh�/6q�ۗ��i�(��-f�bhI���5��"]���?�7b3�*��Ѩ�R#"͋,(a/L"�wn9�Lv��l]��u�V����T;�ˍ�ĝ"z�O�mf�p���vXՉv�gP�J橈��bT`���)�`bִ��Pӭm�Wd}l��d�_�-���������z�')��	r\���t)�(�m��Aۅ�)%�:�ecL��h] ��Fmj.�
�C%���R7R�ۃm+���^]<Վ9#�2��{u��Y֙�$�ە��[<,�!�j+t�@t�*c5���Pz�\F��g��i`�Om�/m	&�gZ�kpY6�9�XlM�j�e�8��Aؽ:�G�B8�*1��P���n̆�Tf��]1`�:��'(%�@�[	�iXp-M�Lv�[ͅ2�4��aӷ��.�:ٺ�]f b�t�6�ZՖ���㟈�� �";T�KR�b�ښSw����I1���v��G�>6y؊w�$sJ�⁯��b�)ؠ���" b�
p}��*�����I�W���xy�I�e�����f��bɋ7o����
����K�����UM�v�߶i�O8����)FJ"��H�m��&Фg�����ަ�m/9c�ty6�\ԡA���� �vΌA4�1�a$��	HM)������=H��\�C���؉���߲�X�̖Դ,Iwa��y��X�{��WY��,3a�P�L%Ys8f*W�ɍ܇��Vf�W�ݲwޝ���y��EwvD-ؒ�X�]�r�.���`d��K&��;`�O&N�Y�z�X]s�Hp��|n7`����!�6{u�*<,F]��w�:&6G �mnPX	��a��c 3���흠 �1[(���u��GC3PiGX�9��	��Ij�ѹ�m�����;?�#��t8:0�įӕ9U3x�oײ��<���m�Gh#l����B���h�
d"e�����>\w��>��VN���2��� �\1 e/�4]�m��pv�7���X��J[>�֍�ކ�)	�n��/0����� )#�t��<����i��;P�T���V+�I�����q`��g$���Hwu2�����㸘be�0f���O����}b��s`�{��7�&RUmK �e�h��wfr�мl�)�vg�mq;�9��k���s��EUR^��܇n�u�;{��x����sg[����� �� �5 ��>w�<>>�QŲ����ye��R��a����+6J�X�-���;����8)��<�dߧ�����A����V��H�B)H�ĳJե.���T,�a�ߟ�qˀN�䗒��Rj�p>u�o����� ��o�q��#%�NY�N�;��6I�lhky��y�w'�lrqSJg&� ����f ���;Λ�q�-�E�%gSj��QP���H���{�M�|��~t���뎴gF�iA��n�̎8~��}�l�eZ�ĐQķ.�ۧ��<�mn2�R�v�v =��`�{ێ^Q��K����{۶�G`�[UL �q����T�(�J=2ڰ5x�{���?P U��˿~���r�0bO1���'��:�W���PUB���� �\�C۵h��(ޥ

�nҕ(�&��m7��P�f��K�`j�t�vÆ攐*���Qu�)Y���.n~���,��A�ky��s���DR�7R�.	�~���D���D�M +���Z�DΛX���񩨩�T���y�yv�C�k�O�9��N�<�t���ζ�)H������N�6�i��ź��>��Y>>�Z�a9fK��
	�On�y�~��A������;vz��^�;�_�2L�"I�IŘ	=��D����}o� P����9n�K{���$�|��˳d�pI1��@
���I�z���i���ߣ�-���l:��\ԡTe����ُ0�ۯ����a4�#k��㎝`�|�Q�g�؉��*g�����-Wŀ����%�Jݞ���N{��);}uTȱ����-�N"�������>^;��O��>����؃��;C��|�L����0���Y��ۛ�>����]����a;��8K�5v��Rp�l��cv�:�zl�v��+'kNw'�ơ�	�.&�nԥ������Gփ��Hy6��~����ceG�34�b6ZXM6��OO�f���:rv7�vD`+�m^ۗpm=���-�.��u.��S���p�n���]��4��N�v�`����V�u�u9C$�s�5���ѳ�����D�����\U.��v�n�8�R�ݲ]�$p\'��ofn�ZM�#eSJD'X j�!I]�^a��@T������w)/-;�Olr�rJEPe���ބc<���N��1w���wH9p��3���A��ŁO�|�${P�-
)R�XZ�T���ŀn���}�n�C�;��.�?}*��j�Y7��3�f&}��y�y�jӝ�f�5a�=2�QW*�.b��&��䆮��� �}����
��F�@�fݽb�!%�
8I�dz\/[i��e:V��	�9۱ג���������Z�~4_{�vwN���%�i��m�I�}��~_w�y�ePkiD[���ӽf�Z�r�����[�p�V�k�׊�����?��o�]��2RC��_��6�鍙	'$R^]�����e�$�����_Pnε`f�򰁾��f/>;���>��"K#�0�a`�H���
�k��([������F�U5eH\̗I]������rj�.�?k�VNh��� Js$xB�75Tf�s��� ����>޷�ָ&���n�AM"���ꎴ�y�����:*���f��%R�R�SB�T'�}���<�5i�l�to6bh��!@^*��m�(�F8�iD	�.F���	�^�O���$53��v�\^�Β���"
���MZ�K$��o���UV��B�+���,���:�K纶��;�n��.l���J�V���Kf7�B'v�}�=^�K��۳. ��>��� ����~��Z�>~�9�.!MbO1�2'/	>]˭	�a�֌��7��ȁ��Fg۰z��{�[��M7s`bәri���d���V���el�)ͫW$�'�.n��R^@�s��9܆���k�k�ln�k�1̍�<���'�O���y��,[��-om��Gh��_Uۑ	"�ib�޶O��k�� �C�
 ۝}�a'��z��]��
bj2��̫���>K��Vާ�H}��,��UA{�|l���k�K�EeGN��O݌��|>���4�i�b2�)u�رe��dBX�D}����ţw!�ڎ�g����RF��:��Y۠E���1j�*T���� �����2���oV�l��w��p�ڒ �(��I��,[��v�y!�y��	t0��>���cYX�Y��z։�������7����n�kwo���{\.��"F�H䪂������!��|X�W�~������M�\ݧ���6�TI^�'+n�n��1�mPfz7g��Q�mvgj��1�v�-��vٝWf��[J�
�G��f���|?)򽜘��r���63m��F����z�EѸ�R,���.�"���������a�QE*�2�r�
�	�'<�w����,��i�$��BWq�v�)l��Z��W��~~X�j:�i��x�֎R�(�Jһ%��clc����MT́��ŀg�u�?ky�{]2�O6��M
�V9��u{L���\����c'��z�9�ܯ�/pZ��iK�Ც)EZ�n����Y��������[��i����0�l4°�a'��:�>����r����~����}�I��
�T��(�6v��9�;��%��2���z5�ݣ��n���]�A��M.���o�����۫xB\�`�}��-2,�]����H�֭]f�����݆hKaf	��"���5���D�#{�#���i"�
 �:���12�r�	F��뙲5R���! ��J:5�Rd�S���CDl�lŭ�m$0Ki�6������Ж�w�ł 2J4��,��F{��!AD�����%�t����� [����:���%��t�s�؎��D��+Op��o��!�	�ł	dX!7�rY��40�O��Y��uX�nL �V�*�TA�ב�=��$&I��Uz��A���A{l�ָ���Si�z):�vp�����X��j��j�
۵@�WQbP�1�գjj�,R���m��Yk� L�qC	f՚鎹�B���Z�����^�1�#k
F��/t�(1@֦v+cF7T3�m�ڬ�8�*���l\�]�j0�݉�C.���,B։�[��qv�M��p��Э!�ak�����%	y�eR��
'�ݝ��'�u;g>NA.;tٳژ�\:�s!�JV��*��6q�R8}vF�;�UYi��m���y4�z�uv����n�)��ʣ��<�o;��]�n��R����X:����\�@�hf.�]hG�Ƽ!�nU�]��=d$CX�M��C�I&���9�8������r��� �Q�:�w����K~?�H�Ϸ�R����)���\�Lb�>N�WJu����9���+��d!Q�T���X7[jsk(�9�2���K��1�W����� 
�B�O-a!�$D���K�S�Q?ݩ5N�=��`�Z'>cv����
��Գ-�Q�����H���f�5`{�Q��#jw��B�����o��MTf�}�X���9!yw\�����<�Â�TUڪ�T��A�����{i��;W;�ۣy�b3Mbk�$��8�'����y|�Z+R�p�Y�;"���B�Q4���O����P۫ݻb��)k��&2�R�1�A%��\*L�C��ը�X'=���$-t�=1�rJ[��rwC�:(�Te�";��	'|��(�'5��d�ޚl��v�g𪪦�Ws�����7l�� ��ŀw����OT��y!��e�״�O�0��cI��~���]����y������T?�N7�:�����IR�.(�>��>�ZБ�^�Q���1�v-�TM��]�	�o�O� ���/;�%8
��/��睗��f1.4,6���cJ�MTҟx�WŁ���=��r{��	����w&Áȭ��q���n�e���b�˴y��Z���A�\���fX�N��։�zwc�}R�b���1��:E_:��}�n�`��=�J&W"&�ɔU�ʥW!����z�܃�����l|��)�IV]�����כ��/������H�	ɉ�����"�$R&#O;ۣ�N�ym�{�M�gۼ���j���X� �*'j�n��<�sm����}����]�!��� v��C��嬅R�&q����Ď��y y�v�{z����N�I"�UB���D�`?>��5�C��l����vI�a˚���%M$)�
�����n��`}��C�ڎ�-	� �Y�r��[ސŖȤ��.�,���q͝�mZ��s���6�8�z��a�\�q�sq�t�}��.��4�yd�:mc�ޕ��9mٴl��=�s�����Ӈ^�)W7�Zf#�QZ�u�mj&�j���;�y�9$�Y8��?~�G��2�VT�R�[��>�m�ԉ�?�)��"B16L���ێq5��J���!����偯�� �u��ͧsUQ5
�^Fao�'�ɥ�X��j��7�ђg�>���!�=�(�����r{�y�h8җ%�eA�����a'��z�k޸�<��6�5�T�*0��˱TM�`y��XA�Or��А�7r�_}��r-�
2ҖS�
Y �X�['=�h1�<�9h�Ɍށ8SR)�71��xI�?o<$�!����q$�m�omQ�a��C�S���AP�����o;���yXx�����]�` !������h�e��.��s�0������7e"��K�b�3��_ʅ�SC��O	ԣ^�zn�l��Ij�1�Y絳�,���5&�v��н�m������ �)(�@�Yr5��'�7��w���>�7�UP��]��N��2���;�*@��%��(�g0��Ǻ�P����ޱd�/o;%�����{��c���f�UU���Z�~��`��}2���Iios�'wF�f�TMck�%w��b'7[���6EO����-��AP[wj�ME%�?��ل��>�����,6���\�kL5���4bB��L��_�>��k��i>�V��qٔg���Ν���-�R�Ÿ��*dQ5T)����N�7:Ձ�ꎴZ��f���^�}[lFM�ҲO}����(
�Wf-Ŗ�ｽ�I�z�{���R�"���+%M�=�V������"?~���U�����Ït.���&��V��~�A�ms�[�l~���9���G�C\
Rc�;08Y�,�O�i���K�ame�t0��EYDۆ��a)\Kmg�}�~�m=��`Q��o"H�@t�#�SV�ʤ]x�k(�fn�9�k����f�2��uGZn�䖺w��w�m[b�*ɒ+s�����}"/�{0���9�'���;��E���%�Ķ�o7������u���>Ϲ��afH%
��%H�(w(���y���{�Q֏{��Ԥ)�ʩ�KȸK0�9���oWŁ�ڎ�<����q�MA�8է!���D�1�O�(c��ȶ���e mF�,�����J��(AI������y!��]h�q<5��+y`H�1��YmPP3,��a&D��$�q�Nn�<��?����e�M�%8U	EY5H���M+A�sy�_�"T������CW��l���>��#9�C@ZE<��$��N�g:�hm6�*f=��H��TQYP�n�9p���b�9������;���j�o�+p�E��m=�Ӻ
�yX]s�I�c2G�9=��ɓ��w-���Om�W��Z�v�G���)`3"��Qڸᡅ�.�ᮭdN���l@�5�0nؐ�V�t˚���6�,s۝:�g��e��F�و�n`e�Z E������wW$�(�x��`��a6��{�P�/c*C:�-�	]��Ye��
j�R�~��R��m��w���Q֏=����n�w�x�y��ڋId�1U1"� �)Q�{����n�=��œ}�h��G.�& Ʀc��wUx��,�ݘ޹���J[�o���E��&\wm���s�Z'��k���]��w�ů�z��>�y���BE\������`��2�ޑ�l�wځQ�r�X��h�vym��0źF�Lj74�[���ғBc�~}?Ož��Z)v�w<'�h�T�'0;��z�|%�h���!������}��g���XKB;���S�!�M�r��]t\t�r���}�]���(í��>&)�Q#%���e6b�^��k�:hG)fu����n�M1�\�}�#7`�c$|����Nޝ���t,[�b�d�o�)�^����n�Ł�ڎ�{M䛨0����\�H*"���k���5Y'~�va'�oX�� U%��ߘpR��%R*p������o[Ž2��A��Ň�Kg��*.n�*�M��y!�,v��:�h��7��j�$�[�X2�'3	�w�Y&��D�5��[��M�ݪK�#��S3	J����ں�cm��:b��-ۮ���y����K���VU~��UA�uE~ݸ�k���1�=�_!8�*q^d�d�����Y���
^P |y���O��Œ}����x=�7M�e\(�%�����<;_G}T���	{��X{������.L���f���l���U�����mo�}���Ds���FH�Nk��]�A F1$��Z��oio �KN�=���n����`�ôy�%�.�U79c�<��,�x��E�u��W�y�7���&7r��V�J&W"&��HU�ʥW!��o>�o���c�J^�q֌ޏ�U2�5Y5V"؁f}�OZ�v�q�� �H�hb�^�u���u�31�$
��RO�h%Әؑ���#��J@NJh�N��K��ID��(�)�	u��JM A�#C� Ⱬ�4%	.�r R�$D
;��dN0�F`ŌL CRP�A	D�����E2H�e�!T����c��p�Xe�F`�l5+� �&	Xf�i(�l�%�!,�K$�цY1��!���X��(K4$�pS 虀��BP�%#�R�2
�� É�������'@2JB�!�(JZA���R���i!��pp�����>�������1�k���1��` 6���͠���^�)����Pb3:g4h��q�n�ct�^��t\[�b+���$�Yֵ�G&0 �1�h�1�b�g&1�[�c cbc�c����D��cŭf]�kZ�s!�c�^�ܤ�X2�t]�����֭���mu:Z��j��S6ݭe�g�Fё;ӗuV�V�Ê�ֹ�*�M3�N��<<0��K���(���6�1YP�+�ͫi�Q�������^��#����/m�p`�@�'U���r��<%�8{$f�a4�Z�;����l�v��v�K�k�`UE*�v=q�&p�:��]kp�EYٷcu%U��q#M��fH9��� �G�u��˹6���2v�Z��u�[[�#طU>m�� =<��X]�n��b�*6t� ;Erd�F��m��Y^�n�u�l�]�׆��Z�
�6��M��ۘH�F&,�s;-�kX0�1��a�E�Yƪ��Ǟ�3t��ֵ��i�0��`\06 k\e.�&ǯ]ێuf�-�`M�c[Z�V�t���ޮ-��"����{Q�_�w7q<�"�x��j���Q"5�[�+����s�����/X�NzF�9֥�e\���m[b���J�L6mCL|���윋y9�>PGZW�Cν qSj��6�zw��W�H����u���]�XR~v�H�CJ�U�~���ʊ�2N^��V@j�t���C����8�4.��5�����	�z�d����,�����@}��ɨ%~$R�"T5T�6��<Յ#�{��o�>��YM�8�8�-Ma�"��P�$QJ8�,�$��ݘI�x�['��'Wۮ�����7��o�Y0=�L����=��)=���F��_���r�r�VI�zi�;�:גs�<�<��ɚ�KIE�)�����
���������䇻���H��1���fvx�f�Cs!%%��.٣l���Jw,"�i�i:�%����#�4سM6���O"�3�����kWNz�US��p#E��u������&��Ģ�ܘ�Tu�p��a�h߸��	<Ģ�:( 8 t �{����[AƔ���*��O�v�b&��x	L�������n��غ)K^�<a�i���Ų�������{�R��7H��F�\��F�"P �	D��Ae��,ih��{�
_���������I뿾���mT���sJf`����S�tl�u�{�M�t�+�B�]���\ɑ�n�xI�:��=��0�2��_�����(�*H��j]ۅ��N�s�O�g$���VO�߽c����ÑR���7�e��[�yY&��%�Cv�rI#1���+F�5�Y�F������ �uq`=��u�"��^�~ECR "�P���h)���h�.�;ì�5�q�+Zc�Ϊ�
;w��,F�
�BX={����vSJ~����sG�\t�d�&jU. %jz��M��#v���mX�o�{�<�f"���c�F��T2��`=uh5n���M�'}����{y�	pe�i��,���ڰ=�y!�<;BM�Ȱ�\�AQswV!J�UVݦ�Cɷ6j[��1k���>��̹I��pXr3 ��e�1������V�z�gR��"f�*��AQu �A�N���v���������z���GP�(Dđ@�O��)�ok�Hj����W�����o�'wL�Q(fd�ٍH[��=�؉����$�q�(P�N��߭��p|�n��ʳo8l�����߿���@�( /�s��_�!�߮,	���=�O�ASY7Y�QH��f�r������y$�WZ�o0<hB蔜Z���`���}1����V{k�I��x\��+�A��R�N7�'��:�.J�*�QVbE��8�e��	Mjj`"�dou�Hyo9���v�����K�^��wu����R+��H��	(�`��3*����� �����L{����u�;�<�D�N<��#p`G05i��7[��3���#^�y8�8i@�f7�B@��6m����I����N�aVRe$� �"a��)$������� ߽��?f`m�X8�qМ!N�d�)�'0�]?}rA����5i���?DG����+�D��
YSWUD�i���ɵ�w��.��.���#n�&f� Pdi����D�_}��̟w�X�I�y�ᯥ8`��W3�+��@l[��v���Ǿۿ��ylƻ�����s�0#Z�	�5R�f�W3QUvg���$y�5`w�_}����Ku?�>��R�ꨄ��#%�s���w[�䛧q`{���;жzeD��])��T�5W'�����9p��缬���>����Gq� ���/��<.mV���NV�hՍ�����ǲn�(��&�uZ�B�=���n��م��y�T�����ϣmz���᛬J꦳����u5���;$3�sҧ]�ǗmD���.Ҳ4�m�M�"UT*������'��5q��53���3	���l�1-a�����	�bf6�m�H"�%A2�{{z4\o\���x��܎L�����j*Ae�h�THMH�
���7]GZ-7�B�{���L������D�k!EM��fަ_�26�������k��Dw�'Y�wv�"ؐ;�_����7y�a��-�Qv�[�ôw������+$s0�ª�
^{ߝ�^��;�Wh#~�o$�AߜQQiZ
]v�w�G����"ĕ
T�2R*gl�w.�U��1��q���������o=�q`���M�2ns#�#�A��v�V�n����md��i}T�{e+4�%��w��v\]��i�+Y�h��1X.p�r�Nn:jo�����6��@�X�Id8�[,P��Jj�ͨ��]1s��9X���v-����h3���3Ӽ� ͘�rw��AQwSE��"���׭� o&�C=��z}��%�>L��	LeL⸜��f����3�\Y{<WT�v�ݵ݌�{X#���q�bvXJ��P�_�C��ޘv�~��R�Mܛ���N(�k�)��f/ ռ��Ap��W�a��6�j��ֳv.*��
�E �~zې��q`F{���:~�FZi����$']-��fr�,���JT�Q1J�����M���޶No��G>� ��6�K�L0��s 5���~��������`r��a>����|t��6�I�`�`��$��L�#��u����[�l3�W?�t*��B��$��}���~���}q����f kMܔ��Xwq(�����LT��Q%d�}�{?���l�RC�� I�n`6	��5��6x��g�n>�?u� ��]h��1�S
f���~7���ަ�d8W���fl�7f�q�h5�<���J�UJ�6�~�eL�����`yx޹��>뇈q���p�8�qc�]�xI;���9�7���
@�UU�
���~���d�_v�'�0�@¨�sP)�"jm��x�#���R[�:�����l����%�ݶJ��e��ߺ~�kvgb
����u	qc�r�ƃkB�/��?~���V���I�50KU373e��ͭF'�r��Cn`LǾ�CS�lݨ�A�z�ޒ��������dx#�h@�8�_?�dﷻ0���:�%��wg��Z���̒�*f�M�;y�9p��k�́��6���#�����m�0��oK$�lh�^>�f ����&��(K# 4@��(6m����Po!�Im�,CEDD&69�Ib�;@�"0�� �3E�]d[�f������f�46� ������rK,��ӵ�[M\���B���Y�p2mF�*:&9�+vhԽ�)Dnx��Jks�ƒ��v��εs��ےvm�6��L�6V*�F� aSh�\�rHn�.gs���8\;��U�3�"6�m��I@b���LO���{�sq��2�ݧl$��Ϙ�M��d�-H2ed��9��6�j�U@�hX�:`{��X���Nls�H�4�$ݔ���!l%�4mnHPH�jU@� {��0����۽,��z�G�F�,���E�#7a�|�>���DBC�Q����}���u[� K�h�?"T��1����&a:����5o9��^���׽o㣐K�TZ���S�2���}�e���w!���a?��o_�d�����pb��ư7nf}��-� �U
��i��m6�I�J�@,#l$�J5�?��zI�������>>D���/���/�`~��0@U���*��7�?ݬQ�o������GZ�b�b���B#J��x�Q��*A�T" S{�QF�4,(kX(�G7���RJ��Qဠ�AV (
!�s�D)D�
�@ &Z�U�DM,�(��H�! ���b ��D�TA�A&@�)�0�GEH� (A] �(!B�(Ҁ� �� ��ߊ#�#�!AH�(A�0�*B
P�Jb�
r@M# �B"4�|���>���k��AU(Q����DG�'��_������O���������g�����	�����3�/������߿��h��O���Oe��__���9�?������������� U_����������_���Q@Eb)���C����~������/�S����E�����������p��������������������_������?��d������|�C?��V�Q�������������v
�P�
%*%**% �J��J�	��) D�HD!�)!K�,� �@�2�! �
�!*��J�0�HH��B+(B)!*�!$
��	
0$"�B	"H	!
	!2
�$"���!"��(��(H��*�$
� ��*���!$��!,�
�*�	@J+	BBJ,��R @�! �H	�	��
H(H�(���*��
��A! 
$$2"#!0��� �@#@)H!"B0�(B���	(H�$�	)(J��BHA �H������� �!����@$!HB�!(�R!	@H	 J0�$�	$�P�!HD%	(� R,@�J4�0,���!�C
	��! ��!�"B�eHV�F`Z�F%�aE�%XJ��	B��AH
B�� �(	�`@�Q�Q�F!V�d��(IB$F�$DUhPp�:���W���u�S�TAU�A/��H��5�z�W����~���p_���������?�������$ Wa�?f�����������߯�������?��� v~����F7��~� W����P*0���?�����~����{��� @W_� U�����&�N�AWO�O���0b�
����;��S	���}�ѲL$T�?��������k��p  ������������~��y�H *���������p����~��?����3��P�k�@Us���?�9��� U\�=QG�'����'�:���>�'����sxG�2�'�ߴ�����G����q�s��~�<����i<#��� U_� ����~��~��������V�)J�t��3�9�������#��TUy�A���?��"(��k�������AWQ��������������������z�o��?�����)���j ��o�9,����������08_ }@� T��&p           �|π]�Z@{�(B�7`h 2 �.���� � �g@�   Uw]�]5���x{�
� u� ���ҹC���݃@;�h����A@42�K�:(rC����Z�z��w��րe��Pwn�����
���T�p���Z�9��+���J � ( U?�R�A� �  �  ������&��d 220�Ob�T
h i�@ �@  ��5R��    @�(�� �1�B'�SM4z�6�m�B��%P!�i���hт4 ��n��t�M`�DB��Iϯ�@Cq���*�"��PO�8�>_⪂1L;���������(k���&��8Ω1���{c-P{��}�_i[Am����1+�m�*��mO��[gO�M�U2� ��U� �h��L��t���蒖΍��RU-����[w_*��t������1�wE=&�AE���v6*�&�iOdͰ�/�)2L yB�!�d������a�ik��a�4ȔC�ĉu��R�[��;��v�{�SBX�9˾ن�f��;SAa�l�����]�2�N-�	�9�`���P`L�۠cZܛ3��	�ë.1ը�!El7"CA�b��(�1# �U6���F��.6&��v3���ӗpq�@�(�X 4u����1'(�H�uf�g}�;wsA0N��
Ŵ18���y<.�=��qРH6�XNm�Q��,'���͘�Q�r��^n^lг[���s�42���bk���4���Z#zxt��ۦÌ�p�����F��,-9�4��de�83�P�*@�)$�h�#ѭ�fg����o��������OS}y��{�H"`�a�Ù�6���vXA1��""0�A���ߴ��,b�!����1aQAd-[�U��Q	�kc:�ߖ�;������Ȓ�����dN���lѤ5a(�
�!���H]�!W�n����㳇�6Hkf�-�:}^Q��k�fbJ�0�3PT"I"��B.�ذc�d���fͶk`�l6Fq�`N��h��3A���UC��O8'���VQS�L��{�Ք^Ř�i�j)�� 8m`c���0䤴aH�* S LP<q4��:.�]`ӵ���Fi٤�4��Fh�iᠥ�&kZcf��&:vZ���FC:�'C���MH`�#	D�iCU!���.+( x_��h��ז=������id`���4�P�5�Z/1�� p0�����,^0�:�����M�8��H�1M�y��o;�G�7xs�ֿ��k�X�EI�x��$"�4�+A[�����U*(+ �~n��<�ì3ÿ��H8f��6g|�5V�V������J�ň&�PjA[�`Hr_g��G�s ٢<�7.I�ᦺ �"�I�Y�B᰿������ t:�C���t:�C���t:�mImԒ		���t:�C���t:�C���t:�C���t:�C���t:�d���[D���t:�C���t:�C���t:��`���v� �:� �EɱR�[��vK^<P%2$��V�(n���@�vI�qs��W�[.(�E����"%�-I! t>���	'7ܧ(��v^vI�C���C���tL$�(���·|��|�$�D�C���t:�C���t~���|����t:�C���t:�C���vKh�Kh�:�C���t:�C���t:�C���t:�C���t:�C���t:�md�����t:�C���t:���C���t:;��{�?��o��w� ݑZ���ؗ�kwU%hln>�8{�D��S��N���{��l<^�s�9���[�S���F��C���j�"J'X]����g��ӹC
C�[d���C���I5�TxR����4�6D������Jұk$�U.[z�ICJ�R�P$��H��@{�̮;�WT\{��{���.�nIg8c:��Ű�ay�H�=���9`M��jj����x^ٻr�=�p�W���I<��jtI�*%�t�nak{�SD����9����7~��$��,�oZ��+�7wJ4Vv(V��Q[�����d�A�Hq#����Uyzl~������wf���|�ӆ��=J����Ude��|]���1x%锒��lI���n[D���	+�*�
4�S��z�����;�bއO,�{���}[a�0�f��0�6��$>|Gq�*C%���Ż��/ ��+W�Th��oW)vL� Pt��Մ�(�&O(b'��n�z���z�Y���'Q!;/
v��A����\�O��hDR�f֮�J!�Ѽ�t��.�@9B=�h'�T�^%įfb�|`P�^{���-��
 �O���2��>$�`̏MS	ш���{�������ZV%ݣ)��ے��xƭ�����t:|�a��t7L�!�ݘ ��w0::�e�i����C��dP$�C$�k���$>��C���y��t_媃D�ΎI��[H*�C��l���`�v��s	���t:$2#o���ќ����G��F)�C���+|�t:�C��0�E�I��k�O7ʅ���vA$�@�t:�C����j��Ht:��$��$�C���t:�C���3out[j�!"��CS[pQ�v�Tzi���\��jG���Kh�Kj@Iv�͆����w����U$�.g0�QS=����#�*�*�uR�fd��@�i �p:�C��������t:��$�m@��0P�8� &�C��Ԓ�ѻ��ܒ	C���t:�,$��RH�Qht:ш"��aC��yШ�^l2U���h�TOhT�^cר5���ws��c��ܖ�-�!�PV�ܛ\Gs�a�_�o�����E��0I$����m�|.���{k$=� 笔�F�^��"��Jo?��b���olm?.^��:O\�r�8s &/����~���;�L��tE�o�}���Յ^ >���Mwz�qAC����(�`�j�K�R@t�\er}-�B�I6�s	='(4��͆wB�o�����y̒$�C���cñC�d�|�t:�d�����P8�C��Qht:2$Im��<�����s�4����9Шh -�l���t"��0��v��|9��n�sIG�9�lPH�!�@���䄉@�w% u�|u���wr��⤯�w���>x|��#�����`�Z�̇�$��Gv�s�{qV��e;���$un�ww6߯��DIZ�̧|L�B�j�%�_j����>�/h�9�k	t:�܇���T_"���HV����k���/d�?}{�lYĒeaD������qx:̿��r�~�!��\9���~����l9��= �ʭB���5P��XA�(v7T�/Z.:DDA�LF��"�S�}G�����b����6+�/H�JqQ��*b=�� t���@�Q	�|P�(J��	�N�{DM
�A�OB	!	�"W�S�AN�$��QzB�ڡ��$��� �N�}G�Gh�@`��&)���C�1K�~_��rrs��B@ӡ~GUF��2�J�V�ê�j������[M<3�1z�w/��î��煘��M�F6^t�%{f���h8�csf�&U]��wWC�w���6�q̽�yղ'�AH(���ph]Ƃ& 	=��y�#�Te���;W���di��IwT�Y�m�'�;�}��� ��3d݊�)}�ݽ�W}�5��^9|��.<�JTP��+ݓ۳m�$�Q@�dۊ��O7����f}��o6����"ۙ�}#'��9���UF�+�tX7a(�X!#͛-	~��ݻ]���6�Vn?4�_�+}s����
���ԤLy��@��Ԑ�m���vba零m��6���9��b-��'-��۽��2�S�Y�"�yw'ZlX-�
g;�v.J#!4L��}�XGvo������L�����跉$Z�m���&궎�st&�$ʳx2�5�wZϩ7u��B�,'�O�p���#i�$n5&�����פQ��=�x�(0Irn��2�K���� Mx׈Y�}n͇ZD5����򒴋 n��_����Zk��&�H�
�T#HƷT4�&˄$�jkH�W�޹�Ɩ'J��@4d�<�o�^�7�i�5���o�$=pi15���t�3P�z`��W�3ZBw]�"�BE���4����|�HFj�7Ѷ�.��hi�#�5�P��֐0��e�ZGw&�i�Rj]#Y�n�D��!��B n�d+1{�����H��sf%Y�CZE�P[,���s��;��7����V����^��c|����$�U9�.�bX�nB�����Tߐ�Ff�ZAÿ�A2�m�%�մ4��se�	���\@X���-�₈f���Ցw�®�5�iZ��&��B����C��1J�Z���a�e"~�0����Z�)�!r4X����r��tk��.2��3��jkHU��C��4՚�Yhe�"��a���Hq5d[^�hf���V�*S��W�"8�����ģ����5���R%ZM
Y��,���!�H�i�4�{�0��F����끡�๾��I��!5U��C$���i�ku"�m��u��CMi�UT{��qC[�!T����Py=�62!|zqc4���\,�1�8�XYh�tlH�$hN0�٢bѽk��}q�Ѕn:��.�W31;j���H��6a�N��v~o�s�"؈���".�E���[��6:� DDDD���g��̸h�7���e�3���BEP�e-�7Z6L��`���I�)�r��I96���L-yxM4���u�2{�:Y�1Ǝ8��ŭQ���4��t�%����$A�|>|�N{u��GBu��:��^x�a�0W̅Y6��dU��Ѧ�R3b�s)�Ҳx'�� �H�>������E�\��pi�F��y��D�u�|���'0B�KphiN[�f��i�I�51?�
�����"C|�5�Y�v�/5����'7�i�k5����H>���ݑ�j#�\�r���ԇPt����fė,�-��l6[�3��q$>C���iˈ��5�1�H**ICu5���~�J��iF�%�|�bI֐�����߾�#�\j5^#F�E}��?
��>%/�2�$ c�m"�^�l:������E�!@�C}uӲ���a`�cp����A�IՔ߇Ƭ�Ʋ���I�,������ i��VE��Q�Y���#MOs{&;k�(Wt16>-�#eD��y�O�?��a�ٯ�[�Zn}rC���bkO�x;�!�{�C^5d!w�끪�0� KU�PB4��c��Lc����ݶ�VJ)U��ҵZF��.Bj���f�@�}s�n��X@(1�^����W�@Q���CV~��� i���4
�F{����E�a���U�,һe��V4��[hx�	_A����0�[@V���D��q7�bܶ��-�V��ςkvj��*svx�z��1YJ*��_|�Ȁ�	F&���iy���-[i�ÃMa@���]����F�P�gE8�q~ �8=��kH�>!�}���/%�@R^�!�W��ĝ��)�m�����L�[�XGkqR4��9��w�ڎ�$���C��9.�i��hx��w�%�Cijw���i�kMm�鄳�bF���|#ET�/�(��̹����i15���tf�U��P��kC3��U�a@�����!��^�E���˺�^%.|1))t�#H���xд�0/�9{��]�E^"��̞�w����F��y��Ȍe?�:w�a
��v�i��4Ր����n���S�K��h��G<B#ƕ�,鎊؉�H�i�5����J���F�+�sD�4��5�[]�B��xu=Ɲ�����\�ލ�(���;�`���q�������ŬkOf�R��ģ��GG.�+�U��K̿��"��@�Cu-��0L#�F�P�gE8�qV�d l�`f���֐��'�4Ր4����>�D<G�^���ͼ	8Ʌ�'�4<F�ӎ���9�l&;}G���c�ǂd� ݖ�q���5�b,Ӭ�p8�`�fP��Λ5�:�7���f�x�N�(�F�\i/K�4C�����/�����$T�t�)p5��UPUU5W�N����e���!zܽ�v+V�p-M��B��k<v'f82�ͨ�:�X��s6V$	v�Wv6� �8$��92�7;�	)JR��V���WF�t���J��0���
B����
����#i)jF��`�u�|��u���?������l�~�5v��x���	F=�0֑f��5����ù�w�P���R���.o��l�����"�C%(<�P����Ps޶rN\������<��(�/�8h�ޛz���?>bj��`�%'�d%:��ͮ�i��ͼ����MBP�����L��#� 4s������5	Jy�?Jz��`�0E5�f&�p��Ò'3(JB���5)E�}|��sZCR�I��'V%'~`�B��1J^��ɚ��\N�(H���JM���J��(JN��J}�b�;�"�44���P$W����*5��u�|��(;�!(Ol$(�r4=���%��@(y*�d({�%)���JPu�&�)���9����(JOa�
݂P�����J��(u|���é5&BP�a�P��]��	���a�Os�(wJQ����/6sBR�^��J�!���I���k��mr�o�!K��"�Z���Xo|}��
Y�R��A�J:���<�E�XZ�|��I�����);��R%�)��ߚ7'����r��0J�{��%	�`�%'rd%=o_>\^o7!������J��)�R$���<�B�뿟{��ԝu��
�d2�$)<�%�y�r$��g�Pjʵu�cP�ێ�7���g\��������+iqj�nv����';D}��%=w���.�kzB������ϟs�e���ff��1JB��H����H�}�Iݲ�a�s�p:��/,������+����L��Fu�̯~lM�Py�&�(N쐡)<�$(O3)J]s��9&�s_3a�JC��)J��J��B���ܚ������^�ԁI�	B]X%	I瘚��z���>]�Ru&BP�fR�����4|��e���w�'R��3�)<�!)�z�Ϟ�Qŀ��\�R�\5��!���i0ħiڔI(�t"�47�MBP�܆BRy 	B]fHP����.s�R'��!I�2R������MBS�;��_9�hP�>I�$u�d}D�$��JR�@wϝl䜹�]l9	H^�%	I�x���<����2�t|���3�b�w�j��lϚ���7����ǻ�
�P�	��.�v^yé9k�����6�nJR�&JPw&BP���BRw��)���|]p�iMHRy&A�*Hd�3)
���5	Bu�'�$S ;�ލÚ��\�(H���JM��� �2��J��J~}1u�]k�С)=�R'3�)<�%( ����޶�s��!(O,��(�k�˛�Y�v����_�u!BF�L�����(��;�qr�s��,���7	I�	B[�J��0P�'Y�P������ԙ	By�/�RD2R���5	B{d�	I�9!N���x�.p�5	I����R�f!O@�.I�9!BZ�J]w�{9&���}�rR��/�|�	JPy&BP�,$(JOodԅ7۽-�����$(|�%(4y��f�֬���Є{/$2R���� �C�@��48��t[���$��u	B^X%	I��h�{���~�|��WP�^5��,߿jWv��a�O9�>�}�5�g�K����+�*b�	�u뷬][1�WV�Mu�"�n@�e⇬��3��g�յ2��VY��{<�����O�.�b�\��>����@�1Ol��*��ѫu�l��{�<�ʝ��ϭ�<j�E�� ������ʬ���N쏨Uy1t�2.�{�w��n�	8Im���kH�ǰZx��@�U(	�r  
U�#5��^ȞU-�{����|��|�N�ގ4��jL%��#O�(�5�*�����|�W�^!�XB��)}@�F���t�gq���Y���=�凘D�d/��՚�Uc7I�B��W	�7~a��՟:����Cb�fN��c05�j����/��������F��>��7�B?U �4�}�烗�@W*�^#�U�3��E��>���A�R,G��Vi��x��o�ڳVmقcH���(�!�!�/F�x��6)���{�W�߆�	9�Z��k5�0Ѯ�/{�l�]�t
t�A"��sJ��c��r7����$'���|�V��kZ�kZ��au<�۰��psP�yU""#h�����".ݎ�cԛؗ�:{a�]�Nq���X�l�8�v��d����a�9�[R���q�:�c2����X�º�.g(\���kvV��$A�kC�@"�c��O;s��*ثE�Q����^��۝̝en�3��k³a+B�ˑ�J��/>zn�CluJR����l5C$ ��"X]�����>����/z��}�P����'���e����#�R(�A��G�ݏZQ��l~���CM{� =UL9��x����ZjZ�P?%�ZM���,�}x���<D�<C��˷��t�slx�1������|��ا�q�[��Mk��+�I�IBt���߽���q�a�`)��+>#H�ҿlbOSTǨU��V@�j�ؠ�i�(�5�U��wdi��>5�c]�F=�0֑�p�{w^ �|��X@�e�"r0��P+l��L�m�F�g% ��M�!��O�P�vF0�y"��$�\�?UU���;����a�ϟs[O=�S���>Y���>
��IP=���=w�ë�i�_�=�G ?B�W�|�ޗA��NI`i�i��������[����B9G�(;����Ƽ�P5�{ϿdP6=���M�'ߘy�������3��)8���K�?�P��k��qV�2ZF@��B�
�ЧZD�o��E�4�1xuT}����q�k�!����p| >5v��a��Ҋ�P+R�6m6�3𯶡�����*��X4�&5��_�ϊ�In�C f�g��ߢ�Q�6����T�5�N3��Ϥ�k�-���rb*�UGք�0g�ԅ���6��&�r$�4j��yq̶`��+�-�HfI��3^��(I`�F"F���}@:ӓ�<F�-jϪ�Ȼ�
h{�a��/�z˱�U�! _��a#�ik>M��N�j4�_��C���	.���Z�4���]�AMHCn6a�J(�W�^*� +�����������5=�/ ODe��,��kg��y�~s���T>�0R�0��C�U
�?d��%x���[�9�F�}BP����{g���fY�����qߊ>��
JF�翟u�����"��]�Ͽz��kOs���}T? J5��>�l���눏��iTp�F~�6bC|����CMє�sr���^dQ�)���� ���E���`I_�i�U@�k|����םo��w�]�2��X`	  
F�	�"��x"�#H��y5���}�whi��d�P��)$_����{�{�{mD���7�A�!��D#�^5k� �qQ��#�Y�/����ʪ��HA�~v�9$.)��e�11l�M-Y�gP�5���J2��v���{���Uv7T������O�6�D8с�W���^��~�'v��+!AcH	������5|5��yv4�>> _��l��p���{�e��ϭ@<G�������*����0�x�����@i!��� J�	�"D�K!JD�wu�v[���ۓ2��u�U�J�4U%��L+3��*6�v��F�m^84����W;��ۊ\�\���*�gmh*��f��Ja�fSF��r�C�����s���QT�G
L��@mU�U�T�F�
C��~L4�M6˔�jr������l�������Lfq_Zhx�4�k�����`����Y������<k�}�Aj��j"���� ��XkH�ׯ-m_Qr��Y m�_����J��HJL`�QX�c����/�������~\���5���VB#���U��5����ȣ\�iR�|A0�gƑ�jp%�:X�$6�i�����^[���C���;U�fD7Pȇ¨�IPE)���{>y�����U}�c��z����4�F���&��B�,'~4��'��І���<@Q>#Hd�l:�B#Ma
�s���U�x�x���kH������SqYmH�ۢ�\ܣ�p�70.�\�l�us��$�M	w�������vkƽ��n"�pbJN�2*�3Tw F�1�Y�\U�8���w���k؇e�7�����9��ٰ<E�|FY֡��5Pt���y���;wN��<�x`�&�H��W�u\l�(ڄ�Ur��A��%4�-�
�?��
��Մ�&��8����cAj�B����<@���x�������#Ma�o�%���u��4#lƛ0@�a;�3od$ �cr 23P�C�ώ��|����P�0��y�w�a�xCdi
�lQ�Po�a��@^��H8{����� ��[Cǌ�6���-����!�U�a�n�_P 5W��߾®Z|F���<E��}���*��Y�y� ���{�~�����&��e"y�0�C'-`��0���ji�!^}�X��U�x�7�a��1j�B��3�ٯ����'*�.l��\=7%V��:Q�iKc6���֠b4�0��$Yp�&�P�� Se0�+٤CCV��[ �����ZEf���EIi��:ns�6Պ��ViwZ��B�4���C�H.o�b:e3�+5T��H�Ti'�)����A��z�3�hy�#���10J
"4��Cm�d���"b|G�_�v�5��о���nƝ#��K�'%i�}�����Q �3���:�H���Iq:E�����Y�j� P����"P��5VW�	aܧ� |Eo��!;��z�خ#��I`(NC��#L�m���!FJ�A�#M��ʹhf��*Z�s^�{��;zt�3�PR�JӐP�f`"�ףG8;"h�GA�F �T��Z�b���(��(�A���Zuђw=�3����"""" ��Ɯq��<�[v����1���5�7aK�/��&y��WV�6�]���Ayp�m3bÙ��@�!]�9㙸�㗎�t��U#���"�u� :5Hk�1���j݋���9\�Q\5�Q1-��˭Acf�̛D%r[F�^�ː�v�6dM�La��-�d�8
�T.�U�PmQ m�T}W�ꊟ�����{�j�!�5�j��M@�@�7�L�7��A�:��4�EKUv;��VjйݩݑQ��H�<z�,�4�Y��#�l	3gp�#��.6����峻1����5�]NEZ�$@ 
��]� �U�)�iD�A^�7Nl��aՆ�M\dx��!���m�"��׺�a�Y�4�"_��M:F�R�N�j�H�UP�7��!Ÿ�$CO��d��UN���>}\��DZ�d:4�>td�SPB۰(\�YL[v)�=�ZC�_j�Px�M�7�-��U�T�%�Gq�"�Pç��j��w!�4�e)�!�V��ٮ�pʉ�Y�\U�P
��ؔ+�4� <P�P	��ݯ��ZEf����$�#�}l&��
_|�`(@������{�U�q6��� xT�/>O�ۈx��Bb^}O`�� 
�T�G��rV�l�4�E9X��>��@ɐ�M�X��Sp�_U

ܦ��5�+�B͛��|�Ȩ�äY?	l��A�ZhZ�C�a�4�������х��)<�{E����q�h���;E�@�����FR.�U(W�!�zD�#H�����P@U���/-27RTE�Mإÿ��Cƾ�2"�o��di�}�`��XEMU}��!�VjٿfH�AZO�>���ނ�W�֮�	7#���bXv����؉��I�"�h^��V���ܷc��T�%�Gq�"�P�C��j����hi�B#���
�5�Da�K۴�/aS[tU�L1��U�U��#ό}T 5@*���b9��pQhf��<_[	���6F�}�U�CuQI.e��(����V��������i��:z�:�Q���XB<{\�þ��� XvB�@��܂���,n��*b��<��#}�n���PmI`ZCN���e�6#MB�H�j�#Ǆ�Mf�� �U�C}'��a�4��C�����i��C��I��������Pxڌ:Y��Y�\�l�e�uj1�Z"�U{t9��{v+	�����[Q��A�GƳn�q�����2�i�D�?\�ZE]���jQHi���.��'�S�7Ui���V��Ĉ�J,6k�����:ֻ�G���V��3Q�	ca``B��	JB��uۼUUA[���+U�UAUTx�9��iZ��nQ�0�g��n6��65���D���R��X��tG]�t�AFѴ0��TlhR�D��s�2n�M��'l]u�����w�t UW�B��P3<�LQ��RDc�Q���'e���K[���F»e�����a5	}���"�Pç����äY����f�qV�א����HD��2-���Y�X@�)��FT�"�P�B{��w��x��F`�҉����G#�i��A�#M�u�r��U�U��>M�����V`*	$��.���{����i�PU�7Ua�#�:�F��r\�y�����w~*h!�A�Y;��)h���!�����"��ǚaJ�DK%{la�4�:%��	��f��V������(�*��p��&�hxU *���2rg�b�C4ﳽ��wٹ��:���f��}u������B���V\H�$Sa��������B�&�]�L#5lsmpb:)(��3@��v�j�$��������9�R�"�P���d�t��ZC���up�#�(��o�v�o�pO�.2%J�z�v���J$[e&Q	H�,E"7�V���G�����l6���Y�a��|u\T�f���Y[�G��گ�!��`äa1U�.|]i��p)M$�iv��m�E�H�敛������PM kj��UY��,)Q���$P�*�Vr��}iI��.Y������
�Z�I�x��ٜ�雔��l8�q��{f삼�6�������5@�D 
��n�}�Uzf�;>�����H$�!���mn0��e��77�P�g��[�y}h|�^��o�w��{�7X�fq�N�u:��:,�X�k�%,j��BYt�<�eO��Nrr@�Y����s�!C\�T�ւN����4>l���mι���ɑk�3f��}�&�ùs�!H��Y۽���͝-���K�L��қ*2!M��"T1�(���ٱ�t8�k"��;ɆN��ͽXM���h~xǏ�)�[!ީُm�
l�!n�ݗ�iI��P�UB�����ݙ�w��n�u��>����$�~��4�V�t��ͽ�W~�":�e� ����<↨`P*�	�M�@�A����+F�%������f�"� �a�T �v��R�QEQE���2͞���e[ޙH��"""#h����*.,ɋi�G�v��4�/Q��a�n�f=F�=ms��Ǚi�`ƺ��4���81%8�i��b�E�v��nl;U��H�:��"�vЙ����G��	���� �A�op�knOi+Q���uq�5�Nh�2�b�F���S :�&��{�ћ��>�v����T���<U� ;�|�G9��s{qw=mf�{�D��b�+�n�x�g��� �|�F�\rl�H����,f��1�d'N(�2����nP�k�mn��k2�m!�9MD�d�Y��1�����B��Rw��/S�A9&��ە���{�^f#��� &g�ϛ�������}I��
(�^�Z;{�ܑ���,�x�.�;G0[������]UP��?�0dċ�U��gy���㛶�	��{*5��N�	��p\M6�h8���76҉@�K���B���3���B���{6�_ȥ�fپu��{f삼�7H�)q��	�<w���p�bN�Iy�o��߅P���߅�9�mUU��=m}@W���W��:3���&�ŶB�(�����-�A��"���~�UB��/����nw���nl�.��cow�NqQ�'�I���x��͹�N���Meu͞4�l�v��I�ˋ�������q�*��0��n<�z=���Y�L�E���L6�wt2��g^�ɛj�~�sN���M�	M��_��� �F8�L��IB�P) �V��fqu��P��X���9�n��{���s�~�l�R�pRf�>�� i"�f���-4����e�4��
4*���7��y0Y:wٳje����n5v��ѹ�E-���oc%:��Z�n{:ͳ��n.穭�ʪUP�A_��׋Vo�U{��}�{9���UA
Gv>�sa��D1";�6͛��nl�.��co�޼Ο`s�3}hto�#L��Qƣ�D��qgnd�nݔ����[L�����k��؛�W�����E/�"M@��3P1�)% L�ɵwpe6b�f������F}�3}�
��w�F/x}��3!�X1;��vP��L��I5�SP�c�[4�&$sF�R��^.�$!0A(T���f`�B�4^g4��kFhf��5�#��Z��PUSQ�Ί-�2�
��j�6輅wC��x�:�j�6��Vs�/�y�]���%3���F�dq�m���n�#����C�>xYW�Ɩ�k-[0���d�>� >���;�򮦋��g-9jKP9���99���wV�u���{<�hyͩ�=�l�A��КaNW��I��B�,.3}�oA0���ͳ�HS�\��U@c�?���5K�ͻc�|��qہ&�"2��Y��l�)�K5^�]�B{����������VN�w�{�����ߜ�!��y>0 [ ȣ+y�t�	T	XƘ[�m�w�l4������w��}w�}}��➹��Jg<S����mr���n��Txa�.�M�`ꪷ,ۓ7Ǘ1Fъ"�yٹ��*��n��;0�6L�VZ�#�y�C�{w�^��j)}�ѧ�8��p�م��s��r\�n
#p�m�ͷee���j�NMSw�UC{�7��?>�L�i��L*������ߢಬ�Qo��HZ�M:a���nEh/��uCh Nڗ�n�� ����~���7|y��c��HJ+5�,݉)D� �=�ٽ�5�z�fߢ�jf��P�@����Rٛf���G7�T(&���H@�>�3XE� ��͚�/�&�ͻ蹻�owݚmɛz�����E$,�R2���� ���+��Qlk��$-6�D�2K� ��d��z�"�3ݛ��2�3
I�L���w)��]Ѻ�`����u��}#}�#|� �[���䞠$�W� �i��Ĭ"蘒(�(�(Q%E�
j-�O\W�P��(r�S
�V���ڳ=����R�q�N�j��@����)�΃.�~�������Dn�%4et=��o�AO7܏6�	Q5]3��є�l���B�ۿE�$�3n��RܿS�0�B��(�� 찈�L���341*�3��6$	,D"R$b�9 �E!f�5$���#"J�`rptw�Y��q�DDf�rۭ2��x[��BDV�a�ؠ1�z��	��m�T��\co<\v�-b٬(B��Qf��g�+UpE�$� �Z�������a�Q���ڹZ��N�n��r�V�;l6�-d����q͟��z��[g1�Q��8e�ѲFzj1rVv�1��5F3R#L׿9*�@�"U@\�.�].�$���8=ѝ�۴ ����Ă�'�pE�n��Вd�fI�f��\�添���ݽ˝��E���r<�TUf�������i�aX�I���i,��ٶ�2p��(S g[�����9ƃ�X�ُM��W�-U�v`�?y�a��7�:<}����pf#u�L�����.Xl��[��J�T �#I|g�������qd���q1H6Sm0�f�����fm���_c	lY��	
vk��Z	{����@�pFSi�_j���N��Ey�P��c�>O� P��-���7nm�}Ч��7�t�p����J��o��%DA�=S6��>Rܽ�fǺ3����B�!%�$� ��b���^w0��o�@fN��I�'�e�b�F��F��{὘77���7/�:9���`k)�K{�ƶ��N�� ��D�=V�7k=���9K��ý��۩��y��5B�j%v��x��	&�){���jF�"E�6Z��K�f��9|���]�\_U 7�=�_�i:���Ci_��[�ܳ��Aq���6�2��fT�r&�`J4�}3�����S�R��n����3ê`44�{��U
��{�fg�7{�'m
jM35��!`��*sw-�Zsw�
��Ч��6�����(W�������G�O�ڔ���ޏײ7��m��o73tٱ�@�se�/��6�
 R�f>��&��y}]����((�U�e+��=��;�����e	O05�Ê��=3vͲ����oP@*4��4��E�I1.�,6kN�m�#��D�}s�",T�ױB���5�uv�O ]F��h)�`E�.Zq,���i��P2Û7V!�3�F
{3w}	�忨U
�.#�{�|3�$����n���V�S@Z4Z
4 ���8ޗ�8q��}B{�~�eUUQ��jTT�f��!�}����ӫ�\�6�<��Q�Вӓ�D^��g9�P�X!��
 :%U�LdP0�QD��riJ��[�^�[�f��ɲ��*x:#(7�Q�A�W�߃������A�9���1���w��2�e�2�F�9���N?U�r����k�Z ����IՋR�������I��m�X���G� 0�`*�>$���=������E�{���E^��>�2����@��V $71�����&�&���l �C`��9~}][o�k�t��e�vtp��PB5���J�TNq�l@A'c����/P�n�}:%�w��Rz�_�����`b�`_j��kZ�ۀ�[�o.��L6��zW)Y�Vwc��ê�I�8G���TPCP*�D
��*,*
�
�J�B�(����B�**)
�	�*B� ȨJ�B
�)
�!�
��B�(��t ��(�RX�2M�.t�S������p��߲�*�(��D �]�&0���l2���:I�`��-�<�����@�o����b��8y����<�:�����u\!�vDUEPBA%���P�T&ڇ�c��u��ߥJϮ����q�,$�D�H�_�Y]�cU�=����;�y����a�W��ޞz�6��H��\��PC��1 ��L�u��X�~%�>��v�]ӄo4wv$ā��,�
!/ A�I��E�|�Y�X;��LµO�#%� 3=�/�!UPB�`��i���P���>�=Q����-c��a�s�E���^��E�ٳyT�{���0�l�a�Ey�C�~�SYk�%J�������dV�~�w�Y��B�GM�O9��!��n< >�w�-G��ƭ{� j3(�������~���$���e���PΟOk,dn;����xx�����l#A\� ��dp��
����V���5��lԁ��
ȝG^p`�����!@�}�yE�}[7���a�Q��a��ǟ ��0��n����b��{�`��[����D���[��Y&��뵴���t[�g��"+�ѧ>L��
��c�8��wT� ƛ ��A1P�tW�wm2�b\uF񌌡��LA����*tX�*�'�\qӫ�h=@�����T�V�b8G_~�?��ߖT�GIͼ:�ޤ<x���|�[؃{��w��yuP�-�A��=D \;��3?���)��q��