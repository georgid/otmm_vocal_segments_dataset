BZh91AY&SY���o�b_�pp��b� ����a��� �      ( �                    0� V�   >P@�   (  @    P  @ P(@( �   R�    	 ��           z    P     �C 6P<�2q;����gG������(zw��ϳ�`�|�At��G����{4qZ���A�4$� ���&�����F���IM
Q�(��@ h0h�S��R�+�V�k��     h� ��
be>��GQj�ۥxm��*� 4sԬgȹh嫋T�6��U��( ��K�t�f��S�44 ׋T�[�T�}���J�k���}����ҝk�J�{}� �JŞ�.m\�y�.6�eR��'�V(��x   ���;�(:>�T�}���S֮}���YB>���(}#>��38ڸ���ͪW7� ]�xU�q��{p����i� ��-+�\ƕ�}��{�Uͯ��G��W��ͩr���O9� w�S-{j]�t�3�J��6�}����@��    @ fM|�e�f��W,se'[�Hq� �V{>��+�ۧ���UŮa��� ���+����|�� 9�ɥ�''R�}�(:9�V���]��۫�/����n��� V��R�q�.M:�Ŕ�˕O�<� ��� 
:�� 
�� }�K-�����l������ p���YK�N�۫̓��eJ���.�,�8�J��(���u^������ ��V���S��&�59���jW< =JŒ��6���W����O        ���MM���   C@ �?%*T M    '�UR�D�      Ob�QM�)@     ��5d�T��&�    �	U�@&ԁz'��Q�O�=4��'���?�Կ������vw��{}�"� B��@ T �   �  �(  O�ԡP  ��`� ���V
  �+�ӥ�$��+'�j7������&��:�e�RsDf�"vV�j��M��_@���A�w�����>e�����Ҏ �AT̎
�w_����n|�Z<\��Bi=�9�c#0a%�H	���
r��tH�U��,xb�#�~�|~0H��:�%|���I�9�yiC���9�O>Y�&�^&B���^A,�����~��i?�${4�=����ɣHo&'>z����=D��G�t̼`f�xh?O�͜؅��2CU�Q'R>o�{�<�G���V����y��!�`�T�Ύ��e�wn�R@�71���ͭ��3�;��O�>�<�i?�y[1�����v��!�f=A�l]8��'�B-�k÷u"}^��Ǧe�:/�7�,̃�z1 `�!�^|e_'�㔟�xp&%�t>"�e��'E=�����ʳFj��z6�W��XJ.!�Lsf�k2�z��{8�h*�c��_S�ȋ�š kxP[��P7r	��? ��}�Y�s���^)x��nr�����z�)�lx�6��&M��um���b�;��ᆺ� �L��0�:���f��(�+W%��>�HߗW�=�<j�Ey5��I�&�	���M	�f�2NY�Ɩs)�'g]%��h3�{&v�|'RB��!NXIrD��sE��n�˳:�+�����c�������Q��>eoֻ|��w��$0A����-�4��ʛ}��`��ڰ�1���B ��ϐ'�B�S�t�L�Dә����|I�9��b�RW�:_�[���R:,hns�x�d�J��tA�����Ji-H�8
42�A��Doc��`�d'.»��Bf,uû��_!7t�3��2k;�m�sh�¾�oS���B�(�H����=�WhAq��es�Ӽ3����	�y#�>� Ρ��:�{�������6}�	���K&�ټ����ox�̰/{e��k��R˛�}���9���F�3����Ӛ���ɥO�`��g��kz��؄��_ P��A���)��̇*�bx^��8#��=�=9�����A�	 %<q�"��%���7ACb
͢P��W�!�,F�O���v/=�{�'�Q� t�J+~*��_r	��!�M��S0˩�Z�:����+�_V��A�z�ɐZon-q��b��I�Jy����X\كՓ�j��sC�)�Z8!޳�5�`��M{{��X,����1xmy��.!fg����ꨫ��h�%L�ga�d@�&վ���b�N���Ε�b�[�����?u`�G^�һ�{�=�#�8!�1K�gwRX���Է�|��Ќ'��<�ߊ��	K�&��E��K���k-ϷFd�gT�K����.���#O��7;��8z���(�ϝdh���ߌfv7�p��
l$��C��0��:{Б;>+�^'#��6���8h�8����ZS�DnA�*�#!
H6Qq���F"Ra��V��,L�>)#��8Q:�3��>3�R�Z"=Ś���>b�y_�7�r�{���	}l�`*k-d��w��ӛ���0�����9���7�b����L9&�v	W_PJ_BR���<AݣS>[%��0{2�؏��p��giܬ����3��)I4���
-�&8j��/Mǘ�9W�Y�!��t�H�:I`��wQ
	���^f%#'�K�H�vB=����(f9����p��`��~a���9at ~%��|��8���D�h>kڜ~����~D��A�s3�L�U�z��4��E�:�<Pb{=��L�5w����Tb �"SG��5�)N��/�4 ��6��?/�#͓Fh$���)�'h�^�B�rn��pa��'�!H����~�%��Bm����qޢ�D�����xfq����b���$�)!�:}4?�� ��L�b���zG^ �Bm�ب�{���~����ff�K��~k2�HH�5�C;���%���zсu�37��w��V�kٰ����n����y�=p��7��8�ɋR5܈�÷��Y�s���cˁ/<>��������n���c����;��4�{�]磙��7>T���Qݚ��7�;lz�"Vёx��VN�p�X�
���3F��>Ϸ��3���SpI�A*	�&`��H$�H' ��j	�& ��H&���0I����f	�$�r)pLA3�I�$�\0L�$��	PJ�\L�5��n}�7u�	�RsB�M�9��c!�����;�>#M�����������,�x���Y�7!OYu'Sq��ڦkŦ��B�LPn��l`;����}�s*͞ߗʪ�a
��?�?(=�i���(�"H4Va���?O�����w|n�c�����*����ox'�z�q}��0�;�sQ����n��5�TY������_�W-�+��LT�̂��#j[n-��d�dZ���Q���~�����\�=�x,z�p����P���S�����`� ���.�/�ׂ���+$���r��'1B8�7��p_fٻ�CN��߷�M�L:�c���2�fEF;�S�`j�� IKl7��M�3���':����[0ng�$6�x��QZᅼB��<AY/���v�p�=u�;�z�4$�ߣ'Վ�y�7����Gb����x7)[�̗[��ٛ��ۃ��'�4t����H�@����Ӫ��K�w�m򒳼�ճa����s�ҎB[�2�:r}�U�K���^He�]ϱ(rl �#J�NI{��R+�HB�4%��'n3u�a:o4x�����hY;��p�y��w\���ٙ��b������pTK�M��PB�xQ'|u��sW�|�?s�]�!�_���E|��fsX����9,�l�9o���P��)�'�tn_�S����`ܘ/�I�%�9����K�|\
�+6%�`y��;G���pA�>��#�^��e�79��@��'½�J����Q�������3}�.M�ˤ���qm#��ϣ$�c{��w�q��7�H`f���<o�ۅ�?t�����7���WnM�Jfon�*��z_��qI�o�4����G�B#�t��W�as2�	vz.I�?4�NC�sM>��}��|��5�d𞺚��?:6���E}��a�v���v3��{>k�n bɻ�0�^wG���?)I�״�{�U)�F�S/[2i����د�-ɼ{CWgM8&Y�9�T�ٗ-��Ao�5t�70��s�{��MA����5	֣�j�P����Q�-�yz	�J��T�ǵ��{�sܢ�6e�O��-ejR��X�H����>Κ�O��˵�㐪G�>�^?J'n}�
�)�C,$��˱ؗ��J'$[X�TdDl!Jh;�u]��l`���st���>~{��޽x8����%>��g�ǖw���ܬC٤+֍A?�]:�s���a���o-R���|�0p���a�1-y��{陼;�#c�N<� �X�� [��~�{ݘo��}�. �DHecJ��&�؃����^���Ä1$��!����(�E�U�l&��Ǆ �W�|CD�6������b`\�%��(2�)��P�/�5h�"w�\ �K�&�H��'�62��)�(5��~ә��Lvw�G�/�k��Q�}�;�i]�1���|���ǹ%�%��=m@9������p���r��!L��B)ɽ�1F0w,���;�_�>ϐyP3��[�ܾ��A��ˤ�Ť�oS��Z�Z�[�{ėQ`�n]�W�{�7-��q�{f�t������i�a�>�3|7y���/|fJ���~�|�����>"WY�����-xW{z�{��-��i ��o�b�&��`�]���d�7��Ĳ�e:Eq�f������&9o�Lw��ɶpd��^���w,��%\f=�s#}��+&�~�Q����י�k9/��ǽ��p9�1C�� ��2׾�-Q=�%rǚ'�G�o{Vz�ޘ��'��1IM��c^������T����@��P~�=��-��]���C+�?UD�S���2xҠB��=��&O_M{�@v�� S�)80�V#v{+��=�*�Ω��2��?���;���7��]������/<	?@���')r�s~����l���O�߸�Y����=��T)�nt�=�vn0ya�`�:��+A�x��$>�F��R6���0W��������x���Kzv������w���I��w:K�z���Z�S�{��' �v"w�{������F��{�=����޾��v��"w�:��w��s55�q�>'�4��/ge{1�레���<>�ݝ��燸���ዼ���g�8h�A{�{78:���|o���G�N��S�������[AɰL鹨d>:�[��8�n|=�����i[O�^�خ`o>Z�ܚ�����_`$�ͨ{�����9�l{���mS��*�H��&Gg�9�x}J��L���%�Dix!HC����$�=���L��񫳠����M��đ�y/�I���Os&v�6�r#��I�H�(��3�/]����c<=�+���/c=2������(Bi�`&A�L�� � ��s��2�k��v�����j]Ӵ��b�36BM"N��������J�I�:ʱ����:\��rtozy�
���]r�.��Gu7�fݛ�:p�!��A$�X�Ɗ$���׽f���ś#�*�`����t��ڭ�*�3-��ot�a����'bߚ�w�o���!~�O��F(4�q���ښ�$��>�>CD "M�00T��f�������
��`�G%Ȣ1��/^��<JY�\�3.(�X�I�%��Y�p	�\�4����qO��Qo!�`��5u*<��H<w�	����v�{����}�����$�h=�Pϳ%�zMW�i��$9\��P�`���uH���s�$�ԝ�Ì;�Y>!�N�0X,#AA����l��02�G%r���*������Oq1�����eݱ#k0#���@(G�O-c�sk�����})k;~{r���ǨMu��[��x�aG���u�\��ЏA���h���M	��}���S7(�U�cM"րx�`��Be�;:����y=�$y�z}1í�d�ouf��1���>���*�i�Q!���||Wc�׺�3ff�Y�ۿl��"�<ժ�c[�9�z�Bk帠5�o��9|H�޹^	�J=�i*���%7/�O�y�8�ߪWE*��������lzl�%��E��!���������u�Җ�C���R�胞�=�|�k�-�?�B�\po����0�-�L�<oK_s7&�`��/���K�2���I��voG�.�i�������>��?|G���p�=}5�M����BgN�e��a����Do��{�E]�#�d�)��n����?|s�K��-���!5>,��"�a��۰�ziY�wA>9$�y,+L߹nݥQ8�hu<�����k]y2��p��P�.�z�}w���L�F�F��1��{F>����(����/}=����6�ہ��yUe��n}�` (�2Ϫ(B
«(nb��)Q^�Ίa�}/���3Uohk~*��9l��Mn�05����p�:�Ñ�:Aes��)y�B�~�L-&h���ڵ���ΝC��郪���������t��gQCņ;_LQ�׬��4e�jå30��zi)<����ǿh՘���h�0-����h+
a���i�9�M(L�h}D7�j.>��x�0B�nh�������|b׽��SU�}�K�~	g.��f�!���4]����-��Hq�<�ޯ'PrnM���>Y�i���^�f^��wLېi��4y,܈F�*��wW}�����n	 ���L�5���	�& ��H&b��H$�j	�' ��pK�\�M�9�K�H&"���u�")J!��r�7�]�3Z> ���0i^�!�L9��fn�ez1���^��9,�\�\�5|��s�wڙ�C�>�n�v�z7h��Qw���ƻHηG���2y�lgSǵE�wv���%��}��ȉE�x��;���3����5��x3��4� üw^��M�8���
�ѫu�	��4��B�ri�*�0m?A>GT��_�t�e|A70i*���G1�֛s���*�)�`C>Cv+ߌfA>��3
w ���>UF
���y�ow�����;)$�h�����[�W��`?��?<csO5��n|Cp{v���j����������
������w|~!`���hJn}�@{����^�ۓ+����a_;���oE~Һ� �6����L������:7~!=�CH�f�� ����B��3~@��P�#ئ�/A��Ԓg>#���?'.���R`Y����SWR�r��ߎ�%^N�y��^�G&�g5T�b&hr๟�`B~N�u�����)E�p���]�׿��U��uu$�I$�p� 2 R��l ߪ           �            �            A�           8            #���H   !Í�b���k@
P`8 �P )@A����� �pf����<       ְm��gA��  �  �|     `                                  8 ΀ )E�)@A�M�Ѧ��wT!�F� gK����$��cxrkl痍�s��l���L�\�w=Y1cQ��=�'M�u���x�4�̉u�n'b������n�Јn�9,T���l.oY0^��]�����ۑ��s�G&�n:��]�p���k��
F���i��\�Xu����ǌ�
��B��ݢ#�������]�d4���/h{R�mٵ��;��q�֬4�h�E�P�*���*E!(!Ge�����+����L����ۚ���'\�cs�cn��[n����(B{:EdǛnI��1��'��b2i�f�f�aG1�rv�ۖ���s�k��lk�J�n�5֬�\�g�ͯC�NXS�&oIh��F%懫�u��Rxv&_;��$i��)\�\uIn���t�`ۥ�\ijvM/;`�l��1�+�t�\pk����t�]Љ�7�䒹�P.6�N�k�m�Ƹ�ۧ[�ugl{L�vr�[��}�k��'[��)F�P��nv�њ{Y؝�k���x�z�<�瓳���m��[g�Ǣz�tN�[����.;;S��oO�͒��H��6X����XX�y[�-�)v(��z'�u�c�v�d�mm����t�ظ�]b:�4m�aV����sۇ��8�u��c�Ctg4�3�=@����\��|�cr/��Y�
W7S�glbj�붩�s��y�R��cl�=��<��:��sj���Q۶⣈�vMhw�c�������tQ��`�3��Q��������.��8�	톯��Sۄ�0�>���f}yvz;��kЮ��v5��D��\��5�厢��f�^m��$q �.�O ɉ�1�v<m�G\ݎ{�K��v��,ݖ�\B^�,�9=��^ؼ.!�x��	b��Btv�#kWv��N�6����n�/;X�'eգ)·c��^b�sr&ݖOP^���n͊gu��\�zy�M�	<��C�j˧v�q�I��]p�݊7�ݴ��0��f�]/�ٸ���>�h�v����=��fbL1�ű�a��ڲ���Gm��K���V|u�vƦ^t��bM�u�Iͭ��f�aF�Ȟ�zĪ�8�c��sV㞺�@j���މ6�;��{�g��	���-�]c K��s�͢��lqxxM۷5����r[2m�d�kbv�l��ɚj�܀�w��֓4���ݳ�o�O���A� v�7��[8;U6�wXŲ&eT�x�E�;tl��\�����+n���۠��R��	g�m���@U��U�km�h��1��ۆ3�� �.F��rY8H�v'h��:�h1�g[Pml��Lr ��FL`8�]1�9� �O�I���k�kv^0�۝K��c)�<����s<԰A��q;er��%N�:�����ێ�l�8��VƋrB�n7Q6�Շu��.�gb47Q�!9�<����q���HUVƙJ��Ѯ��8[I��bx�ǷK��Z�c��Uo6�yh�k5�=�.��������w���k��۷;�qg�ݽDW[Z�m�<aԉ�,mۮS<�C�n=v2p�uY�V�m:〥��	�P�xy�tvte���]n t��Ʌ�,�u��:���>xK�2���y�kc۶YG��͊x5�]�о8U�&����[r�m�\ۍt�����[�;=�-���7+V�������u�(��л�����v�u��gv:�t�fȖ��6=����#ry�gVd�Vx{s�tv�DQ�����P����#�ЃHN�vm3��ȯ�7G W�] N�kV�V�dۄ���-Oh��]����������<l�\n�CR�)��0�<�q�r���4��۷�� Le��ݘa!����۫]����3tF�PB�v �y��L����s�<FjՑ�<�
wf��/aL�h66�ېvC�k&��N�"���)p�aÇ��(�5��Xڭ׌�9����݉u�m�sm�s����q������{-���q��na���by4��8���n���x�0n��->�����O�N:�W�u��[�U���ȓ%���m�o<(�Źm�n ���ۯ�Oà���ئ@u��ļ&8	�ywom���?���ꃪ�o.^@mJ�U�q���k� 'xݢ���2���7W\UTn4��%���h�lu�c��'F��K�Q�^�ۦ��Wj�8�ib|�z<�t�r���;�랧���;N>Dg��	�����8ͻ6�ٴ]���c:��ia:�a2�T��qM�C�gnb;]�b�ے�L�/4vx�,q<n�U��mЭtVS����v��.c�.�z�{��X���v�+ �®��R�Urm�%�s�&֝��pj�&RG��6&굟)k7X��8�{[9�������p�/bG9n�:��.�d���v�j�$���&�t�6p�����5p�9��h�syx�m���u�&J�ꪸ���.�ƖZ1ƁZ�^T�c2�cVne(7~��ﾪ�<�����'`x� ���n����u����f���<��]��r��]rNX�Q�Gt]9������G6�\cq�jOO1f^[�p�ECb�٣���ڎ$L���K^�a�.�����%��m����I�z��0­����c���Q����Z�����ʻn�z�u��*�vjx��d��+�6��Ih�ˇ���h���m�#j�'e�k�\:@/a	vSvxA��QD�R]",�c��&k�����4�� ���m��k�zP��ѩ�ڠ⠽J��>��������	�j�[U�����j�{*�S]��f��y��D���;pG����ͮMn2��ǰO;��v�f�m�N�;Tj�KU.���E�ƴnR�����Z�/��c�&�m8I��Gm�苵3�m���:��7o7��C�c�N��3��!�[[�[��Sj\CU]C������Uw:w�[����|I���n�h;M��ļ�dZ��
iQ��	�;�u�X�Kƌ=�ّ�𚍬`]�hG7i�vMۓ����k�a	�مm�ϩ�k���ݫ�F��69���)�ڂ�܈n-
S�
ͭ���5��V�ݞ�I�5M�-��8 �6���l$��Wcc.Ώ�R{^��uk(潷O�gn�Pl��<���C�u��\�m���[û��-�F}�n�mۨ�oj���luɣ��J��N�)��A�m�=5��������d�I���r�[��8����Ox��گ��� �B��qܚ�M��a�I��Ξ�l�8pj�AYS1��K�%Wc�e�ۧ>����\��q���A3�rGn�W%��tu�sq�!���+���-�$[4�	���Ի��.�f��3�5�ԁ��I��{0t�8�<�����.���1P�r��Χq�#�z� �6����p�[qh6N��7��d:53���YgO֮���9Ր��G%�d�%�rp+E۷�+u\v�3[�e6�JuT<�#̗<v��Z;M�a�q�϶�݇�>1��tƶӐ��Zˊݡ�ǥvy��;W9��k��y夆�:��{+��jx�]kZ�Y�sۍۭ�+S�D i0r@Z3���]w��v��]uv�U�|G���][ًB��m#.ݬ�j�7P�P����_|�y(�vQQ�`�����v�k9�}�z����^�΍�v]�H���e�¹'�e��#:�7�J�&
=�&Z�Z�s�bK�+�4�e^k)]J^�h�Ӱ`�=v�q ���vʸl\hu���G\���'�5��E���U]C�|ګRݴ���)``Uo%��t�R\r�G0�����r���c��ｹ�|3�
K:����jtvz�E�+�fh����-�ٷ:�Q8�.�x��V���d�:�ݕ9�ۅT:�D�X1s{D9��&�p{<�.�[�֔�a2����z���fs`�t2f��H����5g��W�����;'u�wX�5g�C,�6���G�c�s�������y���|i�����g��g1��r����>��g�綺��yg���S��`���a�;�bv�!Cqz�'=zb/A�66^�p�C�+4�C��H�5�rs[KAr>�V�SXY�.ݜ�0y�g��#t�g���&l���)�4��xx�s
s��c����ۊ-��m)7k* �4�GW1Ĥ�.6ݤ��csf`�k˳����mz�V{Y�R5C�:��iܻ:�)ɪ��њ�v�v��=�c�wGn���o7��L�ӳv���^��%Ax�NG�m5����g���ӗ��[���&�5�u�m�U�,nvc�L�M��<5�ڀ�(����Y��ض#442ܺ:�e�Um�wiN������m�٪�;XN�����t~^�����<3n�Q�[�y6㫒��[���'6����wN��6�2c�����U�ٲn�knkض�;us�Y͚�k��#J�ڣ�M���-Y�E]"�������뭍���n:9;�qOcf�v�&'6��W�b��;ae<v�gv�=�.''������۲F���x4�ig5f[����q���Ψ��n�k�ݼgqpwljiõ�Q�;Q���6M�[���.<
I5vm��n�#�޹��Wr���V�����n�x[��=�t<k��'�8E�	�\ɧ<J\�f��n:4qGP�������A��e���hV�h��i�]���h�  ��� �?'�?������~�ӡ�@O�EA�.J��'_ڷ�3�jC��#�@�|Jrv`6�R�CuR`7$U�,	 �d8@�H�;�j�M�	�igi��B!@�s�S�/Q�	�%��6�%	[c(�6�k�l�&�:�d	�I�eI	A�eH%Y# �I! �FEdR	$	 �B$]�H@�/�UT	&"eɈYI���Y,�n IӰ
��w�)��f�IP�ZPفt��/�I"s=hicyM.��{I��.�D*���MN@m9AI8bC-�#%��I"��1!29��]%�	'T��QPsD)@��H�`���M�PI1�5
�����I�<������7&C!*d��BM�7�QI�S���Y+��e!0q9�pP���
a����$��H�B#.R�w!5��V��	Q\"Qpj��Ȯ̓`�w@�N`���T���F @qaC��-�&��e,�Q�����I��������&HPg,M0M�$� �ۭ�������b�*�I�A�)Wjh4#�,rA��\CTa�dN%��4 kd��T�+�J4�o��� ��(�dp�WiM�Sm�h�V���gr;PCHl��s��4#ǩ LE�=^�E�&,"&U���3�H]v�P1�\�! p�!6$����H��¶��PqJn'ᑊM����el�jp�x@I��/N�@�F)+�"� �$j2��AFt[Q���,�^�2!"pVꂉ6&���L�w$
^��M�6t���A�d		�){`��n��-2D����a�t� $��T1@:�XHE؆���n�M�RZ��T�5��#(�%�C b�@2��2����d���7[�ٲH�NDX��$d����hv,��u��H��D HEM茄�$09#!�E@�(�u�Y�$�i$V��Ȅ@�%\�ػ�B a�˰(
7�C�(
)�2,$`���;�H��K�l��M�,h"��gd"az�G�DX̙Fش�_phNo2B��
�r��d��B�Y/4^�2i�
�SH�ܮM�9�<DD\d)��!TQD�SJ�	A�%$�Jf�Dh��iL��#E�ԑ,
z$�H�cm�!ѡ��F�KC��1B���"4脤����:�Uu{P��� X�[;A!��s���G���3��� 
l�T�
�R�+��V�5lN���=+z2�JJa��QBQ%����!:o�JM��/GX��ot�G H1�!"u�Hu\�&��JS�.ү��F&@��H��Ex��9���k��	�:]`����ki�ʨd�!�/G$��5���4�7'BHHHI#u[,ѤNHM���uV\�.�*�	q!��$��{j� � ���U�X016�p�����}�7��+��R�VI&�B'��X�zBI&���$�jn��Ł$��i��hb˗ ��A6S�;���Xe�d���a!� B;ru��(�q�Q��CDTI��2z�"u�,�衢i0TV��ЄIQ��K!��QD��]ZD�*@�"qJ�u�5iI$�K$��җ���h�/j�^�B��\D�inb�(�4gQ��)!�h+0��hq �pl�G��^�jMWh4�2P�\B�/�Qb�j�v�R��,��$RH�R(FFN"B2&ra2��@�%�۽�*3��l�i�GGb1����l���$�$�$ Ĥܐ;S0�B�a2QA���(h�@�E�5r���H	6
�l�����H�";:K2�Y�,HM��8Շ���;Fd�[.I�'Dր��&�@.���p"\z�k����QC��@��:t1đ�J;I9�sa�A$!%RQMM��bj�1
��������awn�uRJ���HI'3o]��b������vJ@�F,3�&���HB�e2���k��ŶH�Y��2Bp1�kmRt��
�*8��D,Lnp8<�@z-Љkf!@l� $�����Z���]����5���LE�&R����h�SvH�a1p�� m�B�P��S��u�-�,$b�����B##!$"���I/
w��wqGtD�v]Y{z������8���<���+��\
`;��,�`�qd��,R�D�	H�4��e�� # ����up����@B
+�&en�2SF*�������H�G�,���t�:T9�0�[�ǹD�� ��H�tl"GU�;���&��	C!����  ��Y����?
?��DB�!REJ��(���pD. 
ȗF@h�I��?/ϟ>wϛI��  p         ��7n��(0K@�#i=��m�       vH69�Y7�q�uC{8 ����Yt䭍j�M�v���F̋+��:M��z�Y{F���(v竱q�r���mv�m�1����s^Mse������=z��u��p{v��raw�N��`R6�gֱ��{tb+��/���t�/h��w(��+4q�<ݹNw$���ڝ\��ne.�M]�\cN��n��m�ζŷF����	܎[���)�%[��S�q랋�s������r������7fgnF �����li5�*#�ew�:�y��&V��ݛ�����*wa����+��ݺE|���.8l�b�����G���^:���:n�6)֠��;Z�͞j9;s��'n7qۆH�Nqa�p\�]jx�y&�c/%�7r� ��ӎ5ѶQ���� �=o5)�[]]8�j�N�.��(�6 ۱��&o �j��$�A���Wc����n^��m��7scMXz����6��<j�I�Y�3ܷk9����c�̛�ޗF�l`G�,��v��q[����θ��zy��a�*{�#��Ʈ}lv��]p-�AS�ڱ�A�.y��=�8y�����&�r�qo8pd�1��X�m@����2�C��W=��V��ݭ�˞6MK�F�y. �V���n)k��wj���on�{5ӝ����]�-�uŦ՞gܻ�o7)ڮƺ�4>;c�m�]=-��S���vM9�����@$����[�|ۧ\wg��\<��9����^9fܾT�mg������&�ی�����v�ۣv�K8�^���urT��.��s���R��f�%�a�.���zPۮ{S`˻<`�pR��t��v��7a҆��.�1��l]-��8F�o�ҺٓG��N��DN5N�C�����]����R���z�m�'�aL���<�����R���@����B�k�g7c��Z'��$����`lq�|�pu:� ��NՄ� N�uN� !͇
`���A:��⽨<�G`�tu�
f�Ⱥ6�G�to�d�;M���'y�&t���M�l��zVt#�$2p���e��]	f�&Ft8�r�C �
��W�p6)Է��G�Y�t7�X:l�s8��1�c 9��4�`�9�����ݸf㛄�`��w�ͷm���s�1�j��8vb�
t/g�m!�n����s��\aJN���:�9�	�{=y�����Cs�����=����<��D���8��v:�['v�7�A�� �vg�d;lw$����uv�q&��q!o���.�-����w\a�u����'��3c��	�d
��M(�ꋔT�B�>��*q�"v�&Nx�W�^�����DpS�9�>[�:I�|a'7z�I���I>މy
b$PrIq�O����p $v�6�w&��u�M��f5�NB&7����n�k`_�,ى-i7���ux��}��j*�RQU$�a�y���y��/��{I>�����l��=I���C`q��k.^>ۼ����6$����"�(
4*���d/=3��wn��۶�hz��ѡx�K�]10E��H�$��]^=��{{[��f-q���+`	v�bm�HP�r���7�w&r>��"aA� �d�s�0f��B��pafJA�p$I	�	'��x�>�+`_k���$�.��OCAJDڢT[;���ۺىi���{���RN���0�.&N�4��-�J���=�{{+˨��s*SC�M5RI*�V���m�KZ��qp�L6n�`b���n�o5�SL]۫s��y79	1�eNk�y���u��=s�E�1HԦHM6RuP�� ��ml��$��y�O���$��/ D��iԒ-�\�y�%�&ϝ�V�˹�������l��l��(��Ru!�>w�[��fȴ��G�F�']�f�Z�����_�f�r���{�n�K~[��zhB�$	���������l����衵#(�J�bKO.�����ml��Z�O���]�kq�D�Hl��������>w�[��f��5�yT���B�U!�ME�:��
�`�˴Q=�ݮK׷�����U�oH�YȨ������D��w&��u�/��f���0��ml��y�:*GE*����qw��'��ƒ{��RO���洓e��x�D��j��UT���s������ŕ�wu�/�]��N)42'U
�l1i��ql�L6���d���d��'�f+6��%�:c�����k��c�4& H�!UD�O�s���,�U��S�*E�/�lZ]�̮�s����lI%�_������q��q�n^h��b�sa�`�3�hôv���Ov�γ����]��IW@�z����ad��%=h��P�e${��f��n���Wo`}uv��6	vլnH(MP�������]����}��{.� _�iB!�#nE�/�{뫷�>��6�����]T�"(�B�qH#qRN��ʒN��)'�ޢ�y��k2K$ ��� HH�.p^_w&R�e@����!$BB@� $IQP���,�X�	l�38�pԫ��EMZA��� 	Y�Ò ���Q� �q�,�wkv�[�{�p�K�����	>ͳ�C�6âs�z��#q�7	d�������Ck��m����?�շۃwӱnX�;vM��YպsN�#r����'a뫯>�˚:�ok�ΈGͶ�uƍ��zy�]����f��3���J����1Ů9^�K��mW<v鎮ݛ�1.sT�����v�v��{n��;�M��D/&9gs��V�ج��^�Xn+�������q�Ŋ��Q���8�D��5RIT| �ߦ��n��k��$�'�G��aFb%(f'&��nY�-&��f=�ܬǰ�no�l�Y2�j*�U)ԕP���{뫷�f]��y0�K���pR&�&�9#�bO���`w�`w�,�f��1��5j,n:%2���_{s`w�,��]���ܳ`b�wv��y���v��!�݅z���ى���0�g�=�nf�N�<���w[�[�/&����h��n�@�v�\�n��xԱ!��D5Dm�6�Wo|�]��r�2]��l��Y�fl6��)�cA���fU� ��ɰ;ۖo4�gWhw��)H�G"�Q��L6����I$��f=�}�ǰ;���SBj��:���&���`]�c�����4��}ɘ�tY�n��DӔ:��&��j��W٘�r��>��������������J�UǯR�G��]����̹���;���vm^:�D1�],�c3��>*�:�����������ۛ�����ݽ��!�&�9#���{ ��s`w��{�U��%z�2��(��M��E${ �^M���m�KzЄpd�	+��>VӉ�JbB ��H��o��fd���ՙ$��Ԅ2D!6ܒ�{�yROo��$矼��}�ɰ��bM��D5�H�~�f��ܳ`_nl��o`f��?���"��-�(l�v).v�=�q�S�vtf냎:���{�uú^&�灭������� �+G@>�m�z������t��� !��$n����7��ux��&�ŕ
��r��t���6{]��;��6f�fL6�y6�.�V�N*N�TrS���y٘�ٓ�_{sa��qoJ�֟O%����P�B�L��J��v�#T����2�|�fI��w���&�rG�8��-$��y8n�����{�m�X�U�<G^���/r���S&�$rt�$Y7M�N�:���=9�U�@i���6'%I%p켔���ʒ{_yRN/{ΒHüQ�Ie��rJI�}�I=���'��I'=ۛ��+/$؊�CP�������ww[1kM�e��ux���>ډ�I�TR�=�i-?�3+`e���v��4�����ƚ�D*�$�R���́�J�^>}�ǰ8������>	���������t[~嶜����v�Wx�q�W�����H ���M>G��{:a�Īޗ�.�������./<����$|	éG�tkoϠ @9Ǳ���{i��7N��lN�6Ht�`�DZxc���[�M��=z.�[���W	Λr<t����Ca3�ݢ��Uc����������|��#���F�����m˞mr�Lľ�!�z��o$Q�N��ƶ�z{n���g��n)�q=6�󭌪�� ��=g�xϋ����aݨM�f��u�����t�\��y'F�v'�m��n�߾ݽ��1��h&�,`�W��j�����3��띻ݓۧm�Y����uN��u�8�o)j�{Vۄ��u<9_m�������w���wu�q��^M�x^5[�:�)*����~���6|�2��^M���m�5�-&Υ�͸�j&�MF�`})*�;�gv�O@�V���uEB�M�%9#�f���%��ux�~���bd�{ K��jE%R�TrG�;���Z����>��{�]��1/�c�ST�5E�T�#��$��<um���
��iK�5��R�h]{e�N0����M�Aԏ�_j��]]��ˮ�ĸ�����WX�����u%E*����+�?�	������B�2�����:�1
����V��+�.�u��k��.�~k�����#�bX($!����~$4T���~�2љ�?��"E�FX�$WUH@���s�`w��߫���ii�.�yI�Ȁ��T��=��U���v�������$�H���(ڌ$mF��bZwr���^=�˫��ē�%���cU�'N(�����{�vY�3_d�|�ǰ>�v���.�m�M�G7-[�_n�aR��c�q���s����1��m�=���]��Q�%�k^����~����`r��ݮ��-q���:�MQ�19(��������l����ۘms�����X1T*U'�$�k����v���S�#��K�T��������w�W��鯵�f�j��)j�;�r]�-X�5N��}�tJ�?�� �a����~sSdi�K�D�<d�Wȁc ���@���|�Z6�
^�D���[� e�P�0``IЬ�uw��~�{z��.�WEz��23R�0��LL󒽒��NWuY9�w�u1��_�^A݀�h/o���R�&��>�X=X�#iN:"�mEK�\ĹKz��V��37�Pw��e�>~���K��=�q"��h�s.%G]�,�0�k�yb�:0J��{��*�+ٛ�a��값Q�^�9K���gX�ZM�4k�������+� $�$��O����"a�h�x�wyMgu�d���uD�0 -��	?-����}���V��=��{����(�p����Bf��M�	��q�^w��W�`�?�2)s��&pr�[b��n�%�,&�lc�xJw�Nۘ��E4<UA�b����'�$EΧ:~�ݧ�{.��uU������9?S��0<_�óE�t:�bH�����z����-����������e8���d��'J�*��Y.�&o{�2BD�+]����IȜ�?�M�R� �򟓯�����zS+�i6�#���d�� �����^P�4�^��������4� �)r������wB��&Դz�Ø��8o���B���/Gc��ÝpM+��h�K{��Q�&�ړ�׉��q:KK�G[���i]��y�;L2,8�۰��L �&׬D; �T�A�FEH1U!�%E;Z�o*H�������i��e�ě���6������?s��#���r��ו$RD���du�>��c�VT�I�==]��
�x��fo��)"���Օ$RC�bs��#���w��Օ$RA���du�O��f=�1U�\1p��8��qk�ڶ^	���#ڥ�qΪ��k����/�~x��.��m���{ݷ����E$S��=2��H>�;��H�+���I�=�{��rb�d���w����)��� 	�}�w�E$S��z�H��;쎠"��1���Dd��oZA� Zϻy��RE9^��*H�!
��;�:�H���>�RE$M��]+�.�ba�n��u��X������H�s��#���w�ǦT�H���*����05k~P���-ƵHZ�[ 5��>-=7J&��fR�@����!$���h�^f3�3d0B}�kE�̘��8R1��0@�P�Q��%D�� ��2:�H���?.}r�X�˕w��"�'���#���D> (P_{��=����Q��=^���,�T*�QW�y5��n�8�9�ڋaj3;���J/ƕ��d�Hax2f,�⬦�1�d~�H��}YRE$o��GQI���>T� TRD����E$R���*���Ī11*�ʒ) ����:����>���I�>���#���w��VT�H�TRA��.]��cx��s����)Ͼ�9RE$O{��GQ��E=��Օ$RA����GQI�b�eb�ė����*���"�$P��}�}��RE=��Օ$RA���du�7g���I�=�{��^.��ܢ��w����)��}YRE$>P"��w�dw�N}��ʒ)"{��:�H��D��C��:�!�T��Z�Z�j����Ʊ1
�56��F��_|���>��]>~?�  y�tث��6�����]yLuR�
�cC֒��_m��:��On���6��^�����bm��6���l:7�c���,�R|w+ǥ��r�v�$�gzm��n���1�m��4j���h��h1��\[�1�n����0Q�8��X�vy�m�K|)�[��<����]k�Z8�Y(�\ro:�r&u �v0����ր$�!�T�wn��=�@�mn���`���8���6�[�oYz���񗳡�㳣W绸��kr5T∦J�:�z�i�s=�N��)���yRE$O{��S� �RE=��Օ$RD�s��1vB�L8���9E$Su�z����H�}�}��RE=��Օ$RA���du䊅E=�#�¾jV1r�/��"�'�w�du�N���ʒ��s���)"��{ו$RD�o�OF�1�e7+�GQI>H
��=�eI�~�}�GQI�{޼� �@P��s�}��RE!���^%Qs���"����#���|�N_�}yRE$O�����)"���Օ$RD��ՙ���㳹�z���ж�xH���5\��<n]Ak2K"Mwi�����{�󖃊[�g9E$Su�z�H��;쎢�)��}YdRA���du�N{���u���IUR�� ֐igݼ���HR=%e%��'M�)��+�kuD���b�^� SWMHB�"U؜���s7�|A�ȥ@*A�X@XB> J�k��*H����߲:�H�+���O� %E$�����*���*���mk���ZY��*H�������!�UZ�v���ʒ)"}�{쎢�)�Oz��(��%���X�eI�"�A����E$S���^T�I��}��R@�T������ʒ)"x9��_�!f&f�8�GQI�{޼�"�	�{�dw�N������H>�{쎢�kK�O�<t�^PhU� ��HJ���np5ݒw�xvAu�F���	QI��IF���f�+.��^T�I{�du�Nv��ʒ) �}ﲟESqI�{�*H����B��SuW�du�Nv���J�H>��GQI�{�*H���w���'���|g��n��R�DnH�� ֐-gs=��E$Su�z��z��`!C�˹l�.U������n\�O��� @��� ��[ ,��������< #PABxc���Y|�\�$aռ�3�Vj���*���)��*��`�4Q��}�wyE!�/�W�i��k�ޫ��P�2�Ss8�r:�I�߾��H����#���s��VT�O��A�=�:�H�=�K����0Y�K�b��yRE$M{��GQI �H"����ʒ) ����E$S��z�H�!���U�U�������չ��s���[d�q�i�gr�'B�g��@۫t�5~��{��%�p�/b��$S�����"�w��#���r��^@RE$M{��GQI���+)��m9RS��ZA� Z���k\�J�v��ו$RD����E$S��z���T*)"|�x��Yd�3w�g#���v��ו$RD׹�du�""�QN������H>�綵�ZA�,�V72�@�UNT��h�~E�(5w�du�N���eI�{�w�E$�����$qM3ChT�LBV��ѥ�Z�H��~�D����ѥQ��ȵ4iI	`D�O�*/P��<��"�&��>��eಛ��1��RE;��*H�������)"��{ו$RD׹�du�O�V����]�� 6��ݶ�r��mvUS2�t���N�Mu�cfc�\�������Y���E�T|��H>�}�GQI�{޼�"�&���)��$S޿}YRE$N�ޙ��M��*����k\5����em%�F �>�}�GQI���VT�I��}��O� ��Ŀ��Ys�Ļ�.��$RD����E$S�������
��;�:�H�+ﾼ�i�tYoYD���T��i@���VT�I��}��RE7���*H'�J��;�:�H��z�_�K�r��G�i��k>��ָkH^*w�}�eI�>��GQI�oެ�"�'s�8^���0I^�r�{�.�bf�2���}
����]=͍� �!r8� ��G6��-%6&�5��?�������o���m��a�^���V[��K�%'TكA	-��:4�	���/8M<pX���l��t��l�L=V���x<부ʎ�9F�::Qt��N5�]�ca�N[�\��y�l�5��_�{��Σ����7uv����3�g�É1�v��n��풰k��63v�9�7-F^O׹�n����$a
�%�7p�d�S��9�:aav�X�$��Wt�"I� ��:O��)?����Da��3�[���E$S���YRE$Oo��GQI�o����*E$O�=�:�H��D�^)�0r*��z�i�}w�Z�b�����VT�I��{���)�_�YVE$Ny:z%��e�*񌎢�)��}YRE$OM����!�j)�_�VT�I�{�du�H�wǂ������W�VT�~bQ>�����)"��}��I�=���E$ Pv��ʒ)"nM�z�V�ي!�U��q��u�M�}�ʒ) �*{|�:�H�;}�eI�=7�����|��}VK���,��܅��؈�z����<�<-/$\��b�z����{����W�N՗�Y���������쎢�)��}YRE$OM��*��)��yRE$Or�>��X��rU�%�2:�H�;}�d�G_p�c���*�U�}��tUG{��ۅ6cl,(d2 D�$��U*)"ngo���r���*H�������iy-���5��1�^t0�9RS��H�N{�`u�M�}�ʒ?"E��s��#���w��Օ$RD�o�Ҽb�.�&Vo8�QI> /o�}yRE$O��}��RE;���*H������E$S��aU��]��X�wX�b�H��{쎢�"��߽YRE$OM����)"��{ו$RM/%�^^7G�UP"B�4���ϲ�v�z����Z�:@���[�kFn�����w}�kɘQ.�1%�*��)�_�VT�I�}�:�H�=~�d>H
E$O��}��RE#���UY�����eI�=7���|���������H�s��#���w��VPE!����V:�tJGQos{�\5���_�YRE$Oo��GQ��$�pJ��`��㢉3+&&��@"B ��#1E0��L��O^08��[isn��4-	P��� iT��!D��@0l�@q���b�h1��!B�lc�0`E(��$RyT$S���YRE$OOs�`u�NT��*�]b��%ٌU�+*H '���#���w��VT�I�|�:�Hy}��@֐iz���r�j�T*�ָkH�o���"�D�;�;�H�+ﾼ�"�'���#���o��*�+1��ꍭ� �k�ǒϭ�0��ۆ6�S�-^8�B:�K}�����n&!���I�|�:�H�����I�=�w�WQI�oެ�"�'��x�bʲ�+7�g���r��^@�X�QI�w�du�Oz�����H���}��^ѭi3ZY��7��S��ʒ���H�s��#���w��VT��"�Q>����)"�������H�zr���+�S��1��RO�"���Օ$RD�s�����o��VT�M�k�}M5av����C�6J+�}���I\�]���X'Z.`�ֈ�YM_)�ɬ�4qM���HĞ�1��E$R<�t�*��V0F���ʒ)"zo��QI � ���}YRE$O��}��RE;��*I� ��_^y�
)�RT��ꪪ�u N�^�t�;*={����à�n����x��{��wշI��T��roqk�ZA�.�����E$Os��GQI�o���� J�CK�sދ\5���-cM�(%JF�*H������� �{��*H�����}��RE7�c�*|��f��K�x��A�m�꣪�Z�)���VT�I�~��:�| �R����}2��H�{��#���t�hĿ[!X�V*�YRA@�=7�{���o�ǦT�I��}��R@� 	,ɞ{֐kH4�iY�D��4�5�x�QI߽�L�"�>���GqI���VT�I�~��:�H���J,��ŪBih���{�_�?-/�RB�y�3����e�*!av^�%��[P�ߘ�Pr�8�r^�x���-�.0���D�+�QԻ��Y<����n�#�Ni��
Dd�U���P�͛AA�Y���/ʒ�!�[�r-��O�O�!��#깜�= �wXù��Y:�����t(�$�b���I	A)�RX@��D�ے�����s"ᴩ�}m�Du��������K�#,��@ �E��	�}R�u�n����P���k�e�����X�2@q� ����h)Lפ�vx}��~ �}0�B�.C7����)vb3
����%�����I_ǅ��S[N���h"�-�A��Р���'��� ����4Q��U������`w1�����|� ����ѵ����ʺ^mw~u~��aU�f/��+ټ����n}� eĄ���#��F�B>$_���0�����<�ē��uZi��ifi="��?S�
	D�y��71����f{s;�A����9	��́���]7����{e"����7xQ��=�y��ťS��;w��X�m7Ö�:c�����o,���^ߥ�c���
9��A��/�Wx}ݹ�J�)$�I$�         ���Am��Y�  �8k�-�{c�       �����ͱ�plSF��r���M�3�e:s�[�簸D��SM���3�a� I	�	�}���O�Ҿ R�Hk�+R<c�l�1�� 7$@�vٚ���z���v�Ȝ�����q�����rvȌ��6�몎��F�m�KO^6�S�f�]��t������<s\��nۦ)�]n۷m�n�[�L+�]��j��ᷓ�F��9~zw�s�v����P�4��ɞs�W/k�)�L[�Ùg�����v�`�ĩ��cV�N;@Uѽ�e�k�+i��x磠M ��F.��Bc��vܧ\�e	#�3t�co:;6nSu�r֫<�n9ӂ�]�[x�9y��&�<�+ɘ��n���:�v��8Y;g�S�;1�]����q��ܸݟnD��[��`�v��yr8vz��G<U�n�q�g��Gfzp�P�Zzv'Y��ۃm";�M� U�{t�u��\;rru���h�B%Ӻoأ-�ݗp��zm�Y�Q���7筻r-��nYy
�����Xw6�r��� ��{��^^З&��[�5�q�of�ё;'��\]�����˛g]�u��[l���ہ�v���O8�7e��"g9�t��I�:f	0�׺�2p���J�����h��lE�:�q[��j��q����$Mx��7D\�tF��,���m��'d��v���t�Gg=��6�]s�xFP.�s=�����I��p���8�v�3����sƥ�XWgm����z��¦�;&��{'����6�n�y��~��v�:.9��� =Vǝ�jm[�>zv�ݴn�;t�YU����Ƽ�wVW���=d���y�S��/]H�ᴽvuت�0�e㞺#L��\sZ۶�\��O��=�A�u��P�"$�i�7mv|�˵��֘��VCu�\�"m��/A�2䥸�WM�6�g���Y�������vb�1���`�:����O���	�v������u��r]�8���a�� �"kb)d�8�h�!A^N)�6P8m,;	�sހu��������hN�c��ˎ��:�db�0dc��&�gk�z��Lt��4=x8�H��(�z	O��ࡼ��x�8����gz�vL�:o�0 K8r@ F.C6�6�1�m��T���v������\��.:���l�r�U��]��u����o���]��i�s��5�h�F����q���ip�p[w�ӽ88T��uɦ݌��+m�m��GR���λk�ZLŴ��y��:0ۧ�1���[��4]=�r�º�m�>�#~knM����3s
M���d9ue��^�Qک*U(��HF��iI׷[�����2��y���\;�t:�x��.��7)�m�ٌr��0{pKq}��ueC��:)9Su!�i��K�{=��E$S��z���H�����CQIw2a�i��K���x �tɪ*I��RE;��� ~����>���:�H�~�L�"�'���#��*D������UUU��Mb���$RD�s���)"����$A$Ow��GQI�oެ�"�'$��_�J/
����QI>b�߾��*H�����:�H�{~�eIdOM����)"����(�rPJ*���7� ֐ie��#���|�A����*H�����}��RE9���*H������Qr�wuu���u�n�z�v4m�j٫�I���x��L�Jݫ��ww�w�}͉"��w�qI����*H���{�E$S��=2!
�H�{��#���x���z�M@����oZA� ��̜����(�H� +_ ��k�:ꁽ<�4T�$�77����mr�ॐI�$���s������wY�~�ZZB�L=�Y�D��C��|���~���۫0|��D�Ss��'x�atRr*��Ca��g�y�wY��)�u^�r&"9���x�eC��*K�Wy�n�S�O9�N�[�6}w���O:E4S�B���jB�������0���͟W��{N���K�m1O���TT[I�ܩ
Ӎ�G�<����̴t�Վ�s���zOF�sq$�H!ʨ�$����{�֍ikL=y�� ̯y�^d級KZe��4*� ::���3��ux�uD�д��=��S%W[*�Va"�T�4Sbവ�@(@��O�]�����7U�y/7�1�J{۾81yw��9�s"�^D1:�)"��#5_c}Ƥ����̓>0շ��
l�US�i���d���s���T��=�ɎG#��}�
�+�ZpD�ING�-�w[4�kKK�iO@Z���Z��8�Z��D̰����m��b��0n��=s���v�;Om�+���JM |#�(24X*�U�f��v΀��� ��S��D ��J��DX�:eHl��s�ZI5��5Ss��7x�Z:�Ñą
���/�M]�������J�qÜe种����8�/�Sm�%h������s���N���V`}��'�IuW�~�����JC9��P�
n��6J�"r�̘�x��UHL��j��Vw�]�O�dX@bDJ�TB���c\��>�˾�"��H!ʨ�$��^L6��R}�T��?jW�>DD$ZsAN���7n��v8[�2l<��7�s�v.4v�x�U7C���{�3���e`9$՝�O0mj����J�A���<k�h�m���s�v����"Aϓw�ySs��Vc����H��n�Ԋ�*8�=����� �+1��\�KԞ`	Rs���7UQ16_.r����Ly�s��� �֩�@��Jp��p��N�${;w����V��|����6���{ц�OL�4�OU��Y�	��pj3��p����Tv��"�E���B��E���^��S�_��  �:�`[ͻzk�FĲn;���������is۬��ԗE�^m�Ls��6{�WT�2�*㛓�v7\ 3oy�p�=umb�;j�ۮ�n�!�nM�I�ָ��i�xr%��A�l�\@�q�j�C����nA�<�����ź�v��]�;q�Ƹü�m�ٹ���݋��t����N�OY��O��{g�;;�ޙ����\=~tX(
��(�����v����p7��h����n��7[FB�1�b;j��n.�Z3$��>���ݮ�&�u&��_�=���̜���Z\L=��� 5�y�H�9$��#��I^򤧠-�Y�n֩���G�$TD�T��r�� �+1����%ȃ�%I�@s���I�ق�UTʪ.����ru�� J�����J�8��Oy�.��ުm��R��8�j���"y�n�Λ����Y�>r#�������d3�\�]s����'PY�6�mƺ�pX�+�^Ά��_��>��|����)Q�Q�}�zp����.�Ip��{�]���&��o{�	�_�Y�*�N�QL���D�)$��Y1�gY�%�E��%2dJ�T���yt��P,B01ID�!+���>�j�����x�<��"G�D^D!Iȝ2H�}��p�^=���OKZOsޜ�^��Ֆ�`�N���T�]��s�ȎF�Nz�&� �i)�8�p�G"|�y�Br8��n���.f��l��^ ��Dy[s�<�y�v���-i.��_oujUi��
{x���yJ܄��#[��s���C"Koi�ھ�{��ksd���1UJ��$���{�`}��0��."9��䂟&� ��
`��S&�����e�s�֒MkZf;��`c�{Ӏw*��-h_c��Sh�m��u9�-�2���2p�XhOI>i[�Th�B��Pq��KŘ0`�zR�A�������n�װ;��s�^
ɍ�MF!J��I[jDr%O�w�k��|�V`�#g�W@��Eu���	��[�� �U���r'��4�~N�]g�����*^˿<tv��cr�rF�gJ�]n���{<�"F;u�u/;P��T�����o��ֳ�p�ws�I��䫠)�%nG#�5�y��x�*c�(&�u'8��V�r ?$� �V��}�1�9��9!�g�䂓�JA	$����g� �*��s���<���zO��qAUrEU�\v��x����5������h�tTyr�ڠ2>
�	���b�$�I�5��qZ���(�IEF��ǽίfu�p���d��a�UD�TZ���g��5$�O���Wt_*�������ڳ |��D+I�@s��Ӏ}����ׯ�n�oڍT�ӣunC���{n-�&��-�nu�.�g3k���^f����!M�on��N�S�3հ1����}�����}�� ��Ԁ�&.��j������DLI����֧��s+~ZBa�j���%:�5O�7��5�s��V`��9)��9�N��"�E��)9�I��Z֐���`
u��
~Z��"&#]�=�Bx�*e*�PrNp}̭�k��p*�=o�f��vb8��� ����2H	���Ii������$Q@r��� -îGY,��� ��@[��v����}���7eS�����9]�-l����\rחu��].�:u���!O���[�cv3��e���=��&��p��ڋ����2c\Z�T��6���JuZ�������͂�����7Z�z�ju�vu���rn"]��<��>ض<��Wn�]Nw��yb�v�5`+�����{����x�n;{���7O��J���F��vn���*�M�����Օ��U䍴��Ƕ�cO��Ta�'H�JA䭁��_��/*���՟�G"��RӮ��z5�P�M\�uuW�����O_	�<���c�/'<�����1
�y:�&�����$� ݭS��<�s���t��_c�c��!CT��s��$���ql>m��IOA���y�&B,s˰����컸�
~I^ ���΀�'���6�w2�EPy�&8T���h�]��N�k��t�\�3���N��n����+����lq�Bj=����g�x�ۼ� ն��DdrAϓw�y)�1eC�:eHl��s��y��\t��֍��l�=�=�0��hZT�p�
B$$�VىwK��3�]-O����E�J�ʉ�݃�-�;v\S8*�%�w�h$$���d"D F,g��0D��0v�g^��5m��	q)�����	�Wy�&��Oڕ���"L�O�y�pYx�ęIʒ�@�΃��>�� M[:�ڳ��;M�gVz�^�UE�Ss�^\�`>DO�}��9�
~�W�o�MASA�l��/=�u׊��e5وO�~
�i��$Y}sb��s�߯~����p���'�U�z��U� ��m[:�|���"��:�N�8e^=�kI�>�� m[:�uf>G"c�.iJg^QF�p�*T�`y�3Ӏf\�ek8�'H��s�O5[��kb��+��[ϐ�_�I��h������T� U������7/?L�Tk���%�2�+�lwD��<U��|�}-�L��#�S�����;r�Fq	O�|�Ӏ�<|h�<��e���o{��[֫8�D��R���J��� �����1)�Q��3u|<�E�P�	��dUp��!�]��>���L��n<0�3�]#����-37�ˉ^pH��>�Mq *M��`.�Ӛ�I���c���{se�`,��Nu�W_�u8�=7>��D[�[�|F�_� Z1W��- _�!��z�w����쬆T!<ʉ��1�d��w�ok�;�����{���X���d�@��rI�`��� �è^&���튟��4b�B���8
�r��݊b'+bT.v���_"<|�7ӳ�<�	�oÅ�ī!x�� �đ�PI��,z��~>c��O�jI���\G��_�^��f�gG��X�"iv�N1O@@7�%����{�2�w0p�r�.b�5��'�O��KW��9|0gp���V�I����`�$��a1$qtR®x@ۗ�ız��]<�
��8<�x��'J�� �w�Oz���`]�"&���x��t�d�x����&���:$З�h4  tzu'Z1���c�L!�d6�^kD�:u���T4��t3jtp��F��Bsl��/B�&���h:	��%�K������SfE:=8�Wo:�! $RVC�s����&�~�fI�<���U�Ae��+���>Ko���<��O`��뼜�l"�����!�۫0��s��'x[h�����*������/C�jv�}���8#����dˢ�v��_���y�5�����%Z��)�u^ ��;�۫0Yx�ęIʒ�DI��뼜b�G@_n���G_9H)=
\T>P�Tu䛜���`gݼ�$���Hڶt>�� Rn�%+���.��f��>r	{�� �'=O�J�/a�ϡ�vD���2�nW	b�ȼ�B�{w�+�f�����iR����t��/ 5$F�@Y!ֵ�˭����/e�TڧU
��-�tȉ�=���7I�@^��ͷ����v�|?��e8}�1Q�=td�rqFͽ��m�S�Ɯ��8�l��f�߮����n��L6U�]ݝϵ���S���q-�z��`{�Y��lq�P�����`	V������`�s����Ah�z�*�I�ϻy��Z���"y.}�� �'=�ݙ�PJ*��Yuw�9ݧ=ϵ;��S���4���s��$�M������U�	RS�۫0�T���U��Jd�j��,��yZ�d=�+����G��NG&Hb�p�k7F)���|  %\� Jv7� ?���H|��dn;H�#�1u@�3�e�f�VyRŜ2�������:�)f8�t����v��'���c�gsjx���Hq�v�`��섭V���<P��k��r���<�;u�'pfs�u��W��n:9JUvV��c�����Wl��\�U�@�ⓞ��^^۷LY���^�I�f�Ɠr�g_���XD��5d�.�6B�\�V��=z�����ݗ��n��I�X{�W'Y]0~L6�i��H��(u�Ss�{+���_n���S��#"Aϒw�8���ݩN8:�����s�֒i��g��s��	V��p�s�ApT��UU��� �7=O۪�qȂ$n�����{��EV1b�cN%J�����*Jz�uf����-���NH
5ʛ��<̭�k>���wy[�y8�FUc�T�F:C���²xԜx��量kmÕ}�����X��P�����2ET㒶}w������U��s�Kn�����Ļ.G�J����V���$�5I4�������,&�YtK�cR��Z �IQ�! ���:�e-1D�oS����`��,�e䄅�n�L�ˡ�n,$ �{R@Q�<\����zV���՘���!9%I7dQeU�t>I�����-�����Y��&�IB���[�M���r�m���� ��f�����~)y��QDIU*��l��� �ZT��ϛw�|�)�"5��uT\k�k&݆�v��6�i5�qv��br���krr$�!Nm	�-,��M�ۅ9t��$�)�%xʒ�Ȍ��y�(�R�ה��I�[ٙ9�%��:��$� ݭS��� �<l(rM�IF�S{���y����i�$�& {��dZ�BI�D���f�BJ�ALA�'n��̓u߻�5$���G�A"�d��<�����8e'=O�+�|��O<���S+���'�M]��Z��>ry��M��˻�pkI-.��S
<�����㮮�'l=�䒶#bb�sW/N���;I�m1Ji��D��R6��R>��{Ӏ|�)�wV8����zOF��qwqr��UE����ef=��w��ux�?�2s�6u;����R�T{��`��z>G"eϓw�y�s�|��US�T���8ZI�L��}�zp����b�-��M�EI�D-h�L1m��ߦ�	�C8q���+w P�kH]�{��-xT���A�9NHM��?n��G#�ۜ�S�v�=���n��xN��$n�'&��8�p�l�S�q]��|�8켍F�9�[��=����\��s�}���}��p��~�K�<�y��2����L�Ȫ�${{ڳDDȕ'=ϵ��>T���-+Śhk̐�����{�̜�ǰ3�y� +,�bLE)EU�t#��ɻ�<��۫0�ܭ��>]��IB�t�����ef>��ǩ?�JN���+�G>"9`���B�*(LQ�����w1��XW�ϸ����D��[�^��ڋh!e���ǉ���|�}�=Еz�]]j�C,�1N��3%}� He��
�����N��0�V� :Wct"�G+�1�&�:2ׇ[v����eb3�X�P���t���lI\��<-x��1�u��ӷl�H��z���:����pݺ����v�&��rY������8���a��㒷V�%"q�<��i�<���!�7��m����ӻY�������Ua5<fԏA�<������\���^���������{�n����Ǩ��89�]�F��2�ٷd��K�WIv�}s��f+k��9���	%JuQ��s�8������̟��a�M�@q�<q.��j�������6wUu�L�|��Λ�����DL�4��گj4')����sޜ�ǳ�m�O0�9����R]EvY�����%={uf�Z����K�&� �b"�Ƈ"�d����s��k��%i� �ɻ�>T����[�����N�gy�b:l[�8Oi��O`m�u�l=q�N��(f]q�&;����~�{o�򓞀��J��%.2A�O0��`T �Aԏ`c��':��_�i�T��?s|f�W�Ii�<�@��j:�YP
z����Mr�̓{��kRN�^=�M�ά�k�EI�ꪪ-�M��M�@[�Y����9�|Ӽ �=��ԔEHrI)�G����s=� Ǚ��
~�W�㜈���8�8�UqW3EEU]U^`;����U�%h�۫��Z������"i�b��P��c�;8�=����ًt:�xݤ�8y:�:5nw�4$�T]���`|���{ug ��ǰ-/��A֥@D9[�� �+G_&G�<���)�R�q"�a�n&�E*C`z�=�wW�f��#�f@��Yui-v�HJ�&a���n�Y%90;�h�d����F��Ii�Vu��s�e��`u.ڽ4��.��eU�`��z��W�|�����i'� B�qYd�Y5w=O�+�s���I<�6}��ֻ�c�/�*Q���ONA JC!#$-]y�Ht����ݺq�N�d�e�fj�#BA�^:�����������j����6}��FHy�����<=Iʨ�1�U)���˽Y��Ȉ��u���x�mG�u��TT�UU��o���1����}�0�}�� ��U�U��7*� ���ȗ�i���o�fVG6�5UP:Z΋v[=��f�"�:o��U_yH8���s&D�p�J�����1s7p�OCPGڻ�+0:�Ǘ���T�A�{�p�&/�� ݭS�ԵV �ɏ%TAT8�Gnx՝�1�=y�-���7G1�������C�u����H�5Q���l��� ݭS�ԵS��<ݳ�lF�Q#����/�U���Z��d~��`n�l��s�
�1��
�{}KU`%h��&Z�� J����>W�)IQUTm�TSrn�֓ｿ٩��Z����~��`;�Q3uqU37sWS5g@[�Y�>s�ĭ9���\�Ɇ��}�R�M98����ڿ��v��c���Ծ�@�~���G�s/!���� "�`�w�������=��w��݌��|j{)�0��/�ô�5酜��p�Z�"Q7���4�yZD�	������\��=q�"ӎ�9��+�iW���co�AZ�[R�����p��(K+�AC[H�]�>�����A��k�eF5�B%�x�[����=zK�ux5�����F��U1T�P5�UzК�m8�SUĶ�B�%�(* C%Q�h�$����'Y�ݔ&��q�21�y,������	T���M]K���������h�@hM���{�F)��]���q�p��ZC�Kb�_�7E�=��xPx���Zd(m�@�{p3)�Ĩ�
�H� m��7��vm�6N}���sZ�I��atxѣp�D�;Q�8>���)���o����kNv��M��B��R�R�>	ƾ H����hw�{ TmsN \�[�2=0"�YVPZZ\�*��L�L�d��殆nO�//��i�{��͌H3����� ��s�Q1��L�a����>DFmR&
`,� U��VZ0�h�i5�T_Ɩ�7q=o��c�5�gݿR��??�H�Q�#�U���Y��U�>�h|���tr�4-���[n�&�}��׌CB���%�O����5T �+h���<�?]�g�� �����1I,�9��VlԴ,�#& V�Kޞ����｟]�>�-`           ��7�)�p )X�m�t��   �    A��K����+��x_�)��,<�+Xq�pu��n6x�M�=z�v�%�Ϸc��8-�;��k����Qk�.�ŦL�Uч��������#�u��N��n���v���蜉���]|��ɸ��lH�i���-]�@ܜ<I�׹�m�Ǎ�����q���qێc���\`FQ�<+x3��d�hrâ#f�/:9����	�1�4=�f��tfڭ�AH(m3NA��Zs�%';��]�W�C�:�.=6^^ʖ��pc�@�t\G1��$;1�g�V���m��_\1ӘDT���n���'a�œ9���������|��!"K:�cuN����>+^M�]��&�nX�l�qMvzܞI�q��{8z3������s�y�&H80�&��9��qk�4��bo;�-�f���s�b�2a���N���ytk��9�ݸ�{l�<�ܷ�C9��Ї�-�;l�.2g	epI��+VJm&���l]���w��Md�ޖҸ�Hk��#����3�b۬j�׃S燎7G]��4[:��θ�&4�Xs���Þ��M�q��[u��h��įs��۷@Fh�G����gc�Sn�[v!S�sH[u�n`2ё���k`���k�Y�a���Qk�$܀M��β/^�m�J�'�7E��%�[��W3r/@nm�
�[h���̓sګA�Y�MXX�jV�'l�v�c���*�"��.x96��.�Ԕ��3Ӑ���=z���Nͩ:֓��|c��������<�e��jRه��`��^9��d[�V���[n�eW\kt��ض�Bݝ�V�/5�c��cb�s`HH�٣����I�K�ק�I��q��˥��伙�������;8Ṟ�9�#�85f.�e�i����:]]�n�NH�1�N��p^}��
�K�\��/�ђ�m��c�W�t������:*����=3DNN��p]��S�q�z#̌�u���M�,��WEp�$B8N&&�/p%�)�Z�v0� ��m,zp$�'x�D�w���u��k�:�m�{����a��-C�܏`�t�'F����N*kl�)�u�#�r� =^:y҇��8�`A��h@o����h ��y�N<�I$�Iԣ�,` �ͽoV���뷥\rČ-����\gom����&;���ѓ�/<�.v[�Ug���n�v׵�a]�v����=q��f��z:7�s �v=C\�')ŔЗ��k.tӲ��l�MkG�\�v�<n5�ʼe��n���ݵ��t�49��z-�	b]q��i5xR{�ʼ��3��p������Llў[�õbUb����R�QsX�U�U�+��E�[���mٻG:{1,vN��5kOdG]�=n���o1�t��'r����m���� ������>s$�y�(�)3G��ܪ$�������$�;�O�I��Z����=�q@��5Nw����:�uf#�����9�ԓ�}i��G(jTQ�H��~��}�%I�@_R�X"|����
$�J�5
�s�[���I-{�������2���Zkٍ�J�� ۉ�vݚ˷V�#��v�rwK:��m�̜t�s1�]u\څI�8��B�J��{ޮ򤧠-�X�#��N���9���N$�pK%xI��ߕ�}I��>i���=&űC��Z���WE	��M��pI!	Dt�篜߯+`gՙ��kM��<=I�QQL�ԧU��f<�6}��8�&_��X�'=G�x(U7@L�*��j��G%V�]��u�}�x�]�s�Z��:x�ܧ$r����U�|�T���0�j������¨C�z�T�7M�jT�Rm>ً�zP牶8RyC����y����my�qn��O��k�<�9�۫0�j��Խ��b15�p)�l�=����8�E:�t��� �V���&M�$(t���BjI���հ3��ep����jih�kٺ�A� ��C�|0��ľb��1��9,��>�в!Q�$�������8 ���4Tne]�tK��� ���/n��|�O*�հ:Ϋ��"H�#nS�n��}+Ut�O�S��@_RJ�����>ȟ�{=�K�l�צ/���28�ɍ�]1�������L��f��^��[:�iJ�����6��l�Ut�$� �V���Ƃ�7(檪�8��V�-&��M��i�@^�Y�9și�$�M��NH�J��g�\痕���M��<��u�Gǹ�(�]ԄNw��ȟSN�Ԟ`>�]�Ôr;P�K���(K@�cH7�M=�zzAN��qV���KI?���p��5�p
��s77u���9
�:���X�/+`{K����F�qA�� �Ym�5��9����"j6�^n�ч�&�ct#v���┝P�Bj���1�z�}Y�\�Z��#��$� !p8���n�\�����U�}+Ut�՘ϵW@�>]Ŕ��F�S�n��|���j�reJN��4� ��'EQ77wWuUW]֧� �']}KU`8�'�ۮ���`9��&o�Uu5y�l��#�֓�����/�V`Z��oBi��M�!��؄�4!#@�$���h�
��=&��hf�1� ��!N��h�O�
�8� D�	�I��� !HBA���r�˼c�Ib��E�2!$l$�z~=�;��� �B�q� �%u�u��kz+�V�q�`��ˈ���H2�`Z�*<<�<�����ӧ�p�q��k5+Ӭ䧜��;rI����rN^7\b9�����ވ�v���]��k�mٛ$�ލ%'s��-�9j��6��lF痆à��7C��n7'j^����ِ�z�FD͓�0�)��tpN���w[�<��趀('���f{��뷻n�����E�m����\ �9�0ԝ[ۢ�4�i�=f���kv�mTm��NHܕ�;���p�fV�Ϯ�ZB�y���~�ב�q�F����>��u�����JN���U`��j,D"*Q�䭁�]�8����֛����<̭��]���Uރ�"v�Ut�i�����㜗��C��HU��+�U��@_V��r#�Ӝ�'���O@q��5Mc���.p�\Յ�l�P��uh.����8S��>�AAn'�C���r���+��'�'=}�� �m��/�uV }���MBIT{>��r��3Z�I��I7�� �$(��EEsR<b��y�>�I1Y;�{�e&1Vt�,�2�x:@	�XDI�J_���S�Xʒ��s�#�9�Pɺ ��UVU^`	+g@_R�XҒ�����p]+<R�������%��u�z[u��V`ݴtG<f�5�j7ɽ� ��el/e��J��ԵV �ٚeUP\��U�N�:R�)m����s���F6y=��5B�����J�4�Q��MF㒸������l�����+`}�v��H��Z���`ݴu�2?RN�Jn��j�|�&B������W.f�΀�M:ԓu�z�26����z�dh�J��O�i��`�(�� ͷ��X���R�x-�6��V2^]葘�# ����w�����>]Ŕ�����:�)ھ��r'�Ӯ�֧��m�o=\��y�	M9Qʒ�J�}�� qū����XҵW@��Jb��R�]��Y��oˮ,�b�����-�ْ۬u�.��1��<=f�g^V�~�[o��h��Z� �V�y ֧�ƑP�My��2HGP��Oݞ�W?$�-����jy�o���2&sG�qs733����i�@[�Y�n�/�j�5�ME��
��7%J�{O�y�fO>�������		R�� ��u�O����	\0^�an�>�1��e�D���j�� n����"����������/�t�*�9/0ݴt�s���i��y�s��Vpi.��SK�)�8��������gv8nJ�)݆3�'3p�S�q�H�t�'�k�B��\���0�i�򤧠-��kZ��fO��~^�N�J�GTE7Su�|�)눉��O0���/�j�|�M�e�ΐH��T�T{�y�p�ګ����i���$�o�HQ|��*�09>�N��4� �ժzO�y��,5�6��$�R�}KU`#ں��O0�ګ�|gҐw5��[�!	�L������B��e��h�f�y��ѓK��_S��֖5�d�I$�I$���� ��֞��ש6���ڵǞ��L<����֕�gh��8��Z���fl���w8.���-�`��s㞱y���=�V�;^�O �����)j�b�Ai7�l��.sW[v�<n�����&�3���{u��ĉ�<�ś{<mxt�Q��<�i�;soo3����\�S�z�sZ�۝�uGR�C��i�$؂��R�H��(� "� �n���@�O�G���j�bM�p`�d�^��/OFG�pG���s���<�{7R.����o�f��Ut?e���q5"��7NC`e���I-6u�z��}�����`}�v�0�T���>�V���^NZ֓}��6�����f#a$�U�NI=Ȉ��N�j�t�՘#���-�W���QR��ꈷ�����à6�?�ө�@S��x���Nb�/N����n��6�-n1!�*3rD����д���u�.�a��z�X��6`jy�}>�]O�U�G#��l��[XԈک�
����elJ�n�eUO�ӫ�R�L���3�D����l��h�c�
,ѹJB��E=BER#�A�s�"v|�� �;G@[�Y�&M抖
��pd��J�}�zp�W�c�"&Z�� =��@�F���L�\�\�_{x����s��� >���8���w���/W��^8��������s��N�>i�����s�X�{��m��:����	�ON�Nl�B'1�\��7GXL��:t�,�|�w|�N�����=�t�՘ �f&�&H�Z�T�`c�/' �na�2�y� }�ɿi���~^�R��u�-�� ���`e��?�U�I}$���z!k=J�-��U_�u{�:�Nr�B;��Q:�!!@َ��Y�I3�.b�WrF1e�	�6�U��3�}E�Wk���zB`�m�ޡơL-�űY�U!{��������O����%�J����,�B���@�A�L��d��b�L�tV&�`�~A.H��̢*F�`�p"IM��Q��c���~^�\���N��`������Z>���PRA��	�� n���	�2��[��ǺP��fl��z�7�z�x,�YY�$�|�h�Z5M�A�$6�M-=5D�����Q�5��oB���h ��q ��>E
��1�q������x���5�~�;룷�:���w�.43�<~�V�<R,�� �� ����3b'�J^�������g��(�+���brQ�,��,!%C8/l�Í�8�/R7
��	�/�r��}�џ���<3�z}D�t��;Cо(����%h�H�!�$����Z9�$,C�mr����+i��^K48x(����L���m��v|��:=�A�0ؔ�U�;�xq&У�$"m7"# �-t��]�����r�؊�H'D��m�:&]�M���Ł��
@��a�$%�3Ǫ#Gc-�&��.�<:P�@{��l�ȒM�ˑ�3��R��tN�.�o��4*=:�\��\����Q�T�bF!=��}{]��33
AZ� �����l?s��DKZ���N�����q�z�΁����#B�"�B�s�c��l.:�N��'=o�f ��Nf�f\Y�܆{�5۰�[tc���^�k	ΰ�o���ٺ�ãV��vv��4��ߓ��ժz�j�Ϥ�u�Bٔj���|����������l������u���^8�5��������MU��@kS�O�WG�re��� {Y�>Ձv�*F*����kKO�x�?5�`ժzn�g��]r&E.\�����9�y�Ya����Y�b�c�[���9���	��X���kBH��2n}� .��$�I��7wu��z��m9��� S���ZZ�f?R�r�j�$"D8e�\���8Y���C�\����n���sw�ʊ���ʩ��������-����*|���~k��Cl�
�Eŗ5E���@[�Y�l�*��F�Z���I�<[X�9�S��հ�z�Ul��6��s�T"
3d�qWW}/�c0):�}�0=�7�{�`bX^Py�N���n�6p��]�5����w��z� �EA{�B]$=M+���n��&.P\&
���2TqT�`�"˪�����'�
S|�"��I$�I${I�îip �ɦ����qi"=����;�����M��rVψ�+�,su۝nɆy^��q�.�Ĵ�sn�#����1�8͸�3m�k`9��n]�x��"�������G��ƻv�4S��n�i�mέɝ�Ee��}��\+�x��nΜtmmɸ�p<;p��u���`�d��/Iֵuƞ:��l�<�i�g`��Q���u�C(@b� $c���v]�sƤ�΋��P�i�[nm��/aj�T񷜺�%m�8�����"�Uyb��-՘�J��oP��:�t� �B#ʠ�$� >�ɰ3�ޣ ����}�1�br"B��y\�������Y�l�UtqșkS� ��`u�.��TQ�P�qG[����"Uju��� �_A���3 <�<R
�)Q*V����8����;���0>�]��=nf�f_���U:�8غ�nŞ����z�"hF�<���c��^H�
�e=MH�J��
���y�z��oQ�)��y ֧��P���#n�	R�}��9�j�5�i4����� 9�we��"��tP��sr�"A�H�0`Ňd�I�@~Z� �__"&E�*A�Iu̅���LΧ]o�f"ge�]��o� �v�Qb!8�R�����Z���N��oQ��*����(s`U\�M���Z��8�江 �[���ڳ q�r#����uUQPY!q̜we��r��l��y:,k2O"z.�=�U�W'H�(��$�I�(�I\��o� ��U��V8�C]'=d�k�QA5aUeT�\�z`>J��"925������ϲ��=��ë��Re@RUr��Z�`U�z{�%��	�� �p8A%5
� �7��x�;/73����5����­-�%A%�bY�gp�Mbg���$0%	�"As�>���9iW@�zy�]��]��Uy�����?5�`��['�����R�W�6�Q������ޣ ��U��V`U�z>E�T!�z�&9@�Q�5�}�W$�^��m�Z�u���k�����h�mcOh�����䯠-���=>J�#����\ڿ&��!P��$�}՘��W@_-Y�%}q2{���&��lPrNpw�V�ϲ󋇓e߽6�����Z/LFI�(�H����^i� n�}o�f��ޗdf�T����F�UCVj��# A�1#��3�fI�9��˺��M�U7�_o >�W�#�j|�&�?��p���&�S��J����P�5��qv��v�n��v]1���c����:vɺkj��GQʩ8�����^=��켟����M��-�4yH�)$UU9�;��=g�%x�䫠|��3b!�EQ�/R+M�tS����N�p�i&���s�]׼�%}n��"6������n����ޤ���v��� ���&�*j8T�`}�^s�w���_�̜ �s&�方�%��6�i���0��T�J�P��/�f��j4��$����Ԏyf�}�~dU�n�64H����Βnu����+��͸ۦ��{�svV���'HĂ㫓���g�ͬpG[]X�un��8��˽e�fM�,��2ԇ>�r�E8۬���pÊ�F��۝��;�2��m��:ݴ]��lM�7&Wf�c#F���իWV�	a��(�i\�]���rv2\#���3�+��DwXq\�t�Hk��29�c������ݽ���ݽ��۽�ۺ��W�qu� ld�G��Rqrqڕ����%���zbiu�B7h�L	8��Q�G*L��_�����^ yj���H{�<�!@�$��*"��z��%x��rd5�}�i�}�ǿii��x�H�T!T�������}�՘>s�+i��>�� >�0h�UJ*$���I����}���e�s�=?y+�|�����������U	"r�8v�������w�`}�s9�<���`��PrQ(c�G	HC�-y3�v���z�Duǳ&�<��d��5���]n�+M��B���u�����ɰ>�����9Ϥ�s�G�� "��9]�o�c���y�$���Bn���,T "��:HLf��u�K�FƎ%��$���"�8r<%m��Z�}?y+�ikM�J���PST�9+`w��s�/RS���ϧ���Ru�=�ѪfӢ��8J��$��{�`[��Ӏc���y���}�xŌ�G���J:�=����^ �uW@��0�Jz�G͹{#�Ǔ��ʼ#�t�9u��5��˙��ԝ�ֆqn?{�~�ܙ�f㽻����t�Z� ^���s�̐���� ;�����AR:�nJ�guf8�D������Z�`
wUu�L��<|P]�U�wUy�=��o��CS��1cwL��)�e\��Σ�H$b�wv����	$RHHH�4����z��ל����cQ:�j7P�#�y-'���W ���l�j��K�nz�[2�"���Y73��� �uW@�����)��-U�>���ρ�����ٝ�y	��@���ɺ��#�\����*�ۮ���`"�=���s�[�T�Wf�S�z����R�N>�i[6u�Z�9C���89'8v���)�z�u�4���ڳr&C�P�H�sw3ʈ������M:��y{V`��{��v�R(n�N��)����䴺΁�S�z����}�~"	��5S��cZ�I+6gH�`*�*��g7�˻X�|�"A�H��BH֗{}�+�e��:�SD���T:��f ��ۜz�u�-�G@�Ҽ/�j�ܔ'h��Ӫ�q	��6�wϰ���2�N��vJpWC�3k=���Y7quW��=��oԵV ��O@[����j�cQ:LjS�S����2���=n��z����D{d�:���s9����9�۫0|�����v�ޮ�w��V�:$�a䟵'� ������J�r9ȉjӞ��@l'7D�Quɹ���z����֛��j������ �V��v��Ó�$&Aa�+8O��ȯ>�u����`��D�xfUL�e�5VFU˧������h2�����e��pKQ@��$ �L2�����	��}= <ApPi	Kj4�z�����ٶ~e�AT��~��P���s0WȢ���}|;�����E�I�@ ��b��P�JѤ����R�iE���ݻ�om���c�c�.x����P�8�e�k�Ւ�C�( � C�
,��$�$nc�g���@�"`[a��{���o��Z�;1È�EX�=�vv��x��@��k}�6
�Z�p"h@-*���+�
-�?@�J>Ls&Q�;�%ޣ"���7/\��fx��ϼQ�ߵ(uC�˼MM����a��^���sw��*��3��M]��?�)2���v�oh�u7��A��i�0��p�~i��P�>�f]��S�ȋ�t��*s��%���*la�$��}���َo۬����Ȥ��
��
qCD~l?�?3nnv @׆M��KD6�\0`dq����|� a.+��`�qG�x��ݥ���Fɸf��-�z���1�����n/���Nb�!���#�$pj�"��s@,�9����T#U��J߷��Nq�!	�K��r7p5��H{R0n02�R���M�.�Uw���ɿ��Z�       �    ��i���&ۤ� J       �[#kq泸�Ӟ�Ϙ�x�ݻ'F��'��Z�O�I`Y���é�Y�η�S�ca��u;�Z`N�ݷj�·%tDS:�=�ζ퓞�e*�h�b� M���^B�C�o셰d�m��b�ܪ��VM�\ܺ�������&�g����9'�>a��Y�̽���q˙A�=�z�ap�vS��F��(�����0�wHw�����,�6C3O9�������3�u�8;B�\Xv�볶���J��c�4�c�W��^�]���ϐ�.s��6����F��۩ۉJ=���A�b�<��#���&놓Y���W%�vg��<�\�qן����;m�ځ8�wV�I�V�eGIΜ���AL�rB�Ql��w7!&��nBy9]Sݱ3ۨ�[r��mfm��8�'n����a�'���J��m��y�Ÿ=���<[�垄�S=c���{h���:��W%��gJ�l�`��ٷk���l�2dȕ��*���Rٵۮ�۝�Y�>cv����O
�67v$S�-nd��\u��T�Ϸl:���r���^�p1��un=���q�����-%t��f�m�wn6]٩�p%m9��GQ��vy��J�zMd-����c�깳k�|����;m��,`��ف�%��r����
�)ʦ컷s�/gj���/$�ͻ9�˺��v۲��r�g�Q�;���a��z%��T�;.�m�Qgb���݃ ��ޝ&s<���5i�&\�L�&��� ��4��=-�����$��Ő0���w.#qʕۗ�t��]�plٻewN�㱷&�,�ar��N{G獮s�t�{r^6�Ǝ^[E��q]�L�8n�ˬ������̡qlaKX�s����8U��vw;gR6X�׉N4q�9���ح۞ی�8+�[GYb�lʛ���n�]m�꺻�AЧ�㭁�PX��'KJ��ӂ;1�^/v��d��'pD�`�PCF���'V�8�<"��S�D�4�7�}]� �ɕ]�!{99��8��;!�(���!+I��Q��8�r3�
uC��,��������Ce=A�0kp0:���c�C�a�"��$Oa�[9	a���� X�TM:�G��5���Ͽw'o�� (��� �N�o��7W&���3;�(�n˭����]ɗN�p͌��[C���v���q��V���u.�olF*y��mی\��Cs�j���Z�K��E�����N���s˞�9y���͍��X:��I�$�ӻv#��s=�P���9C�kzt˧$瓷N�g�vI�8Y�8ꮴ�s�F#�b��04�&�rc-�,��Ӌ!5B� � ��U��N��dx+	�����-��V
@�F�񖙽�R�a6�����=x�E��ߛo������T���0���>���EC��(�r���n�e^=�6{3=��d�3���紓a��^�UUR	��&�zI<��GG/�۬[�líZ4�2(9 �s���=���u�y+GA�I?��"������n����:��U�8�5>� i'����䵗�7TU?"4�*tSi�v��n���pu�o��{M�'(-�ۈD���:⵽T�ODA�ou���6]�s�{U��̐~��`#TM�qd_*B�6]�s�7��_%��g8�Қ�)f���E��Y\@��I�'ҹ�!%J�kh�Y���"�""�"Ĝ��u_�@��u��V���=�o�4L]rnf�� ��}I*�����y�fg��t��1�p�T�n]��~��`���wV`>G9:�Y�:Ϋ��"�J��ꈦ�n�n��m$��N��Ԓ��!"Ә��wN����m��]���>9.�#�n����6n���:h^��j�zyQ��EX�I���/�j��nzf5�'L	���� ��cߒM��6� J����uf>s�#�"��pED�S�G#��g�\�ϸ���h��Va��\��wy���L��	�#��F��=\�;�j�W�`^���SPq�M��x���$� 򤧠��~��`#TM�qd_*`���wV`��!��`�۬m%=�}�˚��ń]��m�A��]��Ǭ�Y���7'X8#��F�
���ST�M�Zq����zx��IV ����$� 9���b��DY7vt�$�"9#T���y�e��~�M�gU�z�L��UDSu7XT����0���Ԓ��7aTUUqe��\�U\�9-&��v́��̮qq���5�i�J�-��[ۜOPj�(�3��S{'TZZ��	���
z�~�l�y�B<�hSQ�C��/&���u�Ss��Y�>:�3Q3..C��[9���&�x�����.���ǎ+�vy�{7�FTtj��&9NHJ� �׽��
V��u,q�} �'=3�K�)�55���c������*�����8����`gk3+�I���PSEI]Zo0�T�|�"em6� rӮ��4�%ʂ�K+��Uy���Kv���۬J�]�7� q
$�ݜ��&��o�%X�9tӬZo0z��̓o#�5PI���8��i��Ye$���0��憖3�}�t�V�Y��:j�f�&�~I7�� ���e�U5��.3�!�����f��G��j�L`D.@.�X�'tv�t�A��m����������۳m#�@Sۢ8$�݆d��q��ۛ�Bv�h;>WFz0m4:-��s�mn�a�x9-�A}�v�kt�vۡ(˰�.�f:�a�no�I�uY��n�9lt�^x,;QB8�ѳ�8�l�hF㞻l����n�����AE�D#R�ޢ�{��g�|K�[��p�Tc\[ڱ��D q'��0�љ-�\�K}�]��5E���Qq}��`
Zu��Y�%Z��gk3+�|˵����(UGQ��6�K3�27I�@{M��䯮"9"�8P2d��swPM�`Rs��%X8�L��4��aۈ�QQ$����7s�q�{m��5�s��Y����˞���Y��SLMMA��7��ʵ=�D4����s��%X�ǒ�v]�;�nxԞ#/.�����]2��� Y����oVW�9��;$7r˽���=��CZO0*�=~��8�}!�M�@�o�T�W&�� �֩�8�EG�8!��΢�6�"�g}]Ǆ��C��������,`�"*�"���"��{���$�w�2N{��9��Vyf���!�J�����=��>�J�>D�Ԟ`�9�I���0T�wSE�jﷀ�'ԛ�����Z�a�'�f{Ӏu?g����PrUBS�]��Y�{kT��ԯ �u*���<�m�9oeS�s��i�w:r\�l�u���sc�D����c�C�vGmΈ��I�M�����9�;�^��U�>�՘�M\J��m�NE�`q��Ny-isUG�7]~I��S�"��ʘwQDM\��w�����t����o �*�!;�
����ʭb+d�-It8̼kU�Mb_f6d���"��� !�"��������'տ_� Į�5E#5	�9RV��Z}��}�j��d�R�>��t�Yb�uɹ���۶���V���<���v�9�<�O��T��R ۉ��9��9������%ݶK��n��n�����ݫ������%M� ^{�� �2a�=�,|��V΁�=��0TԗwSE�����>J��C��9T&�zJ��1�֛>O/���T�GP��6�'���:>D�ө��<ݳ�/�H��0�Q�C���*y��>w���~�=3&�Tu	�eI��#��m��(�`h���i	R��
Q P�@�TBX�TbkIiW�����Uf���b��RT6N�W�8�y�� �I���������إ	����P�D#$`�۳���+m��tq�\��<p]U�C=�"���۠���{x�Z:ۺ� ��C�Ds�!����!"o�T�_����}��1�L����})7xڭqɓb%�����&�j�0J��2wR�&|��;��� 5f+I��!�J�$6�Oԓw�y;g@�wV`>r"u.��y�����9)�&�M����`}w�0ݴt�ԯ ���QW��p�	�a���YDX��#����D$}�1��}�+�n�\�$�I R�ر��Fݥ��V�uZ&�pT�g��md=�ni�s�p�'�"����7n�\f �0Ի����������6��(Wv�i;n���5;[�d��d�[�ct�1�]�/c����v|��h1�Sh� ��t:�ݐ��c����Szۀ�(���l�����z���򭲦m�}99$��N���Z�s�,g�pMӅ�R��]�\�c�AP�QHA $@�D�Ua�c5a.���D.���չ+۱ۚ�+��w����z��يtԛ��}�r��I4:������~�~� �������N�d�`gN���N�����W���;�������n��>��s�ֵ��j�V�c�"�G�>z����n��7v��6#�J�VIʨ"�ns��o�9>o��{S�v�i?�����fj�G�	�:���{V`�h�?{U�%h�����e�%tv:�!7���N��7k���Ȃr<J��g��%���u��}>.������d��W�|���FH}�^� 5��$���5��������ig*��a@(Yr^$�Q�$X��	���	wr�j[��!��]��((H��V�H��ē݅�͸�D6� �V�D��Z4��	kX��l��s�]��~M�gl��EU"JtI�&� �<l}��p��l?�y8z�28�n��*欹�����j`	+g@��گ���΀��dH���wW55y�n�>G9�}^���<ݳ�g�՘��s��A�D���)�M
�%��t�N-Z��t��J��qe����X�5�z��F(���� �}���V���{V`�xl��<xF�U"����8ٓ��{V`�h�p���^>r"dq�o�T�_����=i������ʏ��M�%�D�f|5_nk���H}��Y�$F�_��+�m�`�l�BO\+`��`�\����e����w�U�ҥ
WH?���O��xD����r�� `g��`�CN!�S�q`�~�a`��|�(B�b��&�@�,c@��?DT#)#�i����O�n/[��	
$��9�^:� ���Ǆ	��Y�������{ h{ �bѷ9�{%߷:���ЄJ$��{)7�t�Q�B8lo���LI
�AvV� p𸮄���Xi�>�� �?�/z.+�����g��+�\�"����pt%�|�k���@�l����AbJ0�X����ЫX���BՆ�^�ƌ�ά/���%��P���6c2���/ޒ�B�xxa�s�KJ#�/��S@�`Mz�$��!��ܤr'`A	ڃ�~ܺ�OL��}�����~ �ICXY�cϳey��N���a���>:�
	�� �N��O��l�l����p�'l8�]&�OG�T��ݥ����hS){�V8�ͼ�"��b�u��bp;�D:�E��궽8t��d�d`�	H!��֚z�0k���z���:���8鷂�QÄ��=M�����p�z�;�SGS���Sn{�����% a � "�
}5\�u�I7���2N��x�)֥i�ܜ�~KI�f�l<�zp�&$���=� 5g�$ߩJ�Q*swg@S�J��y>� z��۶���x��yJ���S��JH�F<���\If�͵A�UW���k���#��O���w�eq"8蕺�s�}y0�ܼ� �����}̜�Uu�4:�ۨ� �;��Ȓ�t+[��K���Lh+TԂnIRG'8�Ɇ����NI&���[י�p�5Vj��m���"]-n��l��V`\.�D����zm����:�f������?UB"�t�
! $��lE=n��swW���"m�����\�BX����a��UWai�Q����`�" "�+��~��l=�OB��2>M�s�w�0�ܼ� ��0�﹓�l�z7^*�Tl"$(UTPDqQ�z��w.ç�B��{#��Fȯ
ݱ�V'���MED9���{����`c��N���`u,�Ʃ7Z��rs�}�h눎L�|���[:���|�kM�]�ĩ��J�D�u!�<����n�:8�92�'���t�^)���n��.�w}�>K��Ry�}�h�����;�YYMȊn�����۫0�G#�u��&� �v���l� A��������nzbFϗEƚ4�$kt��y|��$�I$�吹d f�Rt'v�d���k��v|�ְm��O�}�����\4��ٜ��sd�ע�k^�M6�M��WS3����	�L�A'r�k�q�Z�9�[2�v@�s�ic��FF�n�o�^AXxtx..�$|]ly�#���dӇ��ی����/�EA֓�x'!�w!�8ܗf�S��=n�&vn�=�WD�Y.bb��V��o{�n�?k�t�.0�Ocn1�ןF�w�v6��C�M�9��N&!V3k;6e(�䪒9?p������̜빇����s�b�U��I�H��l?jW�92y+g@z����G_#�&��?5�4���#�������`gn�<���s'������ Ļl����j�:��z�� ԭ�Oڕ�8����lK�k�j��Ri�ܜ���t�:Z����t�0��5;?�NW���[E��p�y�)*�Gs(�͡�.��7�*;��rL���[���kw�|���/-X��r>�I[:Y�<�:N ��V�M��W�i`�Д�	R��tH@�I	�'Ƞ�����)�@�ṅA���1DE$��^<���g@S�J��Dɻ-ڥN(�u��`z��� ����&�����=��=��:Յ,��RrUI�`>r"%��t>M� �j������?�r��6Qwug@ڗp�s�=I� ��:�F�S5YOͭ�r=���)�<���7^I�Q���f��yf8�E`RQJ��#�v�~�Nz���-�8�2Aϓw�4�����5R��`gn���l��x��o� ����L�!��sD�.��nNp{'����̜7�LJ�F������0�ʲa
D�R�I�cS)�#PA;��7y�}���jIv�*yR�V�Pu!��ZI������w��,�|��Y�>U-0*��
���w��Z��>s����V΁��̜,�ƤrP�	�ZrB���%˧^3M�dEXL��.s2��15^`fY炥T⚧Q�rM��n��� �o3~�I/�������K�5
NJ�D���mq���S}�Ӿ���Vc�&Er��6E]�Ug@>��pV����ϵ'�j��6#�J�D�Y]D������q-�}ړ�+�l2��h]F�R��|	��C8�oa!0V�q0DM��KZ�[���K����ԒI6��Y�>6�� �S}��U�s�-����ζ����7�eX�[�5�1�u��+`���9�.����g2�$"t�w�u�����V΀g�.�Z��}�՘ �Z����%j%��s��� fZ����V`	m��|�}��
���(����� ���{uf92ڶt��{|���dE:Q�u�I����{��l�>ԯ ����!EER��wUtM^`v��s���� ���>��s�Uh�#N.��S��iuC���.薘�Ňф��6^�����p J��� )d����sv���vn��8����䃧r�r�5u�K�k���ly�u�ћ��-��ڲ1��7v��v�^�7R�5��A�5r��-�k��3�cU�ص�Rs���wa���+�@���ı��[�����8��ů�{v�n��~4u��N�"����Fwm�
�7No�Sj4�hy	z���Z�L����{�{���D! ���*�&*QW����s����qi���k��)kn;׌V�;<�<���h�
B� �*�J�~ٟ� �����V~9�A�l�
#�.a�1d6M��{}� ^J��'�'��l�}���-6bY��P��AMJrG�;i<�<����"93��n�����(�"��i��Np<���7�`|�=�o�)�>G'ړ� 8�
"f]��r�,��:O�+�!m�8�'���6���}���W�!m�4ǽD&���4�g��n՞�Lb�;��7p��Fd�mr�L_?}��c�0**%nI��~�6ݻ�p��<�Z�|�=��-Z��EM���#��6ݻ�rկ�'gD�4�H6���6�mhѠ�i=$7��+wD��J�ً�����-ղe �0�\)K����θ^�jU��5�v�Qhԡ�8 n"!�/��� 9~n��u�&G��(��vEA7wWD�� Ҷt�ԯ�L�v΁����a���TH�T6�d����>�՘%��t�Y�� �&�r�}�yZ:�I��+g@�̜ _e��F$�e&ION1�=m�+��I�� g&�>����D�.�׊�Ot�����U!�>��� �����̟/k]�������ǄRuB�8�I�wwg�ݼ�h�n�� �7�D��D��6˼���&+��q4$�1JEWj8��o|��B�k;�1���5W2��̲v`T���ih�˝�8��6ْ��c�0����ڻ�p��t�uf����e�f�WUedTۈ��:�n��>���wm �j]�>J��y73Q31��q�yT5'�'^����]Vn�vc:ѫ�%��f�{S��g!є�ЭS����������2}�^�V����V`��E	�"���UC`q��'<��g}��`v�=�ws���~���pq���<��t�uf��ԭ� �&��bWn*)��(MA�E��}��}�/2x�wy����)�V��T�il�܃u�=�D^��w&d�N��zI�
AԜ���l;���>�ͭ����8�����cty�R�A�T��6��VP��ꞷI�U�9m�bpb�������&i��D�u!�>y���^f���wV8������yT���j����⋾��o �R�u�"&O$�`���c�̜�I�ժ~�M�'%Ju9��I���GG�93����M�:��j�T�q�IC�����o����7xڗc���� ZC"�DM�YwUg@��J��DG�y�O0����i'Y�m���a�	�eA	�e|�,���Yñ�����M���i"�kX�_Gժ@���JP��b��Hj��L��5�]Vj���-}� �_�L>�hu/mjkpD4�'0T�FH�C�Mŵ��|�o�F�r�`���$
�4\�v�m�0n��ʎ�X}>J���~���ܾ�u`4τ�
J;��*������Yn����P�t������$*�[�VB��vo�;����9�zݎ;����z�v�owv�|y��`�{F�x�? G���v,�~pI��N��41}Mh1�����PKbz��ǼO��`�.ROѶ&so�gO���s �(9�Q٤�9���K�4�$^�I�p�C�6bQ��*b7�{p�2����`��F�,��Lx ��u��|٭ ��r�W�g�FA	�خk��|Eh��	�=u��6�C��ؐ����n��>�N����b��H��=��o]��v>N�1�0�&�uf�gw=
3K��~w���3`X�?#�- �d��Yބ1�O��J?|~-|��� P�D���~59�����FC;A(/⠺K~E�?����΃�UfׁJ�HQ ~���\.�g%�:b�٪%՗d��1 ��aP.�W^��y��
c7�X�0F�l     �       q 	���� "Z ���SE         ��w�,��3ەlv�ְvNmp�zx^���c���`:�<U�I�y:輧OLc��g���7Tm�4���\c�$)vx-�&�XŎ�3N��WE����j�!�OJ����%��k�P=���ӻ,.��M�J����=8S�P����Gnܔ�����/���.�#&J�+�^�L�y��γ���!�'��ˮovT���ýW��l�ͣ:s��z��ζ틐;Gm���!����@ϛ�9�۫͐�0��-�W-���\���Ů�y�,M��Y���h�븙����:F�T����{z�3�gl���x�F��W��r�G�c;;i��x�[�u�!�Gm��]9�bb2#����P�
�BI(��x�z����[;�\�[����d������Ƭ/�"���/n�`�l:��#�q��٦�c�r�K1;���׎,uC��k�v��:�IsmA�v�4�3�K�<;��6�v^U�.g�˴WB��F�r�DH$u�hE�Umx�X%�;:GJ�)��by�.mi	v6�����ۧr�E��0Ό�v-����|�ͻ��[����������8��h�.:���	�E�h7V�7�l��u{m�ѸS��̄wOesdGsz�q�]��Z�"��ϞJq� z�<j9q���DƸ���[a۷�mW����xzqS)lv�ﯭ��e��A��\ku�����[pv���4�q���;O�1���^��\[��k�N��%��nktlcf-�-�W:r���d�pg��n�oe���g��v�Xr��������z=ۮ��l"�5[�`;�^6p���cg�vY�i��*Z;`븺��K�u�[e�);u/*mt<�^��]8�s��5k�p�q�v��WY���w\#��tK���q[lg�_Vp	u����nyn[���{�ﻫt
w�<�~V&s�.�a@��p�YM;��;`$�$ ��z*`�W^4�v���^�u�Ӎ�z�4P`Yh!�p�GoN�"�^@�H
�vʰ�����g]:����%ס��#]1��;�	zvt ��^�S���,;D�buE��I(��y	�:q`D)�l龣��tk�أ�fԩ���_��  �q�lTM�!�P�fj_m�i���͕�WFҲZ�:�\����]7^s�H=g��Q��������� ��1��(	������7>	��2&��ڻ��tz�wS8�흶�kn1D��]j�\^���6���[u�q���K�yՃOZ�#Q�y����=�3��B[vd�z�Ϟ6�ky���z,�m<K!l���ى���s�ݷ{�����*�k'��׭&{sv�r���[/Dv/%�iLrH��Ŵ�N.�{���vر�v�xj��>�՘�m'u+�Wn*)��(MAԆ�����D��y���I��>�h��&G�CL�QUSLY5w��l�;�^"g��:�3��]�j�<�JP5���w�0��t�uf���������j��d��E�jﷀ|���8�O�I[6˼��kK��:H�S\hUN*�VKj۶��7���'|��Z��[u�2�Lc�uϳn�q���&ӊ��NB7P������� �Ի��>��v΁�l�&d�A%���ʼkRN����1�Z���B�>�n-F�)�K�ZHF�\���g}<l��9�%�ٖ/
x�8�T�J�l����GG>I<�5+g@�|G�
f�U�s9��o�9���{Ry�{v��q��'����!)�����&��`}ۼ� ���`q��' ��1�-k=�eW���4�L�P������b�D���'��lk���LK6��-������#B��>�̞6o2p����÷��p+��BO�ƨ5M����J��#�#�l�Ԟ`v���<���4���S(�rM����>��sS'�P����_*j�DY*#�$��Ʈ�UFb��_K�e@�_4�f3��T.n艻Ĉ`A;��6߻y���O2&�GR�@���>����m �j]�7���>^��t�@�%�8r��ִ�����]��}��0l��E���YS �u�5�n�v�qJ�/Q�m��ԝ�	_Z{)u�H	���h�'$*���=���t�uc�G9��CZ�t����d��_o��o�)�L�I<�5���wy��ִ�o�{TW�Rz�ԧ%�@�I��Z���L�)7x�nzt�e�:t�AԜ�y%�;�o���{�}�I;���2lپ��]�,"U"�11��&BI��1HQWT�� �aI/��sRH���R�w��n��;�^ ��-}f���s��_e��'��P�M�5���u���E��T�R39a��-���	q,2��h�h�n*en����O��p��<����3�� �j��n2��UvUs�>�՘�92kV΀|�}�7՘�夛;�l��?M
"�U�8���������Jzۺ� �x���Q�PNH:�a�?�3ޜ.��>��� �U������nPh�8�&�� �RS�r9I?��NzN�W�w�[4��:0z�s��Zu��#���=;[�>�� 8�9L������H�,����gj�)�س�I◞�4�Pq���\bC�8�L�q�"�&^8�b=lc�`��1"C�g���8�N��ݬ�Zk����'M��d��m�p[��g�c68v�W\��F��r��9`׮���-��ޝ��flɫq�r�]v$n%.-�����<�9S���zN �z1uj۰���'���m���x>�8�Ļ�o�E=v�nw��,�H�۷�X k"r%v��Ov\TIJ�jR�������ʼ{��2~־a�Y�/K��y��t�hPu/0�j����&��-��}��1̄Cp−���Prɫ���7�}Z����$�`t�����&`���%���{���Z�΁���Z����7�g��j�?z&�E#$�I����s�v���7���G@H=�t��-�i��[�9c��"�/GZ�ع&5��ָk6T��px�n�t���֩�n����C�#$<�y�uY�y�DNi��:�`���?㯖a��W~�Ih��E���j����%�-Q����w�nj�3b��lZ<��m��/{V`mj����<C\ssS<*ɹʾ�{�y+g\���>�L�Rs��=��J��FJT�AMB���Ϲ���<�9�n���΁��8N�U5Ws�Wy�}��z�'���w3�[��p�y�$Ъ����2uէ�ۭ������7Wufޮ��0��Ĭ�&;�(�L*IJ�PrG�]�o�}w�[��X�HyRs�<�I���Aи�(���������rd�I�䭝 ͼ���I�ժ�z*���J�HG*-����8�s���B�M!4i��U�C4[��8�HQP��m=$e	g+ɝ��O�ke.����E����>��n��H�FL:V`
�E��D�$OI����ԓ��l���7���������Z�}�ߎ�|�}�>�]����$��=2���hj9(���9w�����qp�O0��O@|��!ks5ET��&�&���x��%��a�dƶ回����g�Q�<;L`�qCLN
9T��77���g���v� �kT��FH$�p��P�j
�"�eU\t�uf>Dɪ���|�}�>Իs'���;�MQUe��Wy�j����p�.�@�wV`F�آ&
W1!�&�΃�9ș�&��y;g@�w}�Id>(�$��ywZ��@H���kb��$��Ӗ��Ws��ꐷ%���{�}�����I���9�.�7�<����5#��(M�Ө��β�\�<t%�Z#C:t���C�Y�l�^t3qĩUTP�R�#���w3=�۹��3u.�s��Cʛ���"&yT�⪮h���=�h�n���V����Vg��&�Vx�u@��)G%P��~���Z:8�L�jy�jV΁���B&Ӥ�A�ʛ�� ��a�>��s�v�a�����~��%��ҩ�U:��o�f ����`*�� �+G@P%�V���cР!����[��H �l�2 �uۧ��q�V�[[���`��ϰ��뎼v�g��{EۋZ.��>�PյzgCsY@,;Of=m�>;mեT6�F�
"�t��
��
��F����t��/����}�d��ڋ���[�A��[�F�����ږ��zCGi�,R�L��b�x�&����]{n��\]2g��6`�Z�L\g���8(Ҙ������a�5�������L��{��ݟf7�
2��s��m�=nڷ�#^T.��H.�ݩ�j)Q����:�� ��-g�g@��%x�Z:��Y�	F�0VF�jHl;�d��-kM�~�6r���˘l�W�5��-����u&��V����V`�3�[:ҵ���S��rGH���8ִ�����kV΁�^J��t��M&yT������� ��G@���8�Z:���p����n�o�1��N��*s��m�N��4烦χ�-Ι���=d��k��k:y�U��rQU��W��~�f��������w.a�/^x�� ��!Rrm�I�{���dC�+ϴ`\Dw�F�>�a>�J�53aL�����^���P̲	��0!eBA�a�3��`�t�m)��BSqC�����*��΁��� [���"g�+np���>�B�������ɻ��q�D��΁���8�tr}����(�&vD�.f�΁�m�8��� ��y�-�G@|�֓�������f&C^�ruÝ4ݐ. �/V��ru8א�y�L��=7Hn��i�mDED�[����>�f �m#�!���8��*w3sS)ʕC`}��s�e��`s뙏�gk1��&���<7��B���tUNpfO�\�|���*]Tm�7kkKl+
A
�n�����_�g�,)E���\K�ݹi �@ ��B�c����_�$ń4rƷ`�JRi�6Ʉ�s�|�4���bd�t$�3��C0ݵ	,n��Xxo������-���=���y	���� �_a����濦\���Z�w��{zܲ��/�j���ܾ���n�1������Ћ��N�a�w���I[qf!#&��L�c
����e��|}M$�a�ilKg�A��VD'�SĒGѦ~�.@rd7���1|�)]_l���H���@�YQ�"ax�٦q�O�� �G'h��T++6�lM#�!%��+ģ.�G}�s��X	.�P���>�(cKo;���~�	�����cR)D�8A�+��#`n�L�ά�(��9t�Bh�uv�tzh{�ܽ㤛˴�n����+^��	R�q�b��@�w����܈<��ܳ�)_>ց3�$~�D@�;x���c����+|8�?�DX
�|�����ra�J惣j1���ZHy�{v���ؔJf!�!�h#�Ə�@X��\gs�s�B��Ӄ�ٯ9i%��v�'9X���y�"�ꬻ��ߎ]>��v�?zw��bO�p���vn@�c2i�&����`����ԗ�/:��W@�@����JUQq.�c�"�;�H+C��;���ÿ�~3q����.A��Ɓ$��S��г��ʗ�k�k�e&Zk�P��d��s��!���j&Qzmѝ	�/ �	�@�;`�4�4p1��N��v�W���8�����}�e���r�p������ ��r<�	��i��,a����/C��w/M��G��K^��l�l��@�M��N'N���a� �;q:�����8&�ʴȁ�,�s�x���x�^^s�ut�L��(Pr)Ug@϶Ҝz������0DrZ]g@�tY�Ô���UF������{��V`[h��jU���QT�\PW�h�Xpm�:YӰ�mg�E�8��7t�x��#$�2&K�KjH�'w��0���:}^J�#�H-��yrJ�D�EM�M��嶎�����7X�m����8 �b�Bh��(9!�3��U�o�)��93�jy�kV΁�V�#M�oj"*$�ɺ�{ZI'�=�;�O0-�t>D^��;Q|�!t�&�� �U0*�dp}��c�O��??��m�"�#��w�j�n�:}^J��Jz��s]��&9o(���'^�G�ٸ���7�B4���Ś��Nu� k���
7����l��y*��)q!�jy�n��kt��"�P�w2s�M����jy�-�G_&M�Ld�p����g;���i��}�Y������}>���1+�"��	NH�ZI>��� i[:O�J�s�>v��.C���'JFBT��w0����~�����>�����N3Zn��CIxK�z�D�fj�*�5DZ�Srb�*�eJ��HT�${$39t��]��g����}N�;�~���` N�9 ��i�M�3�;t񴠳qv"mۮzvy9e�	��֓C�`.	ݶ����3�;U�lBo2r�tv������m�M���<Q��[g����D/�܋]���h�X�oQ�N�5�un������ת^y��إ��&9Z�qI�Y�ci�
�neu�qm=�0f��-��;g�3v���-DF6m�q9�i������o{om��0;�+�kۂ7��\�p�K\�7.wX'�Y-���҃��F�:��ꔜ�9h���}���N򤧠}��g�9�J��+3��f�ڈ��*�6��Y�~KI-6{ڞ`	+g@ϽiN8�Dɱ�J��LJ��!*8�����.�a��I��v��t����DLO*�u5sU5y��%�t����*Jz}�O�t�y�Ҩ�M:��J�l}٘�����N�$� ��G@|�`�4ɻ�f�b�ï�Eݨ��{��7+gy�0u��P�ZL�D1�]UJ�)9Z�IM����������՘��H}��� ����AQd�UE�>��9�{��4���'�� Kf��ۘZ�UI_Xk�5E��U��-�%񤐄�a�za�>���|���ߴ��ׄ<^��d$��3'�����8>DL�����O0#T%'L�Q7$6;٘�ٙ��>��3Ĥ�΀�����bਢ��>Iv:�n��7v��3޴� q�����e�~�ܽ9&n
����mG�?m��~b��̚k�ܗ\�#����U�Я\��ʋ�.����ۘlw�1�I%��=��;�l��V���Q�UNp�^=��L�n�s�n���}��s���̆��Q*C�:�:�`}w=��;�ͭ�,Ot�(�J��0�aF��w���ʪj���e{;�gzԓ~�z�$۸�f6��:�Srrm��3k`}��s�w���ZZ]��|�f8��t�P�.&��}���ޤ��g�iN�%��Y�c*��U���D��*h�"��أ�ˌm�k���mҖ��j�����u���d$��y��٘�ٓ$�ý�{� K<��TB��G�;��)��r"d�v΁�4� ��G\DL����4�ڈj����������ً0q�D�J��7vۜ��Wq4Y5Qq5W53Vt#��6��V΁��iV���5l� �$I*��)ʧ�EQP�!$$����yd9eo�E�Q���_ Ai|���>�4+� E�F@$S����&���EPVU5#��UNp��l-%۽���<ݳ�}����by1E���\L�7^}��Ɇ�N�kl!9M�v��v��'Zvr�ӆ��5*��Rr���� ���>�d�`}�fs�]��`}��k1�4T�����p��u�d��y�$�����<�M�J��/GH�	�:������ ��GGȉ��}f���� ��4Eܖ]���G%%�t�}f�S��ٙ� %x��2�5M���yu�"9����m���G@p��$��i(�	T�)�DDz��� �-�4Q,s��J A%U�$�щRʄ�$a�.�^(�����Ӥ��  xر���u�l�f�s�.�\\�k�nl�Z�ی`�^NI��:m���8�9�Q��Ƹg��`̭��FU�*/l�;1�����c��t�[ֻa��a�����nݥ.e��m��l�[��ꬉ�����N�kY�w6 �ng�m������3�m��G8����&�۳�Z^�����t����y�����gnml�&��"+���W�����m���윟��b�:�u����
��O��]��&5�΅��,R���z��j�[��/=?�3��s�aw~ߎj�{�'DR���7Vt�If>rdI[: �+G\Bl��~i����R9:�������yu8��7l�z�`�	Lv��*.���f���>D������:��g �����_Z�n�*HT�N.�V���z�� ��t����9�s����<��X�ݢ��t̽n���vP�t��m���#r%v�DGp�g�־5Wf��������Y#�?O���<�@5�RNp��m����Sf�V�Q� .J����9�GI]}�{���>^K1󜉐�N����(��Ws�<���ڭ��_��y����J��z��jw]����΁�&� ���#���s� �t{ғ�J�%F��l���`��K��=���yZ:�q�S�t��j^(83�����ڛqttv�]<"O�t�=�h8�wOn��UU��+g@��]F ����-o8�^�[�QH�S���T6�����"dz��[�mj�����R���]@wEU��L�t��f
#�^F��H� 9��"�21"�J����G�D��Csi�.�L�l�.�KP$�i�_u��=�8��dXB�JQ�WgA�"}���J��>��Q�㜗�~6q��UCl�P�Np��l�n�g�=v΁�ږ`��[��⽸P�v�&��7�u���N�q4W����F�[�Y[cs$�p�vƴ�u�o�Ƿ_Y�/+G@��K"9�J���y��=n&� �og ���~�ִ�=��`+g@��]���D���	]D�WWuWWQsVt�o0�h��Uj]�l�L6>�v�C�cB�T*��8�KK���}���m�К��}��i�XF3e�E�S�nI\S5<Mv��q�3CZo���a8}0	��qF1�!��F/��=�}��4�5�$�9�=��kt�����P���}�.�@߶���,��>s��������n��x�]&7�[j�t�ӵ�^�qx���c�ջ�l�n�%U�� ��:-K0�h�{˱�:��dUmP�&�'R���s�M�̞6r���/�o4�}V��ScP����0���}�]���m��3�,�]����%)���y�/�[<�<���iu� �58�Qw1E�u�����K���7� �2����2L�������@ ��
  ��O�?�*����g" �'�AEDf�Q A���0��c��p��w�� �����9�����������O����?��������/�?�k � ���y��@ �_��  	?�?�?ԟ��O��s�_��'� � ���G�?d�6~�q�_�������v-TE*!H,H1Q"H AD��H�ED�1Q"�AD� �D��D� R( �H�@�TH�H�+ @� �D�H��Q ��D�!
Q �R(�Q"�ED�ED���D�Q" 1Q"��D� R
�Q"	
�D�$H�Q"�*�"(ED�AD�*Q"��
 �D� �D�)"�"! R
�D�0Q"TH�ED�$TH�DD��H Q ��Q"(�Q"�H��D�� R"�TH�@��Q *�Q" �D�
H(TH �H�� R""�H("(ED��H�! R! AD�Q"�TH�*ED�"�AH�ED��TH ED��H��D�,TH�ED��H AD��Q"�
���Q $TH)"�� �)��� �B(�,*0�"�D ��"�E�$B ��D"� �HB$B	 ��B@$@�BD# �H�"�! ��D B�
D 	�$B(A"B"�"�B*@"	 ���B �"$(,B A" D �)�	 �B$B@# �BI � ��B1E�B$��!�B1@"@"D!#�D!�A#�	 �B� @$B0I�D! ��#�a$D	�	 �D# �D�**$�������@ <rk���'����E  ��k�Ǳ�����?������ <�����?~��}@ �X(  �B�@ ~?iy�r�@ F?e���eY���?�F���,��P  �����O����� ��!�����0��1@� ���@ ���~̘����������_��k<;���?��� Mg�D�_⽾����"� �~��W����� O��������������b��L��q����� � ���fO� Õ~,       Z @   Q@4   
�}     j�� � �   �	   *��
�I   PPP*�� �� �  �  
T(  ��                `T@ �@�0�
�T�y�W�Nm^{u/�;�,���� O|)ݞ���_6����}��gT|{� }g�B�n���7]�]o��Ycm��藶xW��W�{����>����ݾ���׭����tl��ξ���z�� ��ay1_{�z|ʚ�{���|wx���{mi���|  (�   8 � h�֩��=)E��NF��R�.�E)@��)@�%�HJ ��v�ve�-  �)	N�����=� �S  )�c��Ѣ%�. ��JR��)	@��:iAH�R�.%؊R�D���4P�f�ADJR��є�>�j� �@$   R��2�@�R�6:�)u����x��˯l�� 
<�[Ნ�sﾻ���Լmw��_w� �k�*��<YW�ܾP>�T ��3�o_m_;���ϪX�;*�����W�[�`�=R�8�]�uxC�����-J����>�    Q�s�Z������aw����n��{u�yC6w�2o�wT�k���u/w�ԫ�y�UZ�ԫ;w��w��� } a��x6�7
���Gm{�N7��S��<-<l.{��8�y��U2׾���j�L���g��ʫ���5�   � @ �&��ԫu��
�g]����Լ}�/R�|xZ�=sw�K�W����+�Y���<��T��{V���̞@��B =��p��� i�ԫu��i�μYrj����җ{蘒�_>��n���_\m9iWz�G�U�     O��J���  O)%T�@h2d1Ǫ�#*��   4�j���U* �S�	SتT���C�%$D 4x�Q<}��C������3'��c�����PU_���

��QU?�

���(*��AAUb(�����?��"�?�������#�k�ʒ�k�t�}PP��PW��
0�Z�����ƅ�����@��]�T";l�h.����"{���^�?:<\LC�v���m�jկ�6�Q1�y�&�=�I<�Sb�iZv[�A�As�M���SN�\S�vghlwe�a�p��w��==�XS4��٠뻗$4�,Е0�-Peǒ^��4�9��լ��]�qO�{�<��8b�r���8�^��*��f�nv;�3�8����r�
�d�v���DW�ҳT-Υ��m�����#���ʳK����6Zx��#w�W!ՠ�2m��}5�����yLMp�hA�v�ŹL�+���@����E��y����<{{�v'e�����!�G�������}�(��&l�s�Te�Я:�܄i7F�+�B���B��s�o�A�������v14qY(�Ak��!L�sF�(�/��Al���p�^���������K@�k�̻��"�CN���:��������jͷ�6�T��ֹ��ָ�b<-��نf��Y�x�xX�n��8aǘ_jg�+�;:گb(t�oH;�=���1����=����9\
�	ǈb)J��!����b��Of��˸w�x�s�&�U��ҙ�cCQ}QE�6py�ֶ31�}wB�7s^��P��f�SsN��r͈c�׈N_\�����Fv�1ڙ7��M�wOG�ڡ=7�^yd�S�/4n�(M�kǻ��q| Y�����+�!@� 6\�����f��Ĉ@@�Pyp1��:��h��{l����nr2�\�rs��Z���è��(��]Da�8_�JÊ�c�^	�;�h/�v����%�-��m�t��ngV�"����Zg����A&TI;z�S|��`���Lvi�Pp��qQ�v�����fr`�k��	�Yş�k�!���7rj��؞���8Z���x�7u9����� ����̤0NzW�ۼ�L���   YG,��V��������:��	��^S;ġNwn�)��l��g������.K1��;��Y�G;���n%��ࠍ}�-���/h.ٻ�h�
w`jO<\�ɻ�A�-VI��Á�������@��an)1�#��F���i�1�|^���R	!u� ���q=�j��:����]	�Bc�&ƃ���l՚� � 	H���Il�!8J� �K(,4tBv���#��s��z���ͪ��x!����u��a7һ�OJ��ﶜ��\a���~c7��ܰ-�B���.���;0IV����-@�>�V
��� ї���쉡�~^���"ٹ�+k�b�7�!�Crt�"��D>C���T��x`>�'0���t��9W���W�&�e�j~x�^)�v]�~�>9"8�'֡۝�|L�ő2�]d?�7o)��:�-� ɛ��kI�uy�1��[֏c�.c�ϲ�Mƹh!y�a���eb�R��x��"	+��H#����s��Bɇ{{3j��*A"s;i8}�lxd�d��w�|�!L���tN{�]��ۇW�#7����n�������w~�`+��@��g�0���s/��sغ��p�d����EF�Dy��th�өM �3.!Ju,�p��Bc����-��0ӝ��ཌu��ٛ8f����3��NAɘP"M��=�|HC�T��� �@9.gO���h׹'�@��r�A�;��s!O����|5s*�돎v���)�&t�DD�H˙�������2h���!)���D��*F����7ZAX�d �����w1���
VTcN�p>�E�<k�x��1�e2�ކv8^vw�Z)�;r�BΧ��0i���dDy��pWA�z�c���-vd�~%{��x3�=�;8E#�r'7gv̍��:+s��j>A���3�vn�����m��w+����̈́h�Z9����gwvF�N�sm��Bn��B�A�0�,�v��ʤ��,`{��<m[u��b��8B���Z��1� �v������Q�>OHc�����p׷t�44�H�34�6�6������iU���}dr���5x�Ȗ�]^a���;E㸧9c7:�uբT�.`ݓ(ĥ��9���q�ڹk��ٚ��u����{�)��fv"�y4�#u��!���4���0Ŵl)^3��XT�L�/+���w���+�1��8<��; 9i2=�QE��R8K��O�6�é�x]�7K�c'3^�i=j{�+[���0ov_�ϰ��gњ.��^��۽�x�u�$�\5��	9�
О
�=H�\Km����{�U��Q��f�0�[Q��F�j��]��54+'5��vP�����u�� l�ui���A깑�H&�곯D��B.��e�֢S��(q�1�n*�kX�Ip7C�k`��!�����^ѶK�%#%1	!n{H^{sK�p�|NA�E�H'.�T�gg-�j�V�ۨU�p�$w �c�mW�5W�όo5�SfMm�1���2\�����8sx�%���m�aEqx�
�H8� i
�2$Na����.���A�əLPD \aP4�p� ��#��8��R�P�{cn�!$rӻ��a	�Y��N�V���z\��	���C����L���a��9��`�{��G����B�����:K�0}V����'�H/�$�Iì����,��w��P��xk���5�2=�	 ��!� ��"6����)Z$�<:�>
|� ���0��0t��M0\Ğ�|k�r�~](�a���3C9ûΓ��;�d����0c,�{ìtmOs�ta�v�!�t��(."y�k�7Sy�Ը*�������~��Gp�j�3���Ke����$���d,�q�h+����k�'Z��$H���=/c��?yvZ4V��&sKF�\)����t�#r���y3XRx���8p���e�ѺVd�g,�@�x�
[��f��#*�1�Ø/y,p�퀢AI$I/Q�3s�-�hc�`��{�s���TM�ǂ`g�h;��(��>�:��2l}ؠLk��y]A1p�<.���1 �ň!� �B4lz�3H���.!y���'��(�Kw^�8�$��$p�j�OU�.+V����Y�����v.�sP�N+���:�+��'p�Ϭ�j3�����fv�76��<O�3 �F���{e�\]��A�ՙ�nʳ�7'%���פ��b*�K�%�e���|�(\7��:�9#[�v1N�[�of�8�W��Buj�m������y����:��Ȣ}C)�.ݿG�,��1���� ���T�9���z�ϞųgW�=���`Fp�!W�w�f����
<v�S������W��A��ɂ��^������Q�fm�W#�E�'�s�#o�����ơ�〽#{�\��@��p�/���E�e6aq�ӷ��7�ٌf��=>L�6�,��}N��f�1x��T�S�����=(}�vaF#�VB�N}6�wu_9��'f@�MB>��!0�x��w(-��h٬T�έbǺ9ܔG���p$��V{+�p�g_kn�p��ط�A���a\QD@� .Be�ډSv5i)aq�v�=���7Mw�81�nAS�i�*t������JrXBB@�aI$�q5����㉳	��V��ɳm����_q�3VQ�J�yAYv�Yk���8��6mǲSù�Yls���89��'�7 ��.�3tC��<�|	B��8��{f�1e�~�����y��G�! S�	���	*Pk)��(.���j�\�0"|�cÂ�J�S�7�%��œD��ȨRY�<�Nn���tɃv��W{"Μ���_.�M�z=c2q�y�����pW��P+&�D&�2��؏r���H,��Ua��G{ �x��I w'[˫:p7s��۝�S��Z1}��%�I<c��-�<�!�[�@�y�MO�.w[�4�l��)���l�U�5������EF/y��L�`�b�`&nl�{a�c�ݦh;!��Ug� �΢=̫3�c1�/Wřo�� �&�ۉFk왉��7A�w��Օ��[�\���0�[_���/`��c&���$ �Kw^�ݡ`Ϋ=�; :NY��i��۰���8:6�Ǐ�K��si)�	�*ӯ;Joi�8�o�u"��=���d��AD]�Q�p�T+��Ua�/vi���w��(�V� ��7;������A	��uK���]Ԣ�J>�s��©�|ю:�Am�Si�4a4�Aw	�(Ow<+��n,�.����<x���)�Z�x�4a�B%�;gq!�㾯��lE�MM�C VE\�"]8lbr0hoc_NO��1��6T�vc���{26�&8-Fol����ҳ��1���X׽w�GQQ7�RZ����.r�pS��z"��A�� ����?rd��ɾ֞lqe�{5�*o�ܲ��#�}ĳ��ݽ�.�����N�d��i�R�<���a	�[[�vs՜��o��I��MXK���ry�*�L�h=�L
�8GB��>;�T��ok̽���p�����V�5�6�����I�\�&r����/Ց+�`�WBDS�T��.�.B��u��N�`�f��o��0B~ �HQ���Q���W�7uvkDߤ9�qbv���X����@h�q�Sܝ�09MB�\鰓�)���OXa�;}��x��[�ͨ+���/K�̯��⦰k/36���q�Fn�E �A�ҳlm�2�ޛ�$Lc�f������SN�Ag��8ve^���.rX��""�h������1�չ�4�t��i�B ��ff�Bs��臗Z�Z���X�\��p0o��ւ!BB1	w�s,��3� �3h<r��g������ɺ0x���|����<
�0��6ڒ\�f��C3r��m�r����f����逍���mZ��g��A�sp��,�zU1S�;NQ
���ێ�{���Wg-��9���F�����qM-O'mހ��օ�
h���"X湃.���Ύf.ü�m3�|�X�u}�=�r�9�;�/�h9<���G�(�7�a�owtN	��G����\�7���.�rn�gc�ȡC� ��>�⺼�ݹ�&��&@��]��c	��7� ��C �=[;��f��=��+1cݗ3��@�T�:'���l�d8kf-.�S�˾�Ӂ+�#+�@*A���y���O��	��Uh/6���f	��k�fwOiUq$x�|�+AC��$ o\���
�bK��!y�=����W0�v�!/<C��7Qo�X&��2)ٓ5�fh����:-�Tx��)��Iɇ�|�}8g������@ ���psNj����O�e�C��F��`�g��^ͷ�&bfǎ�lC�.�B�Z�';��Ioa�����GI��[o�9.-�\9������޳ؘ˶���L�v�!c�ݰk�jOd�79�f��܂4�ぢK��h/az�C�u�g���dĐ��Nu��b�O*�%�
��oX�����p�˩|��c= ����>&o�*���NFA��`^�R�+
E0SG��8w�d��� �r �%�����M ��<m0�f�cwʱL ���zxm�<c)i�����4d[�&,�BB/u�y�%9��e�/kb(�@���]��ΰ<��2I$�@  -�                                                               �_�|��                                        ��                                 m� �                 ��                                                  ۵W^�UM,�Fe�pJ��+��bW$�܅��-R��$m4�:H��E��r���ZЖ��2�]�KWa�ئRV�jVd���Հ�;WV�c.+���Q��PYEҘm̻Y�0�c���ɒ�]��@��@׬PnVZ�D:�Q+qs�V��5������i�)�:ȱ��˲6�i��K����j��H�.��٠����Lsv���&�0ݑ.ś#m��R�(��3��7�/jE�۔�{�X�i�mڇY�k��={E�tٸ�{v��NYv�h�*]N�U��6a5����꘼	r;i��j�k��j�]7l���K�6�K,Y��k5��&�f�c��qH���#e���1Ԇ�[*5cRdq*�eIm�v��h��>Up�h�n�h�M�i������Lf�nc�k�BT���f.�4�3�S�e��
M��mf��f�ʅ���J�1tp�2����qn{�e��%P9�)q4��|�6�B�K�Xgl��	B�u&�Q��Y�%�\�MR��jM��4�L��LBݶr�uv��BV�Se@ٚ��e�;3BĮᙔלW��52�6Gamn`�,�mv�ָ]�)��W�J@�i�C�bW#ti�h�x�[���pg��%��6:/+I�.l�m�n���ۡ�m��T�6�$J7+0U�M�́r͂]���э�m!l���sLQ�	F��]me��ы]2s�s���o[Z�Yl&����;P͡�ipi�!n��.�Z�KQ�hLJ��ie��n�f���V�'Uå�t.҆ͅWmjGL��D�͌2�i[��*�p�B�Ԇe.��k�7m!�i{[j�Ȳ���"g �b�lZU&5�\�k�nHj]�x���T��}a�K�sn���b-
�%����룘��U�LB�SYJy�,����jZm�m@����hW3����%�k�-6�.�Sb�ʅ)pM�J&)���M1���l�@z��%�q�J���K�C,�v�h����I��m�&5,R�0m���efv��g��4�I`bWPW �v�R��vU	�(�Y��Q�����Ҵ012Wil�ݼ�Ŷ�l�:�Ԩ&�CX�6M6�]��V��mpG�6�V�]Hgl8�Śv�gRv���pPB�Ll]�Qv[��xjCRS��6�\X������;1�z^�V��Man��6���a� I��6u儜��I���Q6�Y�9�ӌp2���[Ĺ�����in��z����� �Z����]��w٢��"���m�m���TF���"��Z��,��B�2jf�ķ(�&�:�;v��m����$I6��mw+9Jk�I���bv��m�b�:���b͛J̫�e���YYA�)i#]�vݭ�$���H�RW4�s�+U�9�����)Wv�-uԚ]T0�H�Z�Q�gR�����k[a�m��nz�9��ؤ!4*7b�*ˠ$���.�<��|lt�����[J��$��%�\i�1--�;Y�˙�l�in���s�۬�ki���eȋ.M�Mnqd�6��-sn̍�kaf�q6�5�ܗsGkۢ��cv����f�T»#�Q��:3�b+-�&�H��ZX�ZZ٭M���1�6ph�ۈM�u�0���� U	`���u�݊E���t�%���4Y�9�3E�1�S:�I�m#n��e��,ί���+�v���p(P�ꨱ!���܂�7jit�f֐4]��d*���lln.4F��,J��\j�Su4K�P�hb�s�i��3/e��Q�$�6�K#����X,Y�-���ڋM�Y�\[`gLjJf^�  JeMz�CI�Ύ-��R㍶�\&j��F 1ssR���� �0�\�6c���/;GY2�{&��۳�zM�����nZ��6���([��&f+ɮ�YM�m�Il!���Ye����]3�B.e��/1�E�X����cA��tԛLZ�05�Z��8��M5���ת]�K�$�:K�)�]յ[����"l�:1vf�Bb6��:�l�/y<-�]��f��^�f�f�q��Q�����e%�Vf�nK��ѡ�aT�K�V��뭴���!��۝�L�/3��,���%XKٯE��9��u�b�l��c(la�$F�ƶ�l�׵���
�-����su�fba�	p0ы�GJ��MG6:�M-�.1�cT�5�6[����f쏊ШRS����h�[kӵ�v EK�\�cj�5�� �&��Ѷ鳛1��a֫s\PQ,n��V۩vW(2�؀ɭ�j7Jպ��S	ja�ԙ�]j�J��M�*������]f�a��*$��`�Y���٘h�-6u�G� ��T�k�cE�ŉ*0�v�p4F3U�gF���b��ˎT@]X:\\����#j���h��C-bq����%�A���ShB7c\`��\!MK�Lmp0%U��k6)���@��͓829�aX�l��uWHfF��a�0�abAM�J�
D�⻠ �l%4���&�d���sI$���nVɳ �����:�[^
�e�h�t� 7�@��Yr�,mL�\��E�u��m�����(���g3t6lK(����WY�D�c�q+h�0ܜ��!�],�3tB\V�M�]����f�m�@Λ2<�hˑ��'Z�� n���h�)�����
�����1�Ĭ#���<B�B袁������aQ�v����e�/4��]�֖��m�A�`�h׭�b���Wi�*:]����۝�Xj��.���f��Y[�b�Բ��fH͖X��X� η&0�P�7S;m3z�5�R
M�
>�n*ʅ
��V�[J�v��h�l�e�k�6�b���j5�v���.��X�"��V0tx����k �	s��5(��ԭ���m�[�L�պJ����s���e%�L)m�՘�j5�	7&�Q�]�-������z�7	H�%��;pR� EF-�a�5�f΂0+Aͻ$ك�l"���c3A�XB��YV��$�t��헫mmȧ6�6�tg�A#���F�䫘���t��b%6f�6�˖�L���Q��]�s�����@ d��2@�	�cR���ְ#lI��9��#�)�GM.Z���i�XS[�Ik��1Jm�&td�݉���^����t	Un��&�Q���LM]
�`&ζ�1�e��\���f@.�@e�&N.��L:WYZ�mi�H��M��,Ʉд��H���d�gn�q�GZ�cKcuy+���֪XL�&��B�b�����Bĺ���l�; �-�����F���)+K��p��CT)�SS'Svŕu�v&vH�S6�m�Ί���4-�˥�v���*i��I�D���5�+c����O5>y�y�.@^�Ե*�v&J�m�C��m�t��K!��4�+GcDH�@���X�u��5��L�K�h�X�;C��4�����{I]���kK����i�umScW��,�/-m�r��a�f�nvo�kt�'��̺l��P�1�4��(��V�]��jMmL:����8�݁�q.f5�(X�s%�F9�nƶ�6n�BЮ6�T���Lkuƫl�j���k��+J;K��i761CZJ��"q�g$��u�atWA�GI�l�++�vΔ�Jy��
u��Ⴢk�f�+���l���0��-�`3Q���]w-!5��l+4�4L�K�Ú�ph��2��.5�����I������Z��c\"�F%�/*Ei�;J�E�Xk���m��ׂV
��q6)��L$�.��֙�֪%D6�L�a���Ў�6kH�!(�V-�bԱ��^
eHi^�ڈ�C�ܤ�M��m�E��Yz���i�iv˺�6�\gm�n�����6Z������$P/kn�(`Hc ���e�=j݉�X���.8)VRQ��6�����f�֏��w��&���� ;�
ѳj"dhl�-���n��iM�탁{]Zޞ���RR&d��Blڬ�鱴�tכH6דn�A���l$�,:�%���^�V�n
bj�aw�&thE�ŕ�0�R�Leb��*�K�j�V�n�ˉ�İ�C:�tݹ���]�&�����l�V��)a\`3�e��m�I�]�nLmn*i���f�m
�%Ѹ
�-ß7f�l�2�S��.���t-S30f1�RXmy)���!�`me�Y�-�.�tU�2$�":{5&�l\��.,-͚]D�&a�&4!em6�;m���-���؆F[i�]Ś��tD��y�Y|�	\l�fٰt��
��Wm�n-�+����k�s*�n��U]��J$� �۶HX`� Mt����˨�\T�k�u����9�5]�r��a�-6�%�*J��6J���5��-���ms-��Y�����Yb�D�T�k��J4M7[l8�L�u����e�ԃ�Z�kuc�pG����X]��2���@���.�;����u/]z+�S��%��K5�RQ&J�8�lVc[����7��/�]G``a�hj@�$i�(�s�% �j�ː%�Y��R���m+WP]��R�iD�v��܉��r��!ȵ6���H��Q�"Q�h�vaf7R�3\!4*lй٦lɬ�cJ��(\�ֹ%�g˯����Y��hڰ�H�N�o\�%��5��Ƿv��-�h���ۊ[إ�4SQ
k�[5�0;LL���&��)<�f�fƌ͕цbE��̘�d�3&1����"
*�����zɏ�Ith���B�~�p7O2��`;�ӓYI@	H1!�0�6��1K��#$$rآT5o$,P����=D�d������΀2���`H�
�qx�&��㧖���V�C��	��` dɈ$�$H�DbH8v���r+ʵ�
�2�E�����H�Cwɂ;�h�K��G�U�N8���d��Ǎ�2H�_p
x6a�#	��@���;$P�8M�S�1M��%0)
evI �l!��<��:�
m#�$<�N2��d|�VYKHL5,*o������!��3�0"�:ቹa��bHl��C��
���y1呄1/�T�@�|:5BHP���$��lؘ<��xe:�#$ �A ���id�M; �~!�.�w�n�!��҆^���;������H!j��� �RBa3�	*��L�%���P����` H:X��Cia"I9�bEF�Ԅ�&��u�bB�I4R�uÔz80	@�W!�8a�L&��ǉM.�@aD쉺��07�w��Ȁm[:V=Y���$2�|�L�q0&�b' vu�8�C�	9Ęp�D�z2@��9 q�NfG*=<�9v	�N'B) &�8t�b�2I���/3�ؐ#qX<Ն^�s!�ũ-]��D�K@I#]Dppq3L��șV�G����K#I�A�9��M��0�H�fO�u��$�@ >��5��Q}А�Ѱ1C�
�
X���4t�D���C�r$�'����Ĥ �8��;J��&���u, �� ��EV$PpFa_�d`(��(B+�8d�f�3N�]�3
�4=)$���uC'��.�@�!�C�c!��A:���1J@�*��	f����� �2��S�P�$"Nu��'A�$!�A��Fbn�RAC[��$�$�N�! FsR.�.@��zۣ%]�<D��=���Z�bH��!��F@�l�s�,��wp3�a�`3tۑ�A�8I*`<f]i"�3�A��oc�9���@9�Z=��iBI���,$r�tC'��	�J�`��2�^S��f0�j y'��V��"�RAӳ`e�`FE���0��p�!�B��� `���D4吐8�,b�2��d6I�w9l#$q��$B�W��x cp"odH���T�!M�5I0s�c��0� �A�6u�`VD���hȩ曞Ȍ�DL���4FA�Ń�z��(ǖǐ1$8<��I
28}"����Xj/d|�Z���"�!T����`F!!���'2��: d�m	5a#C
�l&�R�hRy�i�����Y����W��"�ΐ�� �1�\�,���y��X���z�"2@7�[J��)$��NȯJ1��rI�+��׾��!�$��I�BdA0`Ca�N����"x`Q�!��h��4b�x@��m�@����6���t��*a���Q�ф<�L�"�D�ģ�HN�I!�2#��T��e!!$� �I���Hr�dM����p��
�i�<�dxZ1��uő���!���~Hm�a,O	�/@��'��e4��l{�ƀE�B)u@�憄Ύ�Ӵ�w	����u��@��"	��h�$z��Ր�'i![�ȃ#_9L wpB
q4��P�:$0-62*� F�n6I&㢞P�n"IRPz�,"�bB�N���&P�T��4d#�Jc!9$(Z[�T�BC�hzHq���R�	$��Ғ���M���N���@Hk!,�-G@�]� H��u,�g�2ĝt@`�0 H�D�fL02�#�7�8>~%CQPٲ��v���>@�8B$3���D2l,�$':��ӈM>`j1�Z�3���C��`'9��͠p8D��d���)�$!�Ί�Sa@�>{�紋�Ia1(���k.(bWAԽ\Xj�eޢn���q|<Cϯ���HGM������� v!l��JE$#@�ܧ�(��	�d�F�6Sɿ�!g���8H2 �KD�f@�x6@��	��H���B)�;����B�7D��	"C!5�_L� ֱ.̇ʅ�@���B�p�Od���t#$�Г�]�������2CqH@��`:��*i�z�ș��v��{�/�(\B�4���"���'��2�D��Y�1J�@7'j"��97�Mm��^�aM\�d��.KGY��!$�@a_:vf$�N�#ټU�I 
�0u�E��!ȆH]�p��8D$��FA��p�"�RpD�d6�JeaN!y�J���M$T�!T8��Am�-��\��z�	���@f�I`B0��|�Jl0��.ӶI"Fp9A!�.�Ht�8��[䆙"hS"<�ʐ�q,��"m�n,��9���I<X�G#d�BNF`�B/3��y<�̇�N_mX��,��;�'��$=��i�Go53j������(�q�4�����$�K;������x��*��          �       6�         �`         .�m+��n�4擳��T.wQSU�K���p@�vn�E�.��-�ka����:!@GRQI�&`F�]-�R!�ǵ:j�&�k&Ɲ##]"V�����z�2/)in���s��-3�.d�6�9�v�-����-��4�vњ]4�ضk�`�����b\��V%-l�2��M(bb��M���L6��V�E�Ї%h���-�3V��U����t�����&�.����]Ά���h��v���+�Lic������Z�Yz�z��y)�,e� �
��fٶ(�j�h�v-����/N�b"3dYժ���鱉�QЙ� ��k��8�śh�L��hMe��0+c	]�/)l�L�!��k��`�30\�v����	�XgKńu�Kc�nte�aX���L6�"Y]u��er�ˋ4)-�㝘�k�s��	��]�ŠmU�����m�X�t�9���]��/%ٻ;sv�	�9�M�h�b��Vӷ)f�X��6�L\ˈVkoi���B]�;W��r���Z[eY��,�R)Q�kys`2bJ�XU���qf����R8�[.l�\��n���k-��s���	�k2홥��3��[��;2�vILX[� T��W��`5��������$�����aZ7�w%�ö뙺s���NxZe�%�7mt�a�L��]-�ͨ#p�:��fpi��\�]�n@�0�`p;m`�F�ꅖ���9җX�W�b�3lY^�q&�N��]�Ck�����QXB��F�dcYr%H�Z�FX�Ã�u����լ(Fg���.��¹d�meь�k��+s.���Z�%�k��3e����͵nÙB�y!����X��Y3X�iv��X��J�mJ����nt���5�� ��&hܔX[����K��Q�#�m�ᬚB��`X�Z�8��l�FF���Űخvفr�HЕl��pLg/���l�~ ��|oeH14���`t#��规���y��8x<�&�w���b�E���tC�B�L�_�z��� k�T���]�����K�GN�� y���z&�צE4�8��m=����㮎��H���h��;;�M���c@d�p'��;6>��0)�$�a����yp&�<���ͧCX������߽ޞﭷ� m 6�6�6m� K���b���땛k1*W2�R���`�J6nbn@�����/WK���Mn�3%1���2�,u(�&���p+�.���Tc�f4&XҰslKe�
�Vv�6�]m2��Ҫh�!��Xj�Z�j�v�Zm;2&:t�Xݻn ����00��f��s��`�.�nWF� �mn��3�-����/Y-�e�-��C�||���ش�j[6���m.�b]N���뱌H@uJ�h)6��P�N�q�ۻ,�j(pͫ ��V�r�
]LTUD���rX�v���U_$�����`��|��S��"))$� �>� ��Vw��{���22uk�BRT��Th�Xwԗ�zX�t�>�w�K���|��RD�zb��UU�n7VG�3{���9���=��`w��fE�.�(�J��T�Gs��-��]Gg4n�,J�j�6�]t�,��SsBa�td�4��''�=��V�f� ��g}_����̧��T��'DW95$��ﳭ|���en�.s��b�O6�IFA�&$n���}V����D$doR�TUIIPN���37��o�e���}I{;���w���!��aDe(�E$�脻{���7]Xw�-��`g��T�B�IR
�q�`~��Ձ�W1���7_U��[VDlu4�RJ�������� �]�үk[,�6����$�&�ʴ�Y3��v�Ӷ[�bllwԓ�Ͽ�� ��V�mw�3{�,���i(�B��D()%�{ٲ����#��+7���h�u}�z<�C��2ET�1^�� ���;g�XkwC�lA���Qa�L�W�҇	�X�����Ɣ2�"u�ڥm��
V�ŝ�e�o�e�n掙$�9D*$��G�>��9��`��ý腻]��ܧ��T��'DJJ��[,���Z�W�n�r�>��,��:êfrċjfL��`��]�H�ذT^k�36e�foY7�`�Գv�$����U��-��n�"=������5�L(��	�/n��<��,�_U�f���F{g�UDU9R
���`{{��kٲί�#7zX�y��Z���q	Ɣ�IV脺5�X��`<�j�>kI@��c����,�o�g�y���05> �i�	�x�C ��'g6cZ��c	�� @�0V��Ê�����JbZg���RN>z�U%
�H�9,ٛ,�����1�\X��Vz=ΓIpU���1cG��]j�X.�^y���m&L`��-If�zaa�f�=�xr�������q`u`���7vĕ5R���qX�v��7�l�{6X皯�3)�62'*H�IҊ9V�>� �5՝I�Vk���Kb'�)PNK ���`g�j�>�w�K�}VGK�Q�TH�E���ܝj���}�|�>� �5֤�����	��n*5I"�H	C�f:���ӳ=��S��[��:|��tӤ�b����ߕUUUP  �M��Ʒ.�T��0���5K"�[�썹P� [�v4�쵃S.��-�<�7F]*��Y�镉6����f������c\��y�1��i�6�.�9��(&�6��V�b8։���%����t��ɻ�!�j��7%.����g%����G@�d�����Ê��In��B+�f��-��ߤ�^������_<@cv�4�L�Y�l��mذ�K͛h��ף:D�r7��Y�,�f��F]�Nvq+~�y��,ᮬ��V��V�S�G�$�JH� ����H=����{����۫諭����dU%
�H��f��3�5X��uߐ��Xn�RILr��|��þ�fM�`f�����Xw�Жk�n:bJ��r�TI�`~�mՁ�.�]? {7���<�`u}�8:6ܔB@�$���LF�(������qOV�۶&�N�1�u��R���7*H�IҊ9_�;5t��͖��W}��z���gE���ӑII'7����j�`+'��X	���:����Қ�d�,�1�pb\[�0t@�HF�c��s�]X��諭H�s�j�e)5JT"��v{���k���=��}V��RN{_|�RB pHTrH�?���߰Pc��]XtG���w+]	S�J��II�`Y�,��{7��;g�Xf������$�
����K�[�J�[�H2�ج�kA�5�ҹ��4a��Lh+Q�������Tc	G'�f��Kj��5�w�@t7�`��Sꨖ�)�|����=�}_${6q`[�,��e��n�:dr� IQ)��� q��Ǳ��$z"�����#}��C�	�Md�D�m|J��l�)ZA�(���N�\Τ��z�I�S�i��ʒ8�t������?{6X纬;������΋�'�FB&:�K ���`wݓ�~ٳ� ��ﯖ��;�����ͮ���R5�;3gB۵LL�9U�:u���m�g[���4�+�M�tı�T��FB''�;r�?{&��fί��ٽ,}�8t��Jr�rJVٴ� {�Հ}�����e����i*q�R��RF�`�[,��e���n����l������"�(U�G�ê��oKu�+��ia[V��R �#J�_\4�L�}�\ḗX�h}P� V�#ZV����~��u$���rb��Jb��UX��X�z3]��o.��ٲ������nJ4�� ���&f0R�^k��,@.#^�˶����M�.����29�$�Ӌ�͜X�V� ����Wߐ���̧���ܩ#��¥UE�<iՀ}���3uՁ�d���=Kx�JB|�d"nD�X��Xn���"�uŁ�ʸ�>�;)YEJMTd"rXw�|�n��=�8�7ڦ��U%�ޖ�ݜ��J��MI,�ɥ��_Wg+���zX{���͹پ�|^u|ﳎ�;w�T� ���@���� ��D�O2~���Ś��{�߾�'�$#�?�=�G���|�;�K�d���?�ꪪ��  ��  ��\�]vòZL�f����6ѹ̺u� U��>E�|,��Gv��Z5�3.+ &͆6֠L��\1�e.�s��j/GnK��B:��z��n�AWkn	��m4�P�k��]��65ز����z*�,�$�B��YN0�V"*�G�D���MJԬn�3ڹ��e%h���m1�4l�κ��2�D�KS78M��+Z�,F�+B H:�;�>m���ke�(?�<�>n��4�riZ�7&8�]1�5���ݷVE�N���R��RF�����,��e�{3e���4�2�<zȡ)*��Q4�,��W��H5��5�Ʃ���G�n�RINTbN��I,7zX��K;���8�f��fV�d�6�$*7%�}��ٷŁ��q`��,;�w���Oy�j7*H�IҊHX�X�Y���o���6�`v��x��M�u4�l�)�,K2�l���l�Htt���]Mom:Ws-.��H�4E��UG����3uՁ�m3���UŁ��P�(����D�fl�?_[�#�U�y�"��M��U�}��O��bhD+Z}��4��R)�����͙�,!!��(0����3��H�r��1�#B�*G�(^ �_K�,��q`f���}I�vsDr!*A4Ԓ��l��x�2�>�u`b�s`}�:p�b��*�RF�a�U.�Wŀ{7�����a��Գ6��2�z��BRUN�b�����:<�_O�n���xm2��}����6�n�7*��kvl^Ĥ��FŊ�$��^uGT�Mr��;e�/�)�r;;v��y*������L��;� =���7v��$��(�*D�v��K�BGF�����RNs\��{ޙ�lo����U��U���������ޟER�iv���WP/��6������'G.R2wC'��z�ڤԥ��oA�5�'>�@�&����_�3�}�h��R�bC�!�ܲ���U�l�V ��{�tVp�7)T?�k�%1*�rD�_L��].���"%c�'�MB�%�M��<}۩�����
n��'� 30EӺ���\�D""�WQ�_�`�/�R�[�4�qcJ����
�;��ЗU�<ѹ�=Іr������2�2������>�@&��� Sl�x|���}لE���	��TԨ�"%o����o��w��(!r�>|ΚR
<!���R��sud�`�[_y��AK�CwzI�0}�`���O�;�m�I�o�AL,B�3&.��[/��h�q��]�y��g{�!����3�tMY˝Ӝ�O;҆�/J_�њl���\�j��(�w?���)��@�ڔ
d�a��sY��v�����'8����.ONB&��ؕ�>*���3�<1�ǃc�^�Ӱ���S%#K�P�C+�͇N�8�����D\Ku^��б�p]UeKT�O�okQ���cHA�D��i�Cg:p�������A���o��)��p��^�#��!:�@�b�O�����<kTN�S�VQ�&4�<����bi� ��xdM��Ǔ��μgg�ƀ����#����t� <��!���:��N!����:���|����'���@Ý!�뮇�,@4u��N�WkO p��>�1�ik��i���q�{~��m����> &�}�X�{.������=W�~�i!~�ߧ�Ifӥi/��_��~<��{�RRh����L�������K��y��?�Ԓ_����3IoO�� �I�~����f��l.lA�W:�c!�Σ�)�VP�o\-�,�M��Qw���<�r�!�B�q�ܒG���ʒK��Ē[�过��_����1$����6#�@�Q��| >���ߓ��zI���C����I/���~I#�4�����K+	��IE�b Ӄ1$�}?ERI|��y��{��:r����� {>����� ����h�g[������I����>��|�~�L��o�;�ݷL$ �o��֌H�b�ɜ!7��H5�SD�b�&)� I�ď>�K,�`��F����R!���J�d���:o�?�>���������+nL��gݶ�w>�ն�?�ʧ��ӽ�$��R��K�ٻI.�y�V�t���ԭ6�e�������94s��z��h�Kp\�9�R�m�M������8ʹ�UZ�������7�m��}��m��;�~D?!������_ ���#�r!�\ϟ ���<�I;ޑP����|�~�}������������EO���[F�����5R��N_~��I#6�V��G��U~|�}|�>�}O �����ŬZm��~��z*_}��I%����}�I,�t�%�/&o?ߒK6����H�)ȅn�I<����I/����E>��,I$�����3��T�K�<�����H��	���ΎH̝��k������ɯ�>�?@ �  r�  �&Hl����Vwl]��t���vc�L�r��G�B.�Щ�պ�nGka٦�sХ&�Cda�:�I�7Q(�fYk���\B8�%��iJ�sf�*ԺU�A-s�(5&�ma,a,`��]�#-`�]pZ)ѕ��7&��hNL��v�D�ěY�gV��p�,(��u��%�
2�5�"޲d�H9�*:h�4�	{��u��Ief��c��r*����IuԸ,��o�r:�%�x���]����As����*�5H���h������+�J�Il���3i���~�{*�_����> ���h�g[����������{����C��U������}�I,�t�����t�����t�7;��P]��W�$��_����{�z=UI�~�h�������M��C��n�
�Z���x'����Ē_~��T�\��y�=�N����� ��ﾌD{.�M[SQ��$�iҴ�_���获ߧu$���ʒK�=�Ē���m�"QF}�"^[zgL�����藑,aq�՗9��\a�\U���  VS	P�AA��19$���ߞbI�ʴ�N3_����ѻI$��R��[���Ю[3��9�> _����m����I��w&�����$�a {�߯O�m�w��g���N%���aJB��n��Ī�f�?�����c-�	ۛrs��ov�}�߳�[m�9��|����t��O����&�)3s���� {������ �o��=���$���}��$����2��Ѧs�����DZ�Mn��W�{_~�ն�c߿c{�������I��wE����������K��]n�G�����> {;��$~���bI/�w��H�֪�I~�{v�$��U#[{7c����S.�"��Q�����Y]��f��t[v�hT	���$���5Y���P��ԒO��+I$���}�I:�~�G��w�@�������~��]���F���K�=��� ����*I/��������y�w�H�M��F"=�U�$������V�Kg��M���0���)!��7��!���R��:�H��DA�S��`3�N���� kYރe��Ir��d�d5$�]ջ��x�\��!q��y9�C4��=D�X@��%�������V�K4���I,�T�
Ѷ�j1�����{$迼����/��b��o�;�ݷ���=��\�����=�r٘Ŧ����������DG�{�������C����Il�s��%��o��? 1Ɔ�5]��͑���g��f��YF5�����%�eeZ�+���<�|�h�b8���Ԓ_ߏ���$u��T�]8����?z=�ݤ���ҭ$��WO�)ET�u�%�3�����G�zO{��~���ݶ�g�.�����ٽ�P?"���~��sc�[�Ñ� �����������=�쓻������>| �w�G� ����kgb1���|��ޝ�ܻ�J��_���G�$���U����`�=&)`���5G��|t�V��)�O��w����A�������)#V�Kp��_�$�*7���;������m��s�][m�y�����D$K.&�zn]�-κ��h�gTŋ�3Cfc+R���0���:wyU�m ���f$������Y麿~I/<�q�w�t�����ߓ��������a�An)RIvϾY��a��������� }���|������ޓ�P�����#��u6\�> }ߟq����{f� ~@s��c��:����������&�U�G!W9ǀ{Ӥ�N����������V�Kr�_|������N��ҭ$�֓��"�(UN��~��G�j�m��>��~���g�.�����ٽږ���H�>�� �5e���_��1�I�`���%�0S�|��������  t�  dt����[�ǜj���J�Yua6�6�75�@�����f�.�]Y�.ֶGrե�����Ʉ�!���lo\�0b�½�(�&Wj)�P�]�Ѱ��Bׅ��L�[��4�U�KMt����`�-A�J�mK͉�� ��d�R�CL����v�fuH�:����]�&�Se��-�R��8�����-���<> ڶ��ĮZ��u6�V����Q��� ��L�j2�f�{�I�X�<.lb6�txr? ����>| �c��.�������Q�*w���c��[m�����,Ɉ�\-���?q�{�6��}�f�m�����V�{���{����S���n:�R���ZI.�{�����ߣ�{��E}}������� ���V��U6���>���wI$w�=�| ?}}����?q����|�i����$��N G�_5*ȥ�m�3�]���~�����m���~ٽ���� ���Pݬ���)[[b
��X]���ڷfV�����#�p���k���;�t��甎[����r��߯��}��l��s�� �������o_ߥ	��a��
�����}�26�@qL�~K��z�O�
���O����nL�0!� ���$ ��@��c��:�������m�s��~O{��T>ϵ���"���3���{�� ��O�{�ޝ�*~��� ��{�|�a���`�ۮ+£�����Ͻ�߮�m���7V�}��l�����:s���� }��ݬY��-��R��[��ZI.����k�3H��R�I{�5~��_�W>��nJ! A�u�n�y/�-�$n�mL���9�mv&�K4V\����'wN���)���D�-UO����ݶ�c޹ն�s=����@�sm?~}O ���ʵ��6�f|������:{�NT>�z|� ~��� /���3?x����O�A>!y�!m�*I.��嘒Z�|�K�"p� A�
}qC��Kn�P����HIĜ��]�F�Fc$ֱ�2I��Gbik�J�S�I�K�f�3O��"Ȥ"��[E�� %�g��bI�)RIg��ň�.	5#�1%��}>���$�w����o���=�t_�~~����{��6��1�H��T��y}E$����{þ��`�~V��榒��
	�P�L��D�7F�VS�����#���)l�B�5�G(�����1	(O1I����|�Y�l�7?��=��/����v�ͺ�9<��������=�tɩ��6���Ł�:������dw�$�R��JG`b���`o�M,��������_+V��?"�4N�q��!T��l?z=�ވ���}�����Y��o�l'��?i�3�Y��P	s)���hD1/�.1�6��x8�(������2��$�5��>&����c3x7f���H� ��Li��v���(���R8�$R���G��#��O�N���6�T��~���ͮ��VRj�L�ė2��TјA��ux�U3�.�1jX��$�`��sz��UL�,�ߦ�>���y������UU^a���X���G �)R�i��}����D~�G�&Oϕ~,�+}�{�'��;��{��|��]4uh��`~|��`fN�g���DDDD�O�M�k���o����uH��=� ��}�N��[����~� ����ޏDG�������]�ͥRTp�>Q�`y{5�ވ�ޏDD�����ʿd�Vz*��$�4{^É���+�C_K�8��x��L�"v7
Y�"�XV�>0(W�7�=����V��"M>�n��Qv�K�:�q�Cv�wz��hb�#�ir�a@�>x��\l۳/)��NgJo�o��\�wHF�F�d4���~�����+-�dq�
�b&��x�	LJD�%��X΋�;�e��22���p]�1�YD9>���'�/A0�^D4���_�n?:F\�t�?xbZ60�-$~�{�~�p^`�b����^�S7�A�h���/~"z�ҁ�x�)�A�@�z�$��H,/d��/��+��!@|Z�tR;� ���h�^ë�c���퐻ҋ����x����L����((��ag��c�D��yP}}|�LQ
�T�a� �:f�<���JSى��`m�{s3wT�z�����<H���j,l��y�|��>�M���B��>�'���a,H� ���+�>�����e�cb��g�8�؆��<8�Q(��w���O�bd�X*~=�^>�c������N����尢�ɖ�:�94`*L�L\s$��"Q�����'܂������Ƹ��_E��z�+���~ޛ+̎���8,�Nk>�K�O�;�p��p���3q�7�x�>���==9&d��O�����	��      ��   �   �         � [@            {c��,�Y�Β�]&�.z�j�n�3qi�L mv�%sh�,L��< �g--SCem�n��4�&��mu�Cb�l�E���u(X�[kmB���:i�f�-�mв�1�ٖ�̲��h�h�[+�	)3u-Ќ"ͫZ��[(��k2 `Y���`�XDQ��θ�Ym�-.�v��l��	�.K��2k&�n�P��Ʒj�����DL���D�id/5�䂷Lkf��8��!5��Գ)v�Ы-���ot^�U3JZ�`�TA��[+��ms�ͭ���my����;krc`���y.�LjX�*U&b�x�kc6���HX��'�y�G`F��QF��=��t�G�����/mwgI�t%�ti�䭻v���f���f��d�T��)r8P1�fіQ�.3qX�K�Z�����4Z��\�m��&�:t��zM�ƒt[�m����n�uIR�[�L�KE�p��X1+��mB�b ^�-֒хa�����`�x]6�I����ح�M,X��WLʰ�	i���0:�[u�)f��X,�u�ie�`��{-�9�P+(�b]ֆf�!,�3�F�Wh�:�����[�����u�P�ؕ�2�-5��1v�1��YY�*jb.6d�l��^f.�hITvnҶ�`,�2�U�͌���ԏT%hM0)��wmc�M̥I5�&��A؆�Ȫ^��\�.t�P�]�En�.���H�.��D�([ĭ3jۥ�ٴal��f��� ]����D�@!AF��u`:��9�%Z�Y���L0F�,��[�f��kv�]y�%r[e��5&q�����]rɵ�]�J̔�$����9tNܶy�-���<�|�kz�#k����Վ�-,h�3+e��1����ű��5�)�.�ƌFiJ7b�4Z]������:4�)��f֚f�M0�#Jme��n{h9�č�s��5M6r3�M$:Cb�WK����@>L�Χ�"�1�t��|�4�So`ë�'�u<�c�����tGi�2�et!�"x��'�t|��D8!��@��|�|��׆��R1#7�BlC�-2�*� �A�&�<dB`�õpm^	vNd.C*�<p�9�����D�t'�P��և�p|hzaL��1ӽ�|o@�@�h���]'P���  �� kn  &�ˣ]v�s�Ճ��W��\[���SA��]�т�2l�|���[�v�l���6f���[)2�GGH�gd2X��h�*هJ�K.���c�Zf��T��p���c1wYU�h,�2��P�ka-B�ѷ]��L���Q��2�f6�F橵!q�t�(�A���m*6h��ڴxa���q�]	�t�!'B([E%*���()�M�;��M�˦Anx
4��]L�cv��.��a�Zm��غ�VW�>t�<7�i�ťcD�T�������X��w���,�v�]�'Q��u��KwS����G�dn{��M�}����D~�$��Cﾌ�Y���uə������ō͟����DDɯ��?w*�XC������a��'��$�wM���ym��~��qa�腻O�����
��P�*�U4��n�ޏ{�����}����Vy����dԗ6܁�B��J�et�fe�V)��5�6�e�k���c�Y����>����$T�J���O��O����Z�7%��"#��ђ�ߪ�p���%! %	�"&Hi'�����a��ؽL�)�3���MP�D,s�1�^!�_�R٪P�/��  ��րm >�,K�ݺMı,K����&�X�%������n'�Vb&���߿{�E�m����O��zX�'����I��%�b^wﳤ�K��q?}>���Kı=����>^��^��}����,ZV-�����bX�b^wﳤ�Kı>����Mı,K�Ͼ�Mı,��]z~�羞t�z�z��=��7;;::\�g9�t��bX�'ޞ�f�q,K�^�>��7ı,Ow?}t��bX�%�~�:Mı,K�����m��4څ��e��6U�J��1g#L��'7lI�S�h�N���`Sy:t���eZ�4�s�L�q,K��sﮓq,K��s��I��%�b^wﳠ�$9,K��_�4��bX�'O���ɜf0�.L�c�Mı,K���]&��
"b%�{�߳��Kı?}���I��%�bw���I���*"b%����!h��.O:|�н����Mı,K�z��I��5�$����?Z��7!LD�I�gC0x��a�1�%�7��SAN�X7`�O#���l��?��ysPN�Ų93����	#�]��b""-��b�mc���&"k���I��%�bs����7��zw߿�MhƊ��O��z�\D����&�X�%��g��I��%�bw����K��~B��b'}��SQ	�鏱�4�I)�l��M	 �'9�e5�~��{���O�,K��~ޓq,K��޿l�n%�bX��C��}'���1�Ɍjn�F�j)3"JQt.nk�C:0R�%�ep�֢�W?:I�s�X���*i9ı,K�~��&�X�%�������bX�'���f�U�Kı;���y���^��^��￶�bҭL��s��Kı;߾ޓp��1������&�X�%��g���Kı/{���n'� ���b_�{M�ȓj2��:|�н�߿�vi7ı,N�?}t��c�H�b&"_{���n%�bX�����n%�b��o�߆U��Lg-ə�O��z�1����I��%�b_{���n%�bX���oI��%��Χe�\;����ܧNN���g�������2f$_�[R/�t�S�91��s�u��-d�3�! 4��Ç�."X �P(��J��`�JŢ�BD����|�н���{�szð�짝>D�,K���:Mı,K��\{߿gIȖ%�b~��_��q,K������O��z�z{;�~����Z�N��D�5�l���͸�w ܍�)fl)r���6�����;�n���AZ0cl����"X�%��~Γq,K�����i7ı,N�?}t��"b%�b_{���>^��^���߿{��E5�5vs��Kı>﮾�M�� @D�K����I��%�b_{���n%�bX�����7�,S1��韱�T�(W�D����^��^�~��x��bX�%�}�t��c�`"b%��~Γq,K��﮿M&�X�%������,X���*y���^���C1�}�:Mı,K�߿gI��%�b}�]}4��bX��"{����7�н��znX��S�'�>^�%�b^�ﳤ�Kİ�, ���ND�,K����I��%�bw���I��%�be?c��`�w��k�0���0	$����4B��0Z�z���js��~����Y�V�$��V,$��˃$!+�9!�~}|�� h  ۖ� ��%U�ɸ�KYk۰�v�1�
��4�fh�M0�Z;$�i��;3V�vG��6�7d�5.,tv�Z2ĵ�C=1��٣	�5o&���`oV�����!J�ײ���t���`ь�vHTĕb@@��ec����j�YSZ:�l]6�P�5�
i]fZŘ�9\\L6]6�uٍ,�Ģ��8��&��0�$�Ӻ�E/�� *4Q�Jt�;���BL��|@ZSL�k��I6��\�����έ'd�h�ɚ�R���������7;;:3�����z�z9���f�q,K��s��I��%�bw���A�@�����%�}�߳��az�zM��F":�1��&g�>D�,K���]&୉bX��}��n%�bX�����7ı,O����t�zIн��7���1��5�5�t��bX�'{�}t��bX�%�~�:Mı�+q?{��I��%�b{����7ı,N=��-��e�rd�9�n�q,K?$T1����n%�bX�����I��%�bw����K��$U�O{_~�Mı,K�߽�M���5r����^��^����l�n%�bX~P����߮��,K������Kı/{���n%�oB���w����]�c��r+[@���[-u5��F�o��O<l"g�Pk�M6nM���I�3ʻ�R,�q4L�t��н����.�q,K��sﮓq,KĽ��gA�H
���%���_�4��b[н>����,X���<���/K��sﮓp��;����$ąFZ!~�$&@�3HI&,�{�F�gX[&)�	��0_ �C�A"��*���0�+j�B|�"b%�w��:Mı,K���f�q,K��s��I�����I5�B�>���b݆%�Cf�7ı,K�~��&�X�%��}~٤�KȰ1=���t��bX�'���]&�X�%�z}�Üc7��g%��s�&�X�~(."~���&�X�%��g���Kı;���i7İ?
@W1�~��&�X�0�?���sf��[�3Ο/B�"X��~��7ı,?$}�}�ND�,K�߿gI��%�b}�_�i>^��^���'���}v�PFk�smbcT�;+M�Ģh4�*Y����4�e�D���$�g���1��)6k����/B�b{��4��bX�%�~�:Mı,K����A�*<���%��g��|�н�������4��s��q,KĽ��gI�~��"b%���_�4��bX�'��߮�q,K��;ﱤ�D,K���}�css%əs3�g:Mı,K����I��%�bw����K)CRؐ��0�`0Al����v&L�Q��1a�X��yٻB�'R,iA��*V���P��,Lc]�4��bX�%�~�:Mı,K�f}��3L�3���q�I��%���."{����7ı,Oc�~Ɠq,KĽ��gI��%��b}�_�i7ı,N���ƅX����UO:|�н�����n%�bX~P�.=�߳��Kı?{��f�q,K��s��I��t/B��I��@���L鳆k"Q��juV�%��Rf�q�56�.Ο;�uw��.5b\ƙ�t�^��^��{߿gI��%�b}�_�i7ı,N�?}t��"b%�b{��4��gB�/C����ܹ�ї<�����^,K����I�~��"b%��g���Kı=�}�Mı,K��}�'���:Y;��5�^����Qf��s�sq�I��%�b{����7ı,N��Mı��@W1�߿gI��%�b~����&�X�%��O�3j�W7\�SΟ/B�/�%�;���>��4��bX�%��~Γq,K����l�n%�`cQ��3��<{�~���4�ɽ�u��s�����!Bl\���S���"�a���,��4ಀ���e�[7ȱ�Y�c�z��#��H�j� T�BE��"k����z�z�������`c9�t�Kı/{���n%�bX~ ��_�4��bX�'��߮�q,K��;ﱤ�Kı?>����6ܙ��4��U��L���lI+v��i�tF�-�-�cz�2���+�N���>�F�l�|�Ȗ%�b~����&�X�%���ﮓq,K��;ﱠD7ı,K�������^��^����w�R-�Bh���i7ı,N�?}t���B*����b{��4��bX�%��~Γq,K�����i7�	Q�LD��ٿ~�jU�ˮn%T��нЉ�{���n%�bX�����7��U1����i7ı,O{?�]'�нн��.2T��3�鸖%��H��"c���:Mı,K����i7ı,N�?}t��bX��������n%�bX�ǿ~�q����1�7Γq,K����l�n%�bX~��~�ND�,K��߱��Kı/{���n%�bX�'��7�*kq>�Sw�ɸLa�ޡ5���2H��u���~}UUUTm� �I� L�̸`0*ִ���t9�]Gk�^nڂRĂ݆kZQ+�i[J�c�r\�7�%�Ű��쵣b�`��#���WG#a?��T��8�4"���"����53�:�b�k�kٽ���f��iZ#��@n��;X�`��l�mB:�J��sCZ�[�\&5�%t(B�m��`�+bS��h�V�-7�'���q!ćK,�K�0�o��,�[bd���;f\fف 0�Ω�0�2��L�Yk3R�����wv�y�Z��M�����O��z�z}����I��%�bw���n%�bX�����?���1ı?{��f�q-�^���7��c*�c4�*�t�z,K��Ɠp��T�LD�/���t��bX�'�}l�n%�bX��~��7�0�LD�:����c��%ɒ�\gƓq,Kľ����n%�bX�w��Mı�,U�LD�����n%�bX�Ǿ��&�X�%����t�e���Ο/B�/�$�$���￱�I��%�b{����7ı,Nc��Mı,�Dǽ��t��b[н>Ϸ��ʑ�j�l�:|�ŉbw����Kİ��;����'"X�%�}�߳��Kı>��<���/B�/Og����mm�RZ�kt�$m��"kCD��m��	���ԩ.�`�|�c��L�\�J��O��^��b{��4��bX�'q߾Ɠq,K����l�~F*���%��g����^��^��߽�ŋ��.cL�:n%�bX��~�M�Ɲ4j�\w.��)L�`,IbL�3Q�1<	���������lc�N��#�+������OE����B0㦴 VҐ
@%cZҌO�%���&5۽�Mı,K�g���Kı;���i7�D�K���Cs���ncL�:|�н�߿�vi7ı,N�?}t��c�X��&"{��4��bX�'��߱��K���~��Q�i�Q3<���/B~ ��"{����7ı,Oc�~Ɠq,K��;���n%�`~
b'����>^��^���7��c*�c7c8�s���Kı;���i7ı,?,Q=�~��'"X�%���_�4��bX�'{���Mı,K���߳mɛ��u��Π�[bx�^6�f]��:%��I4���:Y-��Y���$�+�˝F01��q,K��;���n%�bX�w��Mı,K���]�b�Ș�bX�Ǿ��&�X�%���n��s���-�nq�i7ı,O����&��Fb&"X��~�t��bX�'��cI��%�bs��i7��LD�<z�=�R1�Bl��g�>^��^�������n%�bX��}�4��c �>�(L�_@#��~���~�}~g��
�!���f��4�_"L����ۖ���~?�/.�$_Şk�;3s����G��G��LC�7�����2a	��3Ai��y���A����@F+�7\v�W����?Y)��64�Ɍa�V�I�L��o��,Y��8.% ����_L�A�y� ��	X9k�G�}�ND?�s���j�����b��0B ߠ�`��wÁ�~���[��}���� ���  �{X��`�ܓP���^�B�A��C�}���	U��/!{H�'��͓Y��8�O~"l _���z2�4��Y:�����������P�}>��IVx��x#g̀�X7d��!�G�m��)�(�|8ɦ�ZT���4Ip!}�Q �R	L�/��h�~E`ܛ�QpjAHAAnx��oH̘��Q��ݞ^Z
-y>A5�ؘ+���?qߋ����b�
����F!0[		�H=�0fg/�	�?�i��?U�}���]`�ݸ�Pؖ�Q:>��*��$�+�h�.�R1�
[�c,�>0�KS�;c�~50mjx�)'&1��c��=��|���L�P�	�� _K���1�G�1������#j?��b�Β��}�~��|�
ba/�-s��� F"�kȳ���~+ ��IoJ�i����I{�э4� �w0}�����A���M�����$ђì,6�X�KP�f~��F��{��炉C�YS�D�6J�pf�>��0�����S4�M�a1���:�9bm:M��N�]��!�8�SGxGÀ�C�wɀ0�@��T�S�u2�:0�ӱ:@0��<��� y��J������M�t���{��+ Ǌ��9S��H@����<@��s�_D��+M�N{di��L=��4�v��z�y�0'R"�\O<�x���������Cè;U��B!�i6ʞNV���<�IÏ��P\z>A�y�Сh�KZ�hT+ �@�ƥ_��&"w�q��Kı9��4��bX�'L{�`Źɜ䘘��&q���K���Og�~Ɠq,K��=��4��bX�'���f�q,K,N�>��7ı,K�{�9$1��2S��a�G�|5����aKıS����I��%�bw���I��%�bw���n%�bX����ߤ�7m��H��W��,����K�$n�MDLT):�����i����D��'$��7;;:6�&e�q��Kı?{��f�q,K��sﮓq,K��;ﱠ��D�K��=��4��bX�'O~�����!�ڑ���a�G�|;�ߕ��?�LD�=�}�Mı,K�����n%�bX�w��M��� �LF����}��Ɍ݇*�t�z�x�=�}�Mı,K���cI��?������]~�Mı,K����I��/B�/O�}�X~\�1�9�t�K���Og߿cI��%�b~��_��q,K��s��I��%�������o� ���mu���/RO��`�F��3O������}�N��$�[0f���L1Z�D,F��
1����\D��{�&�B�/B������!2��x��y���ı,O�믦�q,K��{_�]'"X�%��{���n%�bX��~�Mı,K�'�}[ym�d3����E���8�73t�04��. �eH�օh�jh��|�,�Wʑ�n�g|���ŉb{����7ı,N��Mı,K���cA�@�Ș�bX������O��z�z}���t��Yu�Ī�&�X�%��w�cI�~�"b%��{��i7ı,O�����n%�bX��~��7�,K�����L�\�%�L˜�I��%�bw��i7ı,O�믦�q, �D�O{?�]&�X�%��{���n%�bX��~��9�vtmZ�;Ο/B�/�%�ק�=�Mı,K����I��%�bw���n%�`~B"{>��Mı,K�>��uGY���[�O��z����]&�X�%�������r%�bX�ǿ~Ɠq,K�����i7ı,J�,�tC�ퟷ!����Z����#z�$ss�g]ͻ�u,�0γ��X{4����y�UUU�  ۤ�  �e�,������k�z%�v��	ˉ�z�I�i�J�R%�%rM
���;°pJJj�HT1D��壳3,ѽ^̶ٴ+�ݢ�z-�-��lPz�[��R�jj]�6o��T�nCM`h-�*:�M���f)tX�BT���X�f4��`�]fc v�
j��X�^�H�E�m��wJX�E���v�L�CuL`�������S�R���U) �h� Q�T�]kx��6��M�B-��Y����ڷ��9:$�W�I
k���(*?�Nc��eVL,�r��r%�bX������n%�bX��~�Mı,K�����)�1ı=���t��bX�'_}��s���&Ifn3��I��%�bw��i7ȱq,O�����n%�bX��~�Mı,K��Ɠq?!�LD�:���*�g��:|�н�߿�=�q��%�bw����K��D�Oc�~Ɠq,K��=��4��bX�'���|�1�X�3��t�z�gB����]&�X�%��w�cI��%�bs��i7İ?)�O�����n%�н>����\,�.�����O��ı;���i7ı,���cI��%�b}�]}4��bX�'{�}t��/B�/Od��}���[t�432R���	�t��+]�3�++��B�jF$��5��]�?$���E��y��z�z��߿cI��%�bs�k�t��bX�'{�}t�B+Ș�bX�Ǿ��&�н���}�7;
��զw�>^,K��~���7
�yK/�'=�u���Xoi0�7 1���o�Iq��f���3��C��"�˨�VGHt4��1"T�RR�bV5'�q,L�;�t��bX�'1�~Ɠq,K��;���n'�b����'O~��1]f�c:�WΟ/B�/B������Kı9���i7��0D�LD�=��4��bX�'}��ޓq,Kޟ�_ߣ*�af×'�>^��[!�B����}�)�$�v���hI�7�ze5�> ��{����n%�^����~��s3�e9�t�z��bs��i7ı,?E�~��r%�bX��~�t��bX�'1�}�&�B�/B��O�~ݶ[T�l�W����ɦX��E�-&���[u�l�ቹ�k�e�����N�y�!2��aW9�t��н��?�zMı,K�Ͼ�Mı,K��ƃ��D�1ı;�~��&��z�����Čy�*;gWΟ/B%�bw���I�~@ ���bw��4��bX�'q�߱��Kı9߾��n'�8���'�}��91�����st��bX�'q�cI��%�bw��i7��;�c�ҁ��
�b�ze0��4<-Z�"�-"�Ƕ�L��&mː+H�`P�V�$`T+H%B՞P�K�ֻn�q,K������n%�н�߿���s*Ƌ����"Y���'��߱��Kı;���n�q,K��s��I��%��B������:|�н��>��nv�o3jˌ�I��%�bs�k�t��bX��H���߮��,K��=��i7ı,N�}�&�X�%�����v��l�L[Y��e(�ۈ�
��s�t�݅���F��-b	v�M�o<[�u�m�����'"X�%��g���Kı9���i7ı,N�}�� �"b%�bwߵ��&�X�%����ْc9IJ9$W��>�#᯾���@q1��=��4��bX�'}�_��n%�bX��~��7�1,O?}����3�e9�t�z�z����w�>D�,K��_[��K�E1=���t��bX�'q�cI��%�bq�����YL®s����/B��%��N���[��Kı=���t��bX�'1�}�&�X�}�Kc�c�g����/��<�w�j]0$,J��@�IA�
%*�<�'3��Ɠq,K������2e� ��:|�н�������н��bw>��4��bX�'��߱��Kı9ߵ��Mı,K����O���-�Ln�\j6/5%��Z�As�+��K1�c:rcV���o<��fњ��\�7IȖ%�bw��4��bX�'q߾Ɠq,K��~���?,D�K^�~��y���^��^���ޛ������s�i7ı,N�}�&�����bwߵ��&�X�%��g���Kı9���i7��D�K���e��2�t�z�z���|�n�q,K��s��I��bX��}�4��bX�'q߾Ɠq,K������0��k�ήP��н��bb'��߮�q,K��=��i7ı,K���t��bX����~��t��^��^��{}������U<����,K��Ɠq,K��,{߿gIȖ%�bwߵ��&�X�%���ﮓq,K��!�L�y�f�S1b�搌�5���Mc\��3�zLju�{����4���z����Ϟo/k{�u������� m  �� m��件�5���h�Y�].��+|�b�i��6�qH��mj�@�.��5�p�)-�%�ݢ�h�qtNl����;�k�\fƈL�A�&eJ�\]��5�-0�CK5�l��T4�6)��虭#���e�6�$u��c�K��KM��GjbU�S	s1���κѐ����F������]��׵�uD�Y´DBe�ڶq�3���ҩ
�ZJ�aV����x��Q��.R	1u5�%��J�A��m��	���r�`�t�{�>y	�Q��3%̹�q��Kı/}���&�X�%������n%�bX��~��?��9,K��߱��Kı:��픵U�XT\�t�z�z��������?1LD�K����I��%�bw��4��bX�%�~�:M�� �q^���~��#u���P��н,K����I��%�bs���n%��"8������:Mı,K�����>^��^���7￴�,4f���S�7İ��Ɠq,Kļ��gI��%�bs�k�t��bX���Ͽ|���O��z�z߿znV��6��q�i7ı,K���t��bX��H�����IȖ%�b{����n%�bX��}�4��bX�'��ڿ���h��� 핰��)W.s�2��[�*]0�R�j����o����m��ֹ|�,K��k��Mı,K�Ͼ�Mı,K��ƃ��1ı/~���O��z�zO������6��8�m�n%�bX��}��n$��0F8�����;����?��9f�)l�X�B�#
"��*�
�&"b%��w_cI��%�b_�{��7ı,Nw�}n�q?$zkн?��}������U<����,K��߱��Kı/;���n%��"b&"wߵ��&�X�%��g��Ο/B�/B���|���ff��G;I��%�����~Γq,K��k��Mı,K�Ͼ�Mı,ʤ\D�}��i7����'_����3��R��_:|�н���zt�z,K�sﮓq,K��;ﱤ�Kı/;���n%�bX���~��~�v�h�um)n�ΖU���Z$�a[�����7Yu�.�[3����y�b6�ߤ�Kı=����7ı,Nc��Mı,K�}�䜉��%��~����нн>���t�,]sq&s���Kı9���i7��1,K�~��&�X�%��~��t��bX�'{�}t�������%��~�33��f�Ս3����/B�/C�ﾾt�z,K��_[��K��W�)I�2!�5I@�!rc�bF��r�3��h0�JF�R�!JO�D�Oc��cI��%�bs��4ϗ�z�z����n\e���\�t�K��9ߵ��Mı,K��Ɠq,K��;ﱤ�K���LD���}|���/B�/O���7��u��Y�g6�7ı,N��Mı,K���߱��Kı/}���7ı,Nw�}n�q,K��?���~�1��"�eu�.���8G"m%A�)k�M���lK�`fN�i�_�_��&�����|�Ȗ%�bw��4��bX�%�}�t��bX�';���I��%�bs���O��z�zw߾B~V�n��G;��Kı/;ﳤ�? �1,N���[��Kı;�}�Mı,K��Ɠq?$�LD�:���ɜ�9%�l3q��:Mı,K�����7ı,Nc��Mı�C1��߱��Kı/}���7ı,N���3s&\�2�l�y���^��t��ק�����7ı,N��~Ɠq,Kļ�Γq,Kzt@���d�o�����Ѓ��]��探r��G���LHew!��!�t�Ή�]o5}�D4iFQ�HB�a,�X�o:�t�z�z�ٿ~=��*�L�D\i7ı,Nc��Mı,K�@�}���9ı,N���[��Kı9���i7ı,O�~�W���m��8�3��%�����B6�v�E`T	F��3n�m����i��vt�]熍Z�fm�i��O��D�,K�}�:Mı,K��_[��Kı9���hwı,Nc��M�/B�/C�~���v�h�֪����ı,Nw�}n�qlK��;ﱤ�Kı9���i7ı,K����7'�z��~�~�����(y�q,K��;ﱤ�Kı9���i7��1��~Γq,K��k�y���^��^�����mٽ�Y��s�&�X�~X�������n%�bX�Ǿ��&�X�%������n%�`~H�����i7ı,O?}���3s13%̹�q��Kı;���i7ı,?
{���n��,K��=��4��bX�'1�}�&�X�%�����<�T."1�&�0|����c��\3�^���^ѧ鱳ͧ��<�?�����5�Q�Ҿ �7��Jѡ��0s͖�Ӣ�{u_S�{���JaY��نrߵ�LL�!�0�nO�~X��8_~A~�c���r!���������!�Ea�/��`�@i��"e�qy�{X�7e��\��N�gyԮ4!C:���n��Iw��=N�����OľۈcdߎOe7y}NC:��=}�{�Ј^b�#FVS0�5du���̹��߳'������>��8&-��BhP�&��"�P<�i��-0��#�I�%�t�I{��<B?BL�!�D$ ���_L>d�RԺ{K�	�+� ���=����}��m���Ԅ�I��#�~���!oo�}^nЉ�}_�<`���(?&	����e�GGS~�����&фa�=IA!"�"�O�[��M�@8�
���ು�Q �vx�����������^'A��>S
��G��C.c��\��ƹ� ��b9�$� �7u��-��phZ)�lA����?A;ޫq��r����@���9�>�Q4��������3�-+��$ly*�$9 0%�*YG�@��B�0�%dƹ�\��&��=sk�(��n�y�7xj����J̚�L�MR�B$ܥ��|	�nx�1��܁f��M�g�}짤���<�������P           �            � $             ��8��XI1,�Z���D˯g�u�kiHfn�E�;cBee�X��SR��5�Q��k�4��Fcml�k7����+c��)s���#*֤�ѥ�5ͷF=�(�X��-� 5u���[Z�[	�nkD��5�65ڏU�e�`��1�͑-m4z���Z�)m@��Y�K[�6���Պ6��̀K�,.a���.���iJ�{RЏNXj�F��k�&�^N�Β�k,ѷ7*i�\[Đ�7SGv�Ǝ�T�YS�]�5�p�bi����K��&�1�L\�B�P�-V7b����MZ��V�!k3�#r6�&�3G����I�v��V�Z�.��I�&��q�3M,�+��BZ�n/1�˷-4`R�4��%��⹸- �+�.¤l�툖;�����]jB���̗XRƬ+fG]*;��JWgZ�]X�,� GGm1rMufe��r]&%k*M.a��-�Yf�f6YZA�.��*Ҡ�ItN�0.i�i�m��f�M�YLdn���R�H��i��Kk��˭%�TI����-c-+q�]���`��.���ko&�9�9�l��Í �Z��,ev��E�\LL����m]CP-�6-�MfM\��u�R��6ݞ4@��5�Eژs5+l���M
l�K��0X+���	����L�<=J��j���[3MR�b��M�1]���6�����[ pa	�Y�v�Nc��XJ��%f�[1b��9j�5%��@ڲ��M�&&Xe��r�J���e	��n�;f�`�[	t@u5�b�-ݵ�WZ�Q���4�,l\Q�֢&`Y�t�J343��'���̗KӷLdoDڝv�ku�uS`1ff����4��2�vv�#�#cq0��.��g]�ft�7��.��^�$����pK��2�X�
���9�-��б�f�rZ瓦�tաZD.�m�V�q���庤�&��K�I���	�Mol�wBܑ�0�TK��ӣ38�\�8���3�������G�=�����f��.G��"i@��vN�^��8>z;z��L������/��iD��0^ux���e2�����ߗ�#�7D��_'��{ʝo�á� ��<�
�p� ��:��8�M�C 2 ��`M�]�2>�z;xS���'>����zՀx���r!���M�z��<���N>�uZuO<���G����I�ψ������s�� m� �-  	g2F�v�K�oi3�y���8��$�;S�Rv"Qы��
��k0+5EL����se�Ւ�a���#sq3���Z�˻��ke�����0k�(�-���ٖ6���pV��2\b\	.��Z�Y�D��'gS��<ƴ��ˮۥ[M�h�n�;/i��v��i�M����6�JK��C�����:
��8�P!���wS����^�Id��ݭ�M��L�9���i��vm&t�Ae�8�4��������	Ụ^\�����/B�/O��u��Mı,K���cI��%�bs���~Br&"X�'��cI��%�oO���=���%���*t�z�x�9���4���8���'q�cI��%�b{��4��bX�';���I��d��Mz��߿�U�f&m�i7ı,N��~Ɠq,K��;ﱤ�K�$1;���n�q,KΟ���:|�н��}��͋Wf�əq�i7ĳ���Og�~Ɠq,K��k��Mı,K���cI��%��b's�cI��%�b_�?c�q��f̒�8��4��bX�';���I��%�a��>��ND�,K��߱��Kı;���i7ı,O�g߭��e��l��K�%͛0Ə ��AԺ�U��f"�G�F��u��癑����v&1�۴�Kı;�~��&�X�%��w�cI��%�bw���~E����%��~��t��bX�'����2Lc1���nH�|�G�_}��"�p~��7�-��f/��r�i�r�r4���	��fs{�x� XK��IaHP�[����C�"X�'�~�q��Kı?}�}n�q,K��;���n'�1S,O?}���&X����:|�н������O��ı9ߵ��Mı��LD�=��4��bX�'q�cI��%�bq���l��Q�.Wy���^��t�Mz}���t��bX�'q�߱��Kı9���i7ı,N��Mı,K����.��K3��T<���/B�/O�;���n%�bX��}�4��bX�'q�}�&�X�%������n%�bX��w�����յ�MMs���[�9�2�V��$�m[��7sm��Yuv 
��6�eY��79�ӑ,K��=��i7ı,N��Mı,K���٠���1ı;�~��&�X�%�{�߮333s�B\������>�s�;�,q,N���٣vN�~��I9{ﱯ���egrl�܍@�'q�Μ���罍Mߎ���~\=�D�w�qIq�!�Y��`�$�����4i0��RLI � ��$!e����Ԍ)J�BФ�o��jI�����^��1��܃r%a��R���1k�1f���Dzo_%`ls�Su
L��Q�#�?/f����{�?���X���:#˹���UL�	�f���YZ�]��kp�3�YjX�u�h�����u�v�\��b��h�|��ߺl��J�ō�G�A�_M��o��H�
�rX��R���1gs�<�y��n�꯫䌭���)A*r�jj�+V����ΏG����VoNJ��-ŠI(���E#�ꯩzu��ouXc����t��zE�(�m3�$LB��0d�r<߰_sYC�k����O��RF�`���R�
 �<|04�F��-!w�w�jI7߽q���#�P�'�~��:���u�_�ś������������6�ĠJ�36Ķ$ʺ�%���4�{**� 0B@4M�Gb2����r5P�$��Μ������f��{��7���ꞥ*�H�BrD܉X^�v���`��,o��'?����1��j7$t��ù}�՝�%��h�5k�3۵	�ʒ�dv�%����%`y{5�u}K�7���z�*$�u>���Xcv��ލ�}?�_M�}�Հ���Q���"�˷VP��T|I�bE$�1�X%���D�����h�������l  m�l  m� �Q6�YV:L��xsq�lK4�2ݥ�s��(��+�m R�]+6κi�Hʷm�i�a%�rTt�4�]����%�ɝD��k���hk�"\�܄ �`�s�nmщ�h��-�m,�Z]�ĭ��d,ƗHM�5k]�eauF�%BXd����Ն�M �e�V�X�R̽m�fi��d�qS���a�Y��Y�M���,'^��K	ץ��K�O ��*�%\�leY�匦�%d��T&��� ��Zf;\��Uf �(%NS�8�,/w;��k��ݝ_W���E����J�H��ٮ�͆N�`{;���]�A��N�G*(
T��=�����M+3��L��hZ�l#4^�2��	3@�����-}6�5͇G�/gt�=]��MEڤ�q7"V�k��������>�M+����~@[6��M��DQX�թ��;.�iԛ<Kj��!&ɴ�-�ky8vV~�� �n���K����l���r���AG�{۲��Ug3W.�0���[�.0c5��%��rK���î(���I4�	��}��֨bYb�.Jl��4�"@��
�*Z5+T�FS�ĬY�6�5��DD$g�넠��8�K�Ӓ�<����ٮ�=��`z�&�PR��rD�:=�w�lZ�l1��>�M+!f7�P6�E#�?/f���������%`~^�v}ݼ��܀���Û�kt�E4����*K�XV�:�6)����ݷ ĥȊ�%r\�RO�����tҰ>X��,�6����)�t@ND�?{f�}_U}IY��,�v��]��I��sMEڤ�q7"T���~t��{�O+8�B\A&RŰ$�gد�d$�tW@�m�7S��BVE�6e�y/t�GA�8&�,`�b�,H�~X�����j��k݀6D��n��ýY:�lZ�l�ӕaޅ�����n�U��r�dv���`w�9��|-}6�5́��ͦ��ą"t���k��M����%JCkH.t���e�s5�ܮ�ۮ�OA��nd�a�@o��rX,�6�5��G�1k�6Φ�)N	T��H�,�ٮ��H���`b��`|�ܗ�		�� ����D�<�y���]��R^��e����?fjp�Q8GJ�q�r���`g>�,�k����>�ϥG�zv���7���Ƴ0�t�~��l����!�,6b[3\�߱
�H >�� �UW�B������eG$�R���jl�������u��-}6�5���yZK�JB��Ң1�!@8��k4ҺGh�7.��:h&��]u�ʱ���\��Q�ڤ�q&�?��������ٯ������h�2��@�q�J'����=脌Z�l��E���s}��RF}�)WG*'Pq�Y����E�	b��`b��`g�]�QJ��Q����w�����o;��k���y��2�gSU��AƤq��5́�:�~�����$|@dx5�`�ղdkh#�g~��O�6�l�w�y�򪪪�m  6��  kQ�̷a�:Xe<�ޭd�t-�jfXV#�-mKsf�ٜ����c�k���fVgn%&n��crgܘ�cM4X�W��{=$ܮdK��&�MKm���d� �����bᬮh�ҹT���Yn���WX��@5�f��5%6ݮB1l̩���lR�F�]n���h���CSK-9��U����q&qs��E��HF�U��*��� ���ɼ��1�Ɍn�].2kflk
B�6�d��-����k���Hm��Gis�eYn��*"�߇����Y�l��E�����>�jh�J�bG:�q�^�w�W�RG���`ygs�?/f� �{u6TrH�IƤv�ݢ��csg{�	b��`j��`<��Zj(��$㉷a�U����`b��`b�saވ�����OuL�ѵ�NH��ٮ��o?�{;����`wۛ|���!j}�9$i�l�WXͥՌu+�2Fŝ5^��Ȓs2��uf��J�jT��@PQ��Y���ݴX,nz">A�_M��o��U4LT�ET�T�cv�=~$���O���$�94j!dCS$�!�R�}j��>�@̆e]{� 1 Eb�"�	R Pl���6�[�77�	�D��Q4%R4㈰1gs�?/f�:��Kw;��h�=K1�(�����"�Ga�舅����ս�`}��,:#�g{��=���D�u#�I������:��f�|��ս�`|�\����\��I-M�8U�Zfi]h�;]�n�v����a�	u0�%�n��w^#i��3[������X���>Y�lX��#i9N5ڥr6�,/n��H���`b��`~����=\���UPIR�����76g�����<���FB(/<
G>�w㠏�}�͉F��~OޫtȠY�Q]���a�eEN��(�Q�F|��޷�9܇���H~|����H1��)=�ʟk~y�#Z�� �K�L�Ϝ'�ĊƬ�{̐{�k���	�L	���ax<}�A4M&�GS�!ԘAS��߭��;����H�A��=N�"A$p�|c�S��a�.<Ѽ{�}����P��FIB���6��&JA}���)��<� R�֘LQ�Gl���'�w�u��5p�.��{�8����eEI���QcJ._@ |DO��>1����Z���d� n�����N��mlIJR�((�#���⒋�;<��.��:�')%+�ԓ�TJ^������0�<���L��`}Ɋč�.9�����ɾ�Z�@A$y|~�?u��U�n�cؔ>> �Ix��I1q�i�'d���ߠ�ƍ��p����V���0�6~B2�@
Ў�L��&v��"��8q�#5o��f�q͓�dٝ��U`Rd�)`c�g.�N��c�:����X2!��T<�D<�h=4�A8�n�/�@6l�ּ=v d�'N���|��ɾ�=�������ؒ*M����8	�ED6pN+�<�"yt��&��!��j3�v:�m�8{I �����<de6��"���T2:g���=�,��
��u;IA27�8�τk��xD�� �p.P�:���go|�
��U�AH�)Q��Dl�s�Y�&�s]��"�J� ((����c��3{�,nl;�'_M��o������T�8��ݴX�WՏ���<�y����������D���4�0���De��k��!{uǞ,��[c����j�-Qҹ���Ћs���o�������Ս��f�Z,���U@6�H�?/f���#Vw;��h�<�5�U$���"Q�GR��'&�k{����Yޏ%��M��_M�e{Ml��Lq�)q�w�UK����}6�5̓���>��>���wX����h�3�#�وh���E��I�y�(� $R E��"�V
Z�no�{�o��g��RhmTn)q����<��՝�����E���V�֗6ے
�e�cH�MR9уD��vBMW��y-�t�Ļ<EíUr��@t�j�M�������s`}��;���5s�7�ZGT����%
8�^�w��${;�.�v�����H���$n��q�L��E���;�K����#v����8%NS�8�,:�X�y�Y�6�nl;�7��X	�� ��
r��q���]��U�;��=�֋	����l��d��s�	�H8x%q�����cF%6IL/)� �{F�v ��>	��>�I#m�-�� ܴ  -��ZM���Z���Y�/Rk6�7;��*9�V3�����h�X�-����1t�uu�̶�(��ݎ˰j���mp���K�st*�%�]\ұ!���ن��9�"��i�+��ˬj��%Z�IH�ʙ��ҙ�F�3\��(J�`l�&��Kf0�V�5�[4Z2��7��b�&�yF�g`�V��Bc&iqr����F0BP��:u���지6��gvͬ�n��F�Θ�P��`�ԍ�a�X�QY\�¶G�JR��v�n���m�澯� ���`Y�6Tr*n)T���cv��6�5́��ﾪH�!�ĚPN����o;��Έ�I��7��`}[�N�6�!D܎þ��^y��Y���ݴXw�o;>ש�)F�
���Ս́ޏFow��\�l�k�-��q����ݭ������0��ks��i��л9l&R�$#r��E�A���YI�੸#�?�{;�����k� ՝���ݝMTR��)Ɯq$��}�c�ǚᵣ�W�>�8� q37�=.}��Γ6R!w~8V,�
��A{�P���lOzl��E��	u�(�>l)�"�G`yf�<�����wZ,Y���f�G$�JR(SSa��-��9��`b��ý����2�xl�$T�%E"R;��,��ů��ṓވ�9�'�m��IѶΚ�铙m�<��0��2�m�aiSY�ʷ8�3�l\!���Dff��[�6�5́���G�3�\���u@t�j���;��k���$j��3{�,no�=	�-.Q�R�jP���ŝ�����E���_Hv&-�M.B!�E0����U�ĒB2p�1����%d�1	�_^�.1�y���3BD�("bKH���^�ԓw���m廬dqҦ�T�8�:��^��Ȱ1gs�?/f���<�vV��j����9N4㈰<����������Y���ݴX�v�i/� J1��HL����1�2ͱV�m"U�m���f"]�X��hQ*|�S�E��Y��/n���m�}U�,�v��lR29**��P���ṓ�7h�1cs`|�\�$]�'��*n)QH����wZ,,nl�y,Z�l[�6�҇UA(�R�QD�E�}�Rǝ�����`y{u�M���(f&2:�m�3��p�1�vkX�r�L�-�4;B:"�R�0`D ��&��j�I:s�Ӫ��R�NH��ۮ���w?���X�������d��IEA�b��e���1x���%Z�ᡫn�L��41*�GM�9Q��JQ�B��;�ۮ���m��_}U��w;�k�BdqҦ�T�8�{v�}T��;���������}�}M����&%M6� ŝ���f��=	b�����Xve�J�6�D�q�u}T���Y��{v�a�o; ��6)�E*
�l�76{w���Z�l�76���:[���[7R�BwM��I���M}�63qM����	�a��zowK|�:I�z~}���� � �I� )�׍s������i�d�Ӵc6�ltô:�k������Υ���d�:�pطb�5y�����6z�f�&�ѩ��\��j֦!�4Fl�ء��W�)�F[
�qW8hJ��6�]kl,�ۢ9{c	�]�����FT�Lږ.ue�X�lv��Ջ6�m��mҫ�׊��X������� 3�4v��f֥G`�3e.6?F�Ţ@�$��wX��嫦�e�YvuH�,I���Y�e"]3�����մ6\D$4��L��v*I7#"�)���R�<����ۯ���<����l]$���Q9IX�\�z<��{��Ž�`f:i_W�$z��:���)D�����`|����K7���5k�3�J��f�RQJ��w�W��;�����X^�vT��y����7Q�I�F�`}��VDl���Z�l�76N�~��֫Z��.��nۖ2����[CF�7&īpFhV�us\��Uf"35*r����,�v���`~^�}�UW�Μ����[�S��*%������][O��ʔP wwdd���t��\��/�rL8�!�K�q��B�	��mNl�)@�D#�#P�l���cROw���I9y�;�H=�͊FG%ER��)���`}��VtDD%�_M��_M�}Y,�$t܌�D�v�lԬ/f���k�������b� 4H�*�8�M��5́�[��́�Zs`to���l���չ�7%�׶h"]&�\����פ��l����ɴ�kn�D�R���������cs`c���� ՛��߳IGG)(�H��ۮ���$oO.�V���7ބ���7Q�I�QQ��3�.v��]����ٓ��D�$a�PϪ`�4@c�t,#��4S���$0Hjاr!��
�`ЫR,�}�I;{߱�?Vd�j����9MEQ�w�RǛ��Ž������9gN\����J�'E9Q(�v�n��������Ձ���`w�wo�� :m'Pq��ٴQ�b: �G4�[��fkf� ���jEt��T����QT�*
G�,�v�&�`y{5��W�Y�����e9#��dR%#�=�5����Hś�����`~^�w��Wԑ����@h��J8܍X���,nl�K�M���XF���t�j�N8�:����w;�{��Ǵ�X_���X��Q'�ʸ�A�xS�$�pn�6�>�2{6���Ӯ ��X���caen/=���ۄ�c���%'$v���`t{��wҾV���́���]�J��mS-�\���^�Qb�
��ZG*��t�Zncef�,F��SVm��e��v �u~�`b�s`|���>X��F�m5QJq%��G�<����ۮ��cs`c�r��{Б����
���D�D�q�Y���ۮΪK;g5`b��`�5�RB9**��AH�:��wM���X�\�w�=哽�`��S�:nFE"R;ۓZ�:�����-��́Q�*�8T�x$� ��(,������F�W6��Rϟu9ąHu�Ay�ߊ���R^b�Jg��`�k_}�"X�pɯ&^b ܰaI�G0vL�QJ$��$�d&!��y"F|E���YleҔ���C��Y��x�Y�$�� �Dc炁����s}��D$bm灐@> ����w���g��~��w\��h����� �A>@%���cÇ
���1XL͔�[�ü��!c93-͇4�w�{�a	�\6��9���x��
[���o`��7/⏾�t�37n�tF�vر���X�j��3�
	�������#B0�30`�s��!�C�,��4�x�hD9��$���UQH4K���hb�$�&���W_G_t�����c�����	h�ޥ��恱��@&rD{�����R:*��pl9Ѝ_��%e�>q�t������zv'��\37@ȷ�դ�=��R�u�k�K��@�1����m�bna�e���Y�7CO�ba[]x�%~���as^%4�<�ǡ�g��hf�[���&@N��R2=P�!��y��8��$V�                         6�@             6j�:�M)n$�5]f�Ǖ-k�n#���cvݱ��6k5b�ѱ��"�- Ga+%GC2Ҙ�0Xm�*�Ymyt��m55n�����].���2ܵ���;��	l���b��d��fue�fķ4η��M6��&-���b�K���&f16�.�t8���l�Y����"KJ����!�u� h� 5n��#vi��ؚ��5�����El,��Y�[,u���4�ͫz܆n���Ѹ�.#�hYqU�ԔИ�-�YaB�����5ic1�9Υkm�1]��Ee�3kK��,9��립q+[l�0qt���2kŭ5���I[�.����"&����^��t��2멵hX��N�V�	*�V�r�6\8�hͲ�f��Z\���0�1�(����շKl�vf�Y�����������3qkXr�cbjg$f�h�K�٥m��f�A 6l�	vp�b2miu�f�#Nel���6dj���np�c��� �-�GKY�&n�5����nՈ�j�(#k֋-��,S�,�GGD���k1n��4��T�;b�\���V�6m�4ά�����Mëe��$̂��D�Z��/��KY�;g��bے^�Equ$n���ٶ�iT�t��e���i�7TtK�B�l�%�4"������=6 ƶXC:]lm`chcf�1�WfR�F��$��5��[�Y��n�X�V卼�0�,L��m�%H[�Ζ;:�S�j�(�Qi5��m^vrמ��h��iu�e�9�q"Vl�)�v����6�ڵ�͖]De*�3f`�.�+�^�-��k�HW�V]f�S\��5����K�A�
6�X,D�k�i�u����5�[o�ڻ.�u�����,�V�nU�X[���hYu��X�}�s4����L��́\Pn�q�ͮ�T�7GJ��v��V^aFb)�De�e�X�0Ԣ��V`�3s�hj�دW�*�p
����|��w�8�y �������i	�r�<�V�_0��/�!��	�����W�"���Ʈ�X&��S�؇@׀���h�8�q�l��d0=<)���ڙ#(��<x9��k�!�C�t<7¯C�W�Oh ��x���&@��9���8LxG�Ýv�8S�b�hh�@ p�7�TI$�I$�D�  m�l  m�%:���jѢ�D��n��.����Jf�&�H��Ҡm��9��n�r���YK�h]1e�Bl���1n���KVʼ�t6�{���J����	i���Fm���P�[U)��pX�A ��+��7Z5�ض�M����[�B�v�eB�շA]�c��������jsq4I��фCX�K����q�L��Yn"d�ԉjU�J'K!�x�L�vLu�$鬻n{s�o.mZnն�oS���cqv�Mȹ�"�R9�5n�?/n����=�5��-�؉N�!��v�́����Ǵ�X�\�{�	�.P���II������`{rkVu%�7���������n��b��m���w��`j��`|�����9[������E)Ĕ"�)j���k�:=;�?�{��Ǵ�X��u0��&�6���Ѻވsi�ԮSL�R�GY�F̥ٺ�]���7*���vt�5?�{���cs`c�r�ވ��}6��tԐ�J��FAH��ۮ�}V���c�x�M�ؘ9�I��0^	�&z��+3����H���4�"�4	H�R�X=�BF��ʰ1n��>X��DBA���e9#�$DN%#�3�sV��]��%������`n|�lp!!IE#�������������a���K;o��=\��!Ӫ�diA���y��;�w�~y�J�1=s`w�뾶�؊��.<m�-̼rb1��t�3{X�0��vky�y�GVm��Tvt���[�6=�*����z>A�{���k�DPtԔTn8�nMj��H���`b��5cs}�BFCu�*)TIH�QE#�X�y���]��оOk$��1�=��LF��D��*4,Z
�!%��Ƥ��Ձ���ޕ>l)��vU�,����ӕa��[<�l�MG*9**�#�1{u���UVs������,nl����%Ԓ��4��2���S��Sl��͵���.�c�S����b��7a�2�}I?�o�V'�l�7= k{����k�h!!IE#���s]���|����՝����֯���H�s��N�!���v�w;�]��Y�9�o;�edZ�)�J���rGaԵ�s�7�t��6o�q�>�/��}��CrNk\�x��BI�a��0d���D	�V��!4Y��N�H�*$f����2�E�h�cJ	b�����t�=����J)�v=�*��F�>��Ž�`j����{������4r��k��n��ڸj���q�:�=��a�InIv���n�顦��*USR��w�>X������DD|�;g5`ec��>l)��v�������M���X����y Ǽ�q�9)��#�5gs�=�5�;ꪤ�v�<���V捔䎛�����u,�݁�����{u�uRם��������!IE$�������k{���:�l	��Iad�1.)��9�H��Y�I�۠�1�Y!!��\:K5�wu���~��UUUR�  :�  $�My6�qNҗd-h�Y�l[���7�%�ݦ0�L������Q�i��J3F�&T%L�X�Qt��l��2�#F�9f��v�Z�"4�Yl�Җf.Qr�P5����9��N�m�2:]������� gr2�7d�.iv�ؚ�W�*ыu�.��m2�M�ck0��d��G�ma����s�.b$õa30�13&s�`h�H�b5 �(T���H�s{Ż�1�g9��,��H�i��J��j��j�3K��L-�.L
��]745�e�-�￦�Ս́�u�����3�I��ETQT��rG`b��=�u��s]��f����=�>91T����8��ޞ��6tz����k{���3&��ȈE#v��������`b��ꪥ�7��2��o�%>l)��v���`uUk����Ձ幮��ع%� F�����M��6TΗ[��1�6��l�1�2�F�E���.�:1�MT��)�5gs�=�5��s_W�~A���6�xl�$tܕ$ �M��iʾ��B����T�LLZ��|Ƈ���[%��Oi��:J3��k	����)H ���E�D@������5!�ws�1{u�$v��tpP����U%`j��`|�����5��`n�rV�ו�48|�D��uR���`5��`f:iXw��y����֥D��F�RQ9#�1{u���J����`~^�v}K;�]R���ȝE�mPs����R;!��*[\��8^�T����M�k�R*p��8���9+�s]��{u�}���v�vu����*A��1=s}��D$b����34���#+���S�¤�����;y�cS)����K�&"e�5e��Z�+s�1�V�	d��ٕ��T��X A�%��
��@�����
�������t8��U*2
Ga�_Rם���{Ԭ-�vT����o��T��$ �v�:�X�DDl���[�6�nl[��v�ej�a��m3�X�<����42�S�
V�at:t�]q�tݚ{*�M�UY��`bz���cs`j����쾅`z��tMU$ҁ�v��������T뮂�ź��#�|�ڕN�H�D(ܑ�����M����v�<����ZF���I�I���5s�>X��O�0S7Fb��x�S1�wxơ'���}�:E3h��1���B-���`*�y��[�hd�dD	R�E���́�;�? ��M�����2��!"M�lVecmu�+��H��%p�%
����멦;^�ޔ�=ƻ"Z��q$����V76fӃ��{�����y��nT�N%#�1{u�}I��W>������8��̨��M�Qʂ���z��幮�����^�v�<U�D�*Er��,�}6-�V76�BݧЬ�����J���B9��{u��k��������f�9��$���HI �.�
�� Ef����@�.�y�K+�`<I�H�׿�� � �-  	gRƣ��f�u�k�s��9�m����(��{���u��Nu� ,L�WKLl��X�b�]�m%Z۳.��m���nf��؎&ܭ�*�)���Y�'fi���i',;^�1pف�������3B5�m�b�ؚ�`ٳq�F\k[H����	��l����to�n�I�[�	�"�DV�7kjԂ|����EX$A`V)HTݮ�F&�k��I����$h�E�#�K$6Z���m�[1Sn�ȓMB�����?�`fN�V'�D|�w;�.��H�$�N8�=�J���́����Ս���#��A$�����`b��`~^�vu}Ij��`f=�V��zD��0� n�l;��B�����3'\+��-}��ۼ�q�7�T�����6d�`bz���cs`w�ѽ�TͲ˥����%-��.F���ke�L��l�Rf!RM%,�v�6iԚ��v�3�����+�6�����5��`v��\�CEIPj(���<�5�aG��9���Ja�j�L�x�0�5.B��i�v�ɘ|L���_�*9���`���B�=�=�H��1wt��د�##��FҒ�*d#��Y��^�vd�+�6y�e�RE!T�#��Z����V��������˨�\�G!$
q���������>��Ž�`j����n�$�V� ��f��s�I�s�]�iA�4i��ը��	q5݇I�t�ӲGGe)�\�l�76�nlOZ�#�zD���*@����]��ۮ��%�X�����	s�UT�j	R�8���՝���횕�)b��̂|F0Ǔ�DKԥ	F_�n��5���X����>���0d#r(>�A��"�X3��>S++y�����P��OڒA�� ��0BY��9�<�po[��v�H | ;�=c����
}�r�w/&��/Q���PG�v�Q���b=L��O�Ԋ��>��E�؈Dl�	���,��>A O�
����@p�:p�J�e�Q��]J�dR-"��S��=��0��?�02��q�ج�����~
y>�l��ɫ������O��{廡g�~����i�}�@��d��/f0b���_ۢ ~>y*��v{=%�HY���>Ub����8�g��sJ�����?h�]��&0�эnB�.�M�p�n���g�~�|:�M����>��OR '� ��k�����$�d�1P����q�+u��ŋ;:��}�" ����?&�+̀`^,0- G���8�3�p��;�7�zY'W��\�H��-��7��rs��։p�CB�@6�§�	S&S��y(0���S�<C����|9z <MǞ�<xh��j��2(t�� ⯜��y^�f�a�ˊt�^��»@u:y���{�8*qG��CO�5�1�6'Tb P�����˴�#7è�:����Y���^�yMy6�x�Ӏ��x؜�:C%[�9��xG��M�C�6� 
D�0�0";(5F!��\�5$��}�I'OwA?�r����#��g_%`b��`~^�v_Rם����H�����QI�<�5�U_}��������J���IlIHS�Д�:�p�FۖV�V�zOI;L�c��f%�F6#2m`��*d#����]��ۮ���j]_�b��`g��u:j}�rG`b����tҰ1=s`|����H�.��r@�q��9+�s]���%���՝�����)ȇR��*����G��>��M���	�1}�q~��m�	�7�Z��B ޵����C�'ɾ��˟��_l�cJ}���!iBZbj��ĥ��\�� ��ٙ!�\��b؅X� ��-���rV�^��)�tT�7#�?,nlX����V'�l�����m�`ܫ�M��f��`���.\���2�^�$���nF��N��v,��W;-5���1�J���́����6�'�S�TR��v��R����#o;�;���ۮ���H��H�J��5RD�?,}��,�vuW�}Ij��`ft���ciIT�2��:N�M���M���`bz���7�R�MJ�J7$v/n����:�/��Ϧ��cs`c����<��<� nO��dHu"� C���wA~����J�x4�>g�b�(���` ��  ۤ�  �R��U��$�4��o*3LBZ�f�0i�sf��;Z�K	���u�6�L^lˆfXl�ؤl�%嶢Qi.��L��F�d�Iv�(,�ڗK�eFem�l)��َ`��n��I����[ḾS!�m,�]V6�SW:�5V�u��H:.M䈥i^�-���31[����t�e�[Il`��HkẌ�c�i���5]E�@ߤ�I/wY:� ��V�� ַm�1�!q;P����on������+�#�� ��p�ѹ��st�4�M=t��Y���3}@�ι+�6����5��`n�S��"J�J��AX[���<����������IX�7�IO�����������gWԖc������~���Br����uTBs��`n�p�O\�t{�'{��v�'�S�Q%A��y��ꯪ�����w;�]�ۜ�%�% �����pq�hB�ٸ�0���b͝���LMD�kF���4&H�`"��->[��M�����Ս�G�� ݞ�XԺ6��$����qo�;�j�'޿'9�ma��z3�J�'�,�J=\g.!�h� ���A��P��P"��ɋ���s�4V���Hϻ��*t� ��ʩ���3%�Yބ�s�1ot��Z�lQ�I�q�a�_,��+W>��͇{��s��`n�U�D�)D�D���幮�ﾯ<��՝����������GM���'`s�%����R�n�m��n���nn�6�mx����D���*@���;���ۮ�̖����A��M�c}!T���̀�R;�]�Wԑ���`b��`~^�w�RA�����9NHT$�����ԓ���5 {epZ� $R��J}��,I��;~�ԧ�0w.��4g	b`�*��(R*Z!E`֠(�ou�j,�v�<U�D�U%A��r
þ�B���`b��5csa�[��+՝FҒ�*��v���`w�Z��1�
����`g�jJ6܄Q�Ǝ�Y�0AJ��ebt�5ic
$)p��L�:n�7]��a��+����u��-�����DG�>A�{���t���#��8����诪���]��,�v/n��H̭��S�a*Q*B)`b��`~^�vuWԖ��vc�����ޑ%>n���vK�;��k{��̖�ap�}��ޟK.0���J�Gv�dIk&-�&Bh `;�R�uLg6&"���e�� P+H	Q�D�J"An��w����9���������k�_��M������{���.Iu$�n�ɣn	�k����kvɜ&��16���]Iqr��m'���\I��;g,9��n�p�O\�,nz>@��M��%��"i*���Q9`ynk�?/n��]��=�X���Ғ�*��M�����Ս͝�zݞ�X����wK�:tԨ�%7$v�ם���}°<�5�uR���`{�uʎ!�$
����=�X�}����<������/��Ue�H����[w}^����9�n�ϟ[� m  6�` Z��6,���\;%��i�&����lYa6DQ,ŕ�*;4�T��]e�ap��mKñ3��iR1�j�	L�}vDN��S���-U[�T�*SLe��n4&*4�f�?�'��ys�\���72�kT���YYf�	G�h���Zʈ��cdȄx��m�Xd�/E�W��f�Qڗ�5p:�鵴�2kj���&m���X�X(�V(���Q��Τ�m�3���n��2D�2󶱪-�Ƨ��
7�u��^U� ��rɌ:���;s�E%��~_����̝k{���n�p����x�)�tT�7#�?/n��Y����+�s]�~���B��JG`j���̖�gG��	j��`b����l�c�R�vK2w
��Ϧ��csaވNw�lq-G)�2�IPj(���<�5���w?�j��`{�5+���y�Ѷ䂩)�JS1��.;ur\��ně�J%��t��멛�k�:7iG*�CR���Y��^�v=�+��D|�W>�}��]11*���7$v/n��_~>�tpf�V
�ۣ&�Ip�Z���C�>�p��3>��J���+�B�PK��k8�`T�!b,Q��B��1=��X��z��cRM�n�ꪤ�}ιW*��r@�q�κU���;�	b����3#j]*�S�P%HH�V�����1{u�w�;o��2��o�"|��uS`|���:!��O�o:�V'�l/��}�k����3���jL�f�n�l��R0��K��
�PY�;��J-���J�lX������9�Dd�.� 7��ک$��E�G��Ȋ平`|���5cs|��%��4�R�!D�9�1v�?/n�?��~�:MX��VM�;���ey�h��P�~@#��D�s�L�K�����Yy��B#��)���^��ԓ��}�jI��ϱ�(�P�%*���ۮ����`{^kvKo;>��.��R�%)8�����>s�f���́��s`t-���n��&���n`��3b��60�n�Յ�h"�f��a	�Չ�[��555?�/�lO\�,�6�nlh��H bL�n�u}�;����<�y������}_$ec��D��)��v�o;�]�_|���7`b��`�5�9�i�8�:<��t���f���̈́��(���22N�w9>��aq|�A _� D�1���}�I'{ߦ1�RH�(���?k�n�着�����o;�]��U_V����rQ��a(j���˝՛Fm.5��$ΨV�M�Ӵ4��YM`�2l[0���-��￦��f��5cs���gK�#z�jE�D�A���{5�U|��;���{��[�ﾯ�#>��.��R�%!MMM���M��s6w��s�1k�`~�]j�P�*9T�8�:�^y�M���M���sa���9��3a��(��:�T���幮����<��k{���cd�D��F"�PB��I�[K����×����ł������{�����}�\�ȒߞL_!n�о�D�Q]�/>�����`Rc"T �L�$�Ӎ������ ("PU�b$C�b��KC^[Bd�H�	'�	��1����jC�FU每�6xvN 4�H�S&�w�4
��`��lx�7C��@�$a�L��Q_&)� o>7��dRKFZ����b�0h߁�g�#���y��8A^$��� CI[#�g��@0��1S��.mG�r��0^��J�������>��Oa�n��ߣ���P}H�o�
{��	=%��� �����i+|/ˊ���A �H�/K	�Ab5 �|y��K�� 6z�����0���߂)��
N9\��H	_"�q H/�`����@/����ˀ��;��$#�����va~�pY�a��g�v��X�����i@�b��|#��hF@1����ٰ�Ho�)�7������UZh�}e����Es�V,���eNW<���Q]��R���_��?Ju�����)+�_S[T���A�z A`~,3�������D��I$�@                       8 �             \�S��Ŧ�0�bRe�vK
,ƔYrͦ%N��Q6�i\���mX63bk�\*�k��(l=�3\�У���F��k��o�>m��	ue���B��y���]fAH�քL�k{Z�VgB���`Mq��ݭ�������a��\�M��3k��h�
v��<�z�v�a5��8�Ge&�L-���Q���u5�J�[e���K��֖ۖhF�k�B��uir�BQm]��fQڸ�%�y��BSC*��i��3M��Z�a�	\+R�(�i*SҌ�b�6� 1.�YHk� �����W16#]����j��1���	`�GR��#na�;��D�bT#/cr�l`&0շYN�j[�`�Y�&n�5�o��ms*jn"�
��cFT��6˰ІY^�j�:\L�h;M�M�MI�])�ޙ�m$ɛH���t���^y�ԒE��6�Ѭ�-��V�U]�����.+�s�)���X��9Y]�`��Z�5���mj!�S,(;Fb+l�0���j�պ�^e4͚��T�l�77�� ���+m괘mmaư`n����J v�ْ�k�f(T�qB��ubM�N����mRm����ز�,5MZ�Ė��*V��h���4��G�-��cl��nI��۳mі���Q���^�!6,Ηk�t,���*���t��՗:;6���F�V�]f&��ٺ��``,�
-�J)��gu�K�G\K1�v�&�j˘cR^�2���l�Knc�34�k����ҥP���6��m�<�|�w��r�5�R0��jit�+k*٦z��]���f��V�%��]�M��/Y\�u�i�tM�q�Fع�	�0���<�y15�b�A�/H��,�6���2�$. ƌ�i��a+��,��3]�R,�YH�Vi]�/.���]]*5���]�k�*��Q�f���V�C�m)P�n͚�P�p�����e!��,#�6�CN����D�ê| x��$M�����<9������`!y�Ã�`<la�^F��BO'Wt�/����4���jP�Q�#����/Ly�*Ca�|�`A8�|��8��<�b�'����]��U3�r�W�"'���6&<�D��U����x_-|�ƊyN�ߐȏp x��x���ڙ��t�'t���O'wߝ���|UUUTT ��  ��s��\b�4�ĕ�:���ں�z�M�.���n��cj���F��#kn�B)�l���[��8���`r:��`ݒa�^�#`V�F�(�A��ManK���+.��R�Xh��We.�f�b�6NY����$��Xl�m��)���ݖ���#k��l�a��ޒd�:�uX���%ܝ=�D�7&q./!),b�`�C'�yj�۲E�2�l�)��'�i�uY2K��5��qb�����q�jVk�P5S�|�t����>X�6'���fk
r"�:�"N;�]�z1oq6��X,�7��BA���$R��2T#�������l�������`r��`o��N&ҩ!ME�
ýK��1k���áf�p�Vt]�B���ےX��]��;�?�=°����yw4�RIl��a�hWSFi�лc��mQ�I�n�RޒCbj@�Z�4M��V7M3��s�Zr��>�lV �]w��b��`g��*�
����H����+�RU�>K"��1�b�!��B$X$A|z�H;�Ձ��s`<���z�#�[R�*0�T�R
�;w���{5��v>�`{p�W�&���B�(m�,:�������}����+�����ޖ^���EIE:�"SS`<�Ձ�Kb�����f��;�7�?GM�(t4:N8��TB��Zj)�\]0�Ћ0ܒ�-]$N�)e�6�iI��U9Dd�����+ �͖��������X��W'iT�����+ {����$b��`v�r�>�lWބ�Vt]�B�)Q7$�<�y��O.����,�u��w:���a-	��>H��I������gYr膈�J1b�A�E������9���l�=���:t�%%P����y-���`uՇ,�|�}��W(T���IV�=�X�z!s}_�_M��[VD{ٽ�/�i"��v:y�:ls,Y����4iGV�p:���ǡ̵-݇E�μ&�Ύ!U�o���n��Kk����A�{�`ec��QShT��%��fk��D$v�r�1�r����=	k}!N�(�D�vc�V�{�ΪH�ޖ-�v��62H�9Dd��ý去��s}V-�6=
1YI1`e�H�.VS�hV@�Z@,��H6�!��D��N�rD"A1P��x�,W�$���q�$�5NE`uՁޏF�}?�{���e�`~��߿x��M�un�s(ծ ��vuη
�%�yZC�r鲁�(�v�&�u�d�j��3U_����nl�[]��zX���d��d��i�`j�뾈���sܬ��1ks}��$g��*�
��qR$q�`f��`������`j��3+#�U$%J���R��D%��X��l�ڰ7]2��y�oj*%&%NQ�X[������]���q`uՀ몾��TLfAy�t��
58B��3�MO�C���,�5��ׯ�O{u����  [@ �&� ��N6��KM�u]#t�f�F9��Xf!K1�=X�9�4�h6�j4D���.m�ͩ�jl�E�.�+�e���р�][b;E�˚]��0R�0�\��+a���K�=l�cq�ٷ&�^%�J4�u�r^� �z�.�YJ���*�X^�掛�:���*m7#^��ku��=��憶k<�(T�fd����3e.(��Rc	��d��:m�ݰnU͸�۳7F�J�2�d�3�VM�et���dm�x^�/c)���(�Ev���`f���73g��U_�j��`��e9"t���N+^�/�o��k�M��[W��BGu=G'$iT���G!`���Ź�����}����Ł���lc�U
��Dܒë�;�������ɥ�}U�ԗn��=�i��'E8ȅ�;r[VD{������5cs`s�}mm�!�:�5���|�n�n�1�3B��9�`�%�[��i�{W�^�$FŃ�Vi`���`uՁ��� ��`fV�ԪH:R�pjE`��� n�>��LgY�&�S�RgWU���q�۝i����& d�3eL	)����cRM���I�c�W�|���S}Q|Jm*p#RKVw;䶬�D%�/��s}V��"h�IE8%#�ꯗ<�vs�V��,:��;��wo�䉲R���ls�X�����l�ڰ?��D��v��$���R��*�l�K]RmLm�.��.K��҃)3],�S+�+`�*��X�u`j���y-��|�y�+՝F8�P�
TM�,^�wޏ$v�r�7�������F{��$��dB��������y�ʰ����6&G Gȇ ��D��_�,h��&\f�o��nsrc0���59�͔�^��x=$�i�!\F=�vFY|M��� R	`�j:ĀFFNТY����I��y���Z�تJIϑ	$,;���gM�`{��Ս͇DB�wŁ���EH:��I���g�e��W�k����Xך����ݜ6�F�o�*�W6�v!v��d�\�+�9�ۻTZ�Te6��uM�!Q�NjI�Y��=�X�Z�G���`���+�(�D�v�&��RFs�V��,�n���Ნ�7�8X�����>���Ǵ�v'PԒH�I���+�������I�w>��2rw�J���A�9�@1��J΂���Ȉ<b�jyz�|7V�H0dH5q��I>;�ϳ���5B�)Q7$�ٻ,�����k�V�ݖW�Y�}I(�rD���F��5pA:�a�X����Rؖ]�1c�(��\��vɸd��aN2!E$���8�=�5X�u���}�`g��(:�UBUD"����͝j�7� �[��/���#2�>�RA�d�NH�s�X��YވKy��|��Ω����j�ԒÒ��K;g�y�þ����[��)�}*P�@�K�,�t�| �����VFz6zѝ��`�pSܗ��CP���~���� �  m�l  m� X�U/���.�p��5�#��6t�	`�[��hJ96�`�ME&.���׮�.Զ!�T�t�ɚk�x��m�l3��,��&�u�S]�m���E����J`9$�ܣ-��m��2�/�o����G�4�٭4�[LD�-�]�
m]r�z�p���j�sB[�6n�6U٤-��3�4V�F)�}��d����,�u�l��ǀx������g0�g��띲�4��5�����3\Mu�\��ԚGX�C(�NH���r�4�?��`��`�6XܚX�yKFI"U$�����n7W�=�A��Xθ�>ݦX[���R�"
TM�,�f�۴�;��K�,�uXy��J&B&2$�#�þ��Y�|XݜX{vX{6X��Z�تJQ�H����e�n7V���{L�.;���a��ښ�+nxF�0Ga���˩�X8�X�YcU��H��\�îμ&慷%TѠ���}�V��ވ�Z��,R�����Rm�p#RK �͗ﾬ��u�g�ɋS0Q5r��fR�Cd��U϶�Am�y1
'_����y���t�ъ�v"��A�!G��A����gS,q���GԐV��
p�J�8��`gl����e�	{��}V ޲d�����1�$p���U�]�ŀooK �͖����;)�s�H�*HE��z����y7�_ ��7L�:7~�o��!dR˙\�s�έ�I�P&u̦Y�a��E��˙]Vl���b��U| �uX��`ct�� ��X���d
q�DrX�4�=�4���`����#�c�TtU%F�BI;���,�J]VF~���"\�G�@�4��؋����|�$�gcsOx�������{�R��>��Lj��iK��WQ:j6.��V}r:PU�L� ȸ �o���%(�Cۙ'pö��)?�5z��m��Rs<���y��
N���&���!��FE�n�x���g�����$�9�n����3�BDg�߼�/��x��&_1�Z2�8�N��V��E}��<p�^o��G�켁>�@�%��^�n��a���#�7�g),���ɢ�&�%���M%�SNgGI�	�Q 9�5z�gQH�|�?;y���7-7�t�������Gc+7�g�8w�'�B�PĮd�X�v= �A0��䘇߿v~�|go�	˹��&���{�����e/�d�n��Y�=��lA�����2Y�+�
Mv���3_��� ϧR�t@?���9���od��O�#x��8�@q��}����%I�a��`kQR
�A�iu|��ED��>!�0��_9@�}��y�my�߻/T>\6o��NDz]�I��(�}��������4̤�ݧ�#�T�g9;���jh������+�?J�D�|J��Q���Ĝ��~�2�� &<�8�HB�N��~=ss{h~,�����	��}�������~	�ݬ�]���s!H�6��*tr�O#�I���p�G��HI�+�0��L�|�����g$L�w��L�:��&��<�Y ����x�<����w���^`��8�:&����^�����<d��4�z�y:��Thi<}CÇ��@���4���=^�|�ȅ!�����8T�	$:flrݯS�u�"&9˽��=GT�  �b0bŶ]n�ۓK�Yҩ �2D'�,q�����Ǵ�����Ł��S}QT�4�"#RK �ݖ�&�7L����y+RL*��DJ��b�TҔG�(d�&\ky�<�M��1�[@*jf�)S��@	Dq�ܚX�&��ݝ��_~A���;���rD��(�����4������`yn�=�4�3��GL��D�j'!`�u`|�\����,�\X��%�*������Xw��/<�vv�,��ԟ||Ie�@��1D����! 3�>Ґ��f�2KCﱡʹ�e6[�aM��p�b��A�����`�o��u$�������Hb2$�JG`{ri`~�M,=�,�ٮ�ﾥ��.�)Pl��l������6�X]��ɱ�E�6e�ˣW�4���c�+*����� ��=�8���?/f����3�q`{k�U�$)N$�#p����""1k�7�q`}�L���=\�7�JM2"5$�<�y�ܚYԗ��+ ��Y��)�} �J�ê��Y�|XǼ�=�,;ﾥ���;��ʒF��(����'Z�:���Z�l{L�D�HL���,� ��x��!�;#�~ư�@��M��3,1�[o^�/��� m  �� j��5�l��r���::�f�[":l��k�q�h�vKG���*ԚF��jSm+vu`V�K�u�F2��X�v���V�LV[��i���wR��thV�nR9@�]A�tMmc5\�S5�trU��4"E�eLT��cZfZ�dͶ�3�Z��c�s��-�9�����5c�6�L3$�;)f]�;Z˙��\R�1x��D�A��o<��m�V���J�ICT-��0S\��f�%E0k'N�`�fu��u5�6u��&�R��`�~����Ǵ���{�:�aқ�U%FDܒ����o�=脍�\X��X�u}���:��DH�����Ł��5Y�U|���,,�v���6:��q�(��,;гi�Ϫ��f�������u_�AҔ�I�'�f����������>ͦX��rK�$ݔ���^��k�7GL�Y��q������].n��n��/q��^u�k�s1�����Z�>ͦw�Ϫ�!��)�} �H�ך����:��:&��$�L��
f2F�7��2L�5������ �%q�
��)��=����nn� �n�꤃�k�*9r��(�E`f���3se�U�������Ł�Ou��jR#�HȜ��f� ��V�֬:>�,��\�&9T�U�K �f�|�U��6i`��`uW˷�]R��*���ڻX/Kck�p�!==e�Բʻ35�@�T�֦�K� �SR��E$�c�V�d��7ٳ������oK�c�A�J�$Q*��iXf�/�	k���`<�j�朗=�˪���IHF�`���&��gS�q
sal��!��Ӹ�3}���3��D9�9���F E��5`���q�]I=߳�ԓ�牽��RT��Tq�`��,�Ƭ�i���DB]���!��R�U1T@���y:Ձ��f�����`��,�w�?GM�(t�N��� �l�.6����K�-�-[RPumv��vP�����c�Q�ӔF)P�?�{6q`��`��;����o;2��E8��G�"���k�舄�5�X���f�/��H�gE�29T� �NI,۽,�\��cuŀv���8�h��JQ	��WԹ��=�8��nu%;L�|̓`�t�R[!!��h�Jtf��V�i��XX�yL>���jS9<��'h�>Ǔ5��4��D(�,F���p�@kh��Lw��I>`�I�9�F����4�?��v�O��U��[Vz3_$�IUTQ�-f���S,3+n�iA�hݣ��� �hB�,ͫ��h��p*H4Jq%!����`�]X%����1�����jg��T%���K �����;�=�8��l��� ����} �(�K�_+��e�H�}V��X݇0��i�%5*5"���^ݾ,�zX�͖��=O5��j}�P"���k����|l�V۴�I>{�%ő����3�\�Өw@"oh�T �9���I$�I%�  7|�~|  -�@j�E�Q��îA��n�ͫ�Ǯ��f�솅�qؚ�lrF5�ƌZ�
6���4�K)N"D�v��#�s���s�
�8�m˭潋�:�I]�����f��E����I��ͻ$̮4��8���.xjc���	v�+��&��e�t6)	�s�d�l�ʉlf��-��`���=c�V�LRc9���G(D{�@��N�'Y:>x��l�`��U�f���ST��h;:y}IXu�.�Zmn���DDu�U6⤢rI�}����<�`~̚W�f��=�V��#aIJ"!��y:��$f���;_U�}����H�c�Tt��9�G#���l��7ٲΪ�H��K��+��T�*H�9IH8�a�_/>�v�ޖy��d���y�Oj:��60��q��͖z����q`5Ձ���7m�6��I��l�9���6p�궎�0�l����s�ۗ�n���vt��Ҧ��;e�>ݦX�u��G�o��;v��㍧(�9Q)��7n�{�=d���DY-z��m���HG��V ",AB�}V��� y���=���>N%>�D()*�;7��g�e�o�e��sn���R��nEB��%�z"z����X=w�_U��uo_�4F(�5$��l�;���g>�> �}V�������J�fj��-��>��>L��I��f,u�s����%�SJ����7��l�
��ŤL��[�����k� ��_��k�3c�tR�NRR�V�͗�UIn����`~�۫���2��O�BRT��UMMU�k}V �]Y��mEA����b?h�.(	�#�B����$��B�/�6K���Dق�4�� #"$[Tm��w�RI�ΖY��t�NP:s�9,:����}V>� y��;Ж��`��6��P��I,ٻu`w�.���7zX�6XU_v�D��1�b%&�Sh0��ʥ���K]l����1�;hT@�#�����R��1��I_�;7��f� y��=�}�C}jR���7"�D��=������ �ޖ����7ض_U}I��ޔ�AR�#!$�X��>��,�V�����I�u*J�U�K���Y�#�]V��X)���y1"d3Wމ!@���;K v�c�I�Y^=�C��9�p��x�ג)� �-I�˓Zq�t�ݕ�dd/B^�:����m��>��fR���UD�TX�N�7]Xcu`}��<������o�M��ۑT�!XJ#m5.Dɦ�4h��7=�����v��f��r��60��O����=��`~�۫ �Ų�+=��R2��u!B�Xcu}��� ��U�fk�脃y��HӔ@s蜖����71l�{6X��,z�k��)RG�*��脹���7_U�n7V�Y�ߪ��n�����1ȨM6I,ٛ,���/{� }��fՀ�DG��W�`(*��DW��(*�AU�

��PPU_� ����T@��B
����� �@X*R
�"�D
�P*P �@ �DE`�@U*@��b�@E`�@�� * ��*@��`�E�V
�D�������������� �D*
�Q��*V
�@ �@B*�Q*D*P*E �EQ��X*Q�� X�Q��H* ��*��
�`�EF*�  �A
� �A
�D`�A
�E �@A��@��D��Q��P �DQ`�E��
�b�A
�Q �@V
�E��`�A
�@ �E�P�� H*Q��*D��H*���@�� �D �D`�E �D`�A*�*H*
�
�X**H*� �A�� ��
�`�D��*� �@������
�F
�B
�*�
�T���� H*��*��H���*F
�@����
�*"�D*
�����* �B
�H���
�*��
�
�`�E�� �� ��
�R
�`�D��*��
� �@��* �A��(� �H
���H*"� �H
��� �H**���*
� �H*�� 
�_�AU���W�V����PU_������W� ����U�H(*��AAUx������d�Mg8sR�	��f�A@��̟\�7|`                     �              ��*
E(�DRUE
�B�J 	PQ@R�R�(QP�I*�	KX�(P�TUP�           z  @    ��QP�"��P0��Zxz<��|�}�}^l{���������$������ʸ��w��|�����J�g}0=�'�[��Io�� w���'�y��v���@��y��ӽ��<�"���S��>�9��;���}}����ª���n��
tq�%I(�)TU(�p�	7w^{U����ί�}5��Ư�Z7��W�W��=�;7�ڨ}�yï}c�&��<����9P�\������Ƥ�;m�z|`g�ǟg�|y�Q_G�y�����}�����]��<��$���ۯA������ہ���}g*|��{T;� �
@�P�� c�������|����;�����O�����|
��g�R�%�������g@�|Ϥ�R�A�IV�R�l�z4��t�� 
	����|Ɣ��I���J#�f�:�X��=z�=}��;��OO�ϲ�O@;�E6�)KL� z(���)OO��Gٔ�:>�(��:���@D��P((��	����ѹ���O�����JYo�o`<�ς�����<���|��7`.f=�o	Uyk����^��>�c�����zD����)%{���u��ϣ�0�^GRw��yꨟf�	����S���y��ﯸ/���v}}��[�z
P�T�A!IU*�p �
,ۀY����O�� ���U}����0<�	�y���g$���w3�`w��ѣ� �w� �ן`w���1�#l��}���`x�� {���p}>�|���}�.v}����_Wy����C��OSEM�T� O))S � #?L�R������ �i���5R�z�  5?I�3*T���C�
lU(A14zj|������8_����Y�9�Nc����3�@^q� ���AO� �������X� �����_O����Vr���0,x�G��b�Ω[����s�r]����
|�^G�7[��'�\���)?NӖ]|��&��/oiN4����1d\޷���k��v�6p��& c|�C�gJ�^�F��	ݼFÏ����x�dbN�B����F��q�`�[���x�O7�q΋w7���xk�E�5)I}0��=|�B�&�]� Y���M�{�d�xM�XL޶ݼN�'��J�!¸�zp���t�!q�ȶ�9���>7WZ`�v�����^�\#������fc�ֆS+��ɵ=Ƶ2�滇hG�o,�SoH�'�T_����:d_p���'�y�M����=�0B�u����1
`��S�;AN[� 	뼹ff�N�b{�=�ޞ5�����9�N�T<� �M��:��p���T�^�UF�
����.n	��T*N�]p0�H^T
q��s�������g��e��K�`�:ǹH[�n]f�=EG+xv���� ��8�zb�=��+o��$5��#�>�Sڳ+�mm��'������b�i��ʏx�s<,�Q�u���f���i�	���h��<�8��:�Q���ot\&�4y�&}e# �$c5�Y��+�zA{s؃���t�����I>!˙&x����3�t�z�n�"����M�q����oM�9�M���=;q��Ue�uwx�D}`�Qy��bNm�����Rp�`�dH\�طbܺ�V������|���`s��r�z�©%�-�P�)���֠nAn�qfk+�~�j ���=��CZ��Ŋ�H���Wk8�a��܇	za\#��.%�X��͡P�����n\������VFa�T�Sl�{�N�Z3�����$�������#B�Y{�����]��bȯ����@�01^a����_n�bk�M����U�ʆ��.�r���ۤ�f�#�ؙ���m��:��x�/�{�������q��g*끼�qr�yt��^����]R�2��h>�x��lW�N�)1fW��`wW��[Օ��Kk�ir����Vb�x��N����f`bIkyEk��7�m�ݐLD��&�˰5�Oh>�x1�uzs�+��a�6�t�����Σ�O�g���]ڮ[<u墟b#�3�³��W8>��-�7ߊtnf�����O�.`�;A�ct�3���M�>�=�8��<����7Ļ(�px���8ucJ���_�W��"���9�R(&I�@S�B{A�q+��x�>�|W�ڂl;�<��',x�h��hB�{�e����f�@�wm�S�?�����=�TV�!���}�1A{��x�m-ܵq䠝	���>��.��$�uk�5���5fd	o`�o�(�ĻO�3���,�Ȝg� }7}��7}� ��d���	�/s�c�]�
�HRe�a�E�s9�k���V�i�郼]��x�����n��B��
�o����H��A�4^͐��3�2-����(�Y�#�31�X��p��e�k#{���f��-#6h�4I�&:w�����<�]����p7��w9P�{��(
(5����	`�e�N	�1����%a٠�'f�5m���!3�������Ё:�\^��t.駊�@��pٔ�0�u�&#���tvH&��s�=Π���\͛R'٨m͹�V�cy�Zn���8#��v��o*��,)��)絘�7T�j}�t���W�{�w����[�8k��<0u�D�Ģ���<Rxܰf�\�p��뫰ig$x{��:?`�VcoR샮}�iܗ��Q}�w��돂|�����5���3nܕ=�l�ۇV��]��۶�ķs1T���fb���2+�S���1)��c1f���.dA֓7:ֱ�+�2����w�;�����i��q��!C������nGDs��)��9�Ҽ������"���H-�I7e1!�#��j�6�_nvnnq�	�۹���9l��W���!�q왞:�ld�x��:LN�m~&�c�sݦ�,{��<�`���L]&�t�t\��1��@:࢝�V�Sv
]�;$�TZN_vu:Чnh̴o��1�ؘ��32h�{YE��k(��W�-�3�'t͙*�˕�#��T�3��Mh8TOv��{r��և/��
�9n��K��ˣP��2k;���l�t��h�J5�G�feYH{��M�z�H�u]�}�N`97ݷ��0^^�+ڷF�EocT2���5�8p�c�o4;!�Fn�-Y�n�Aq��\(�cXAL�Jy�41|�j�]��S�"�/Y�����[�*{�zicZM�[U*��ٵ{!M،�u����gB��*�(yJ�q	����pNP��-�aHvB4�0��Ѫ���ѥ��q%�;�%���Z����<Df'�{�љ7p��{c�c�r����j�vv+ky.��!kU�A�ky���kq��(m�x��(��w�$|-�{�!�Pe8}��a���`0�C��;0_�9y��BL�ʞ۞��
��&��=��o1��x����Re�0
�Ý�B7�ta���1�+�/׵)ٍ��Z��ݏ�um�A�H��D	
.5.�!x���m��{w#�sx0}�f$$�P��<|�>$�Wo�J��:�O�c��&��,�A�3'���dמ�S4�r�һ
 ��l��������tx��s���ˆ���`q��^�`̷���w�C'0c�Sfo��I�J4˻GE��=�7`!5j�#����S�^�V���lݺ�\�Bc�I�Vcр�
�沭�]�qf���;�M/Jk�D|�33`�����<)hó���m
ݕL����|W���/�?!x�I�q敹�X�I/!�pH���x��IP�
��� ���� ��O��q*�$K�\$!
ּ@+S�����(�T��
�7�!&A���e�0�YN�����qb�f�jf=k����+2������m攃 �`�*s�#S�1��+�TT���9�m��ރ��g��C"�U]'��y�׬��;άe�d���kL�9��߰i��4ݍw�T��o2���J(`�3�[����ـ�4�P�FN�f���
w 8QF�v�g@ �)����n`�9�nc�<5��Ijg�5baow�����6�x{�8�=����ì��`������+���,�%��N�� r!V������nQ��������m�7�K8�`_}�}�Ǉ���t>����y���u�q�祼�-���$�^e1�{Y8�Sl���s��B����/���]�f"��=��m��`͎e9��.����J��p5�N{�^+9�,���˳L9�hÙd��$�K8�>V����sg��fn|d������@jc(��+�d<b9:yK�å{[̌Rax���ru�"��u=(O��3x��Mf�Iź^�3���e�V�w\Ϗ�]��ݔพl�εnZ;GI����[��+��32{tww�' U>�(����xl�=�`��-�3��
�Ef"F��GN�p2�z���Z��펄p�0#�vpo5V��� �}�X��i�#u�i�;ڮXj�n��{xz�u�$}��3N���`�|B	�'�\�^xf���C`�I]����س��b��MJ��Z��� �kV�\
}Q�P$���؎�m�3�	��!4�����<��g��� �!�D�$��
\���-| A:;S��R��Ƀyl�{��D��I�$�xU����o���	��KGsK�������(gM��7v8�Im�Q�,�.f��R��0K	����"p�3^�<3���ۇ��oa��N;v&�Iɨ�
QY�6<�tu������F�[[ȷ�
�l77c�)<�x�j%���w����N�
�D���{!t���
��R���3W�5���
}��D�6Z�n��p჆`���]�)�oO{��w:��s���s�Xh���n�Nf�P9�w���\f�|=��F!�O��>Y	~�Ƥs��
�7pt�Ƈ	�u�H-Nf��{�/ ���M���YO*��ss6���M83iۻ�+v�g�a')t͝��>%b�QN�A�`�����g_�g+n�|9($�vf��k�5���AF��௜���7/,�-.�Sm���!Ob�{x��q�wݼ�F�|�yL��R��.޾A�@�;��N�YGkj7�}�2���D�˜��ޝ�.�2���Y�M�td�rVN�ٝH,�Y�.C
z7#<5%�g�'�0��/�A�-��b�=N��G���*z����ٽw�E�t6m$�E]�a�r)��;���KV���SNR�`���Z�nh�
d@'<Ɨ�4�t�v��[}pm6>w!܈7w��Gk���{	Z�d�ʃѴ�mY^�3Q��g�:��w���{�ޘ`��C�K3xB
Ow:�E�'b�zF90bUj�)���pM뻍���C;��g����8cT�b���0��S|��H߳���=�p;�����p3����澳`d��g�,�;��Ԭ���rmqֲwn�:	Z��㈌��@Ȑ�!T��f�z�P42��G@��Y��b�f#_��Q'�hB�VGx�6�L���'�e#��+|Y%l�P�zqu�fu����wj��Ǘ�������,D'�m�6nG���&�ɫm��n��7��ݛ*�&b/����*��l"��}�4E+͊ug�]��xV�%��X�1�q[
���	o������6�>Oɧ��=�M{憗��-X�l'�CcϏY�Y��p��/U��p;�����f�1�pѭJ����,����Ib�0}xDҔ��ʸ���[�+	p�S����c8�π ۘM���4(#�d�376"�V�n>&�"��b�}��s�3 ��5Uj!f��G!FT�f��n��#�ՠZ�v@@�=�\��I��y�p�Jh����v�������=�v
�<Χ^���7��.���^���\�n?s�i׍yy/r�*!<%;�}ᬒK^-��Le���C�N�\sǪ��󀷎 ������>�C<PI�si�3�_1�P`��ưG(��vp6�
%�*G����|ƺ�;&71��s_^�W2YUY�f|Ryw�|t|۶��З��c���&My��4q�J��E�N-�sV��2��O^P��ef�I�z��Y!DV�A�1���5��A�I���,���ߜ:݄e�r����z��<�� �Wŝw����!����8�U��I �rnT(h����$'♠o�|
s.$( !�:h)���;]��CިvգV_��������x�
1����Bx����A���w����3|S�
�,��cr��HOd�;�׎�����/�*Ѱ��/%��׌�+Ji��p��P×���)i��AA����4s���Am�IT���l�C�W�ݝD�`4�
�0�ť��3����Y P��2��-� +E6RX~"�	 ��Q�����,r���u�Qu����ėE86a'�l{|m;��LV����p8w3����PpT��j=⍀��k.F-4 u���zr9��i[0�ޝ�ksO
f����d$�P����wO^��|�>���B�@$�cBW�/�BAhH�;���>]��a:/�rH
���3�Y���(�]չ�&f���w��2�:���z
rMѧ�`��E��i\�M��3si�b���C�������\Wڰp�/��љ�'H�k�P������'+G7�AyJ�'
e�/��`�h7>���bvm����9��*����hg�>:��{��(�u��Wd� �xت2�]����Y�����0G�zt�f���'~����ov�����||K����t��o0V��2��&�<v��5oiq����4Y[��2(> �ˬ ���x�+8��q��RW�JG�|�r<ZLCu*J7�%,����|'��a$����=>�W�&}6�)�`i�+Ӂ'<^j=.ɧ�VB�m��;�u�u.gi[�Lc@\�&M=∼��·i���6oZ��Z�ޯ�$�KW�i%�r!2)	�0j[�fΰ�H���t�!<��
��&>D. �v{iU�	`�^�ķ����&�Jea����x�N�K�GI��$~�؁L���U�k[i�->�;�{�M���@	��8��� �G�Bq��ԁ|S>�u[7�k��(FvANK�� �����<���t���-Wɭ���fWӹ"���=0|���3<v>�N�'��6=b${Vsvs<9��B�y��3U�ʬ� i1C}�I%UUUUuUUUUUUR�jU����������UUUUUUUUUUUJ�����UWm�UUUUUUTUUUUUTUZ�����_UUUUUUUUUUUUUUUUUUUUUUUUVڪ���j[,U�7��/�bƠ�7@��Y\W )v�a`���h�W#�F[�荸�Z����(�ںX��yՊ�n�!3΢76����`u�3Xj����Jcd��]�2�3f�h�v@��J��&��"F|�׭0']�r�Y��^a�ɣ	�,�c2�ŦfCB��	I��R�Lac�4]4�Dj���^v+lH��7���-�`�W'@]M�gh�����H�{���ƛi���Y��Lj&��tl�@1�ђDM�q�>C�&w:g��\-��{87��l�t��2��2��:�ä́=��"��j�k�m�y9s+:%�J�g�w�w\Ց�F�6�Z��f�MW0��Ɣ�T�KV$��g�Е���h����ca�H�a�]�W��e���V�BkH��-�:1�{OkAǆ�hڀi��730K �#Tm1M����L�b��5��ԕ�  U��l��L��V��[6��<v�L�L/�5·��,Z�r�Z�Y���Y5Xd�5�ѷi��% W(2����2�ٷMm��UiQ�'��A,���������.�4�����U�F���u�؋�Z�E��Y0�	ƛl&2iV��#������(��5�;!�EVx�͖���qT�����9�ַ'ex1ÌCn����CV�em�u�(�BM�Tcdg�f�H��h���h7�=�t)�mu1�Zu1*b7m�� ����B X�F�2=��v���؅nѼv8�\��d���63��z��ν��ں3��ļ-m%5b�Ù��!l�؀]s���.��0n��q�N����v��-><��e��e�f�+	��]*����&�mI{a�g�mM].9�*6�3���$&M��mm; ��Ӱ�\d��%�w�7���tMԣ��
6�R1�g-����,��ѹ̍s��օ�!ͷ8M��4�&:݅ݭr�/bvƺ�աMڄ����ݞs.���TTj��k�,���˭se�'�K�; ���ʹ�@�Fe1�՝�������W!�n�pUÝ�Wi*���\�jz�'P<��k�׮ ��3eل�0��UR�=M�j�sռ��"�l��̄��;\��:�[�q��Ϯ�.C�7�� �۰�Ŷ�ֵ�HQ�O�����������Kb��q�ʴq�v�/SmM̏�(���2���n�%�۳\8sS^�r3�ᆺ�m��.c�&�ʓMi7�H�f#q��'dp���.�5Ϝ���\';n��^v�Y���6��6�9��x��&�k�J�kK�,;F�h<F�;:e�{%̈��WnS���n&���7O;$tCG>��{	�7n�m�Y�JF. ݴc�w��s���ʝ�dZ��a�R7۝ؤ��qB(����3%��fs��c������γլ�Riu಼θ&�6�
B�^<�[d�Q�2�v1*��T]�'�tl@����p��vv�/3�"�3���Fj�z�^!5�Y�n�Z ԰��et�I�MYo������q���s���/��k����V��a�������vf�72��f�܎5��5̺����HCU�ֵ҃D����ވmH�<�<%ӣ���e����Cg���Y������t[`U�	[���Eu�?/��U���0,�˂gR�prs����i1􎶎6��ڑ.N9�z����tZ�1�M�&܌򙍪a��]����GY��-�l潃N�ܪ�8*��7t�����0Q�׳�p��^��Ǎ=�ϰ(���V���8��v��h�#q���a[e�簚��� �vSnֽ�|	ׇ�v;g0�H{l3��MmZb��۞T�CN����'A��Pp14�Zv���em�\h�]Vl����J�=\����<��G�am�cMUJ@t�z�:�%�x,�{S��<�sOa��J��/k<*A#�'0���,u/bvr�Yu4u���s�V%r��zN��=����GJ#����z���Z86�e���%;^��_�e�q�xۛN6�f������ɷ;��7-�� �u�^H[,�*ƒl�:7X�k�"�n��f���qZ��8��V�I6\(�.F�;�P�Ë�Qx���es�'>p���wM�%ɫ�J{m��r�	ݣ&�s����L&�A
��	Q�1ʒ������:������v�ͦK����%����j����=��,��y���ǓtH:�k��`W.75:	����;e�^n$���*k۝�q�rbh�탚|�t\�Xn��|��]�l�,h͜<��%�6]i^M�&�ge�kv���b��e�G�NW�Nn��6�h"��s0���[T�6��v,������YAZ�ap�1����D2<iɂ��������zU lm��\b�v�2p� �=���q�IU+���e��Q�v�;.��9ը����C��my��ۑ�5�9$b�2��k\���N`jY��g+�3X�-3�n\��T�	��m\�gq5z,��q����69�r[��v0�=���#�݄V+��[��Xwm��*k�Yc�c:HW��SPf�Sa�#�u�Xoh�{-��ie�赜	�ؼ峈wl�w��|G���nIϞ͵\ú�9�p���j�uך��`���G8�GB�Iov6i�P��������,�A��\q���g]o�?�8~ZP��w1�k{r�a�n��5�<�n�ݜ�68��ۚ|�5]��[�l�����O>/BGS7m�.���@�P�v�n�� �)=�a�-�Ad��Xx�:C6Z���kmfM�����j��hiCQk�in�yc qT#F7RjSf,���8� '%�>3Ө7<vƸkG\�MKJ��f�4p���p��Ku&\�pB�P��pL�vݭ�mbm��4��xL��@=)+sO]W�+�I�́wB2��4���0k
z�([�@ݭ���WWS��c����t�x�F���v�kuC��1�H͜�g��]�{��q�1]�Y��I�V7nZ.�7#��wdn��S�i��h�Od�U�ݛ�O7TX�Y*�SJ��(Ym��!�}_UT�_9��}�?��5m��J�@��6`��X�bm�!-k��q*R�LY�Hz��uk�6ԇm[v�����.�eUp-�A����-<\iZ��^�g]A F�[6u[GcK�6p/���pvU�	M�^�&�<1��n��53���U309,fecN�J����ґNc���Z���i�w���T)v+��{V�kN��]/h�"Ţj���-�q�� ��m�	Ӛ1���@<J�d}����AՒ����,��r[W�C����,j�
CY��Q��f։
Y��Є��Be`�+��5�u,0h=�h,V�إ���=�#��çׂ-s�ۣ��B�7q���uvͱ`L+-Z	r��יd�`�<������'rm��YU�b���;y<�m�ҶS�9�,�Q����`�ݝ�9Z�bc.�Թy��ʽlA]bK	D���6]m��&��#��8i��Z �L������W��qT��,f�ٴ�8�#����YI��hj�3Ji����3\̂c����^Bs���9�ձ��).� �&f�V�-#�0����^�飃�tlYx�6����8s�]TV6��Cm��T&��̄�Ƕ��9s���2��2t��۶��:�o2�2��rŖِ{ۂ�
�iI<,�+]��M�\"9$0(�pB��Oyv�fv�[,m�&�B0/nӺJ5�J�t�2/K��,']�Ps��\t�p8����p�5�=�<�1t�ayu�Z:�"�n�=�.lpV��Ρ�8�<��\&�v�cuV䓱�D�p�N�-�M�>@Gm��Q�۶����;B�����t��@��V͕��:�thL�:����8S.ݍ[v���9��k��+���R�N[��'&��8�\��<�y�2� ���X9�=m�,!�ZK�[2X#���ճ#�H��!ڥ�Ņ� ܆pK)6�:�P2�;��h�����F�̓�!���vB-�j��.`M�,V�۵Bŵ�=4m�R�Ш�a��8���w\��ĺ:a�1�(�#��Z��6��S�).�2�v^\��l�B�1M\ό��[�klcU�(�s�eS!�9��.T-��[M�eX��d��؋/G��7c�(��4��K���W��.Gv���,�P�m���"�6"x]n�c�M��$��հ��� ��65v�f�J��5Yvssg���Yɳ2r�od�I�9
�#���c�C�{.�0=;Y�-q�H<��n�	h-�%��.��pƪ�z�!	�b�h�E��kPe바�����X�ɹ�$���)���������:�;:}��Wd��u�}�����p{h���1�`ɼv�#��Y��fU��z���S;mIn��:�n���#�s7g1�&:;gD��n9���%�8�0�:8Ւk�:���c�[��Ƕ��-%���\m	��� ���P��k�ˢئ�!i4+*��%]���b�� �Հ���ݗ�y��,���g��ڕk����m<C���y��1��4+��SR$�L)dguЩ�-�L���ܲ�E��ki@������ݾg�8�v�v���v�.�A�v�����ǕJ9wc&�x��G.;c�
�v�.��V��&뜀�m��Ҍ��LcMe��6�1����JJn�x��u�ܛ*�5p䞷n��b�����B��!��+/�z�n˩78k���:�4Ν���ۭ#p��Yn��x�����F��_HXz��z�a֓vݛ��ۥY��!vu�c��lk�����-�n�X�#��\X\Vm�z�a�c�{]vh!+��da5ͧ��&*T�N�G&y�V3�.�su������YfZ�:U��u)m-.# cGVP��S;8w����Iӻ�}�GeCq���/�a�I$NB�@�@2H?�`A��+��C�5�T���	�"@�AHGa� �$G���g3r��0��~>��RS!��6�n��	1x����*W0	�4��BO�~ࡠ2�F��b�44�����$�T�Da�$	1d�1A�`@��<Cʚ̉�L��XJ��R!D��\�"|p2!��xD&g���I�?
� I��SS2I�HJ/ ȜM?�Ⱥ�hFmM��ф8�d$�2�$2I	�q�	�5tS�̐�C3q$�2��Q"j���E�rl� a%�r2%
L�IwL��0�B�[0�j!����Jp������$�'����2�!4pNy��H.�BA��0?I$vՐ���If�Ê�4��O�!"��
���$�;��CH���&�lG�H��!��jIɀ���"!'��dX$�	D�4;���Ә>?���N��t�p�.d��[k��`AҫJ!H�a4�h��VI%��t?��p`�9� HHE�ۘ��CbB!�$E�C�!	�?I���萋! i��H�>�'���� hP�
Y@aaa4+�i㿷�cm(c'#���3*Y6	���ןH��1%h>W/$H0�~�𴄓����lL���O�����S�O�?D�c!��!e8@���D�'��A~�:��$>�3
�D9G���	I'῏�m?�ms�ʿ~.��#�� ���$%�1��2����L�E�q�|;�B^ĒN��FVd��g���qr��+ VHD@?�E7�	 &-?~�Ȭ�%aX��KP,`Ǌ|��7q�ar"d�d�2�L�Ql�t?�4pn�k8a$$I�	-�� D~�"��O�Ȁj	Tx~�?1N"�ec @d���˸@0�@����9�I!�)M��6�8B�'�� �`�� c�` �� ���� G�@�%] m�r�� ȁ"� �8�����$t~��bp�B� ۬����H,�2,��ICm4���BHD�HY$G���#8��
Yai�6d�_߬��R Hm���� ��!!"8� �ȖHO�&6B��$#��@4|�L�����V��B�PB$�$��tf��9�5�IQ���c- �� �$�+�;��Y �0�$ � :n�G9�lP�1�C�<U΀�A2��		"L(`�Ć��?H�(�E$X@ȿ<�O�)�Il�`�g��H�<6l!?Yi�0n+�$��HE�C"|;7���(~�$� ~'�1��dP2'��^KeR~�h0�C�$KK󽪼ݴ����1a�<��&��1�6_��A�%B�W�N	cI �D�'�H$a��D�dg�H�`��&@*3�s�B�'2H�$�"8T��$$M�x��Uن�I��u��ĶXX�ၰ^$OƧēR���HIa�Á���&�����S����q�0����91 �����B!)��X��1�FC��(��D�m���ߡЉ<BG㌰C���!��
�u"!�3�E"	oC��{v'����L�g�h����	a��'ژmm!:���LQ\<�r�*�b����0d�!g�$I#6BH�H@���	��0��BD�6����"�:>d��$!8�E���H��}�BD�F@����9�[i�%��<~��VBH2}Ɉ�4���y�6Z
Z�JD���2~��ȓ)����p	s�$ HB0!�����$�\0I��R�@|�+#�1� Ѷ���%А�qV�t�3��b�$$$�Hd?H���n�#h��H����0�mvXH���>�T��!	4ig
@?:@�dm�HBHو�d�-bS@>��A�A��	�@	����":@�p����Ia�'�!Dd܄B���;�ȅ�"d�0~!#�!
P��� Hd���R`D��!��SP�iGy؍�l!o&��f�pp�?!+(؄@�����/ a"�$	HE`M'�Z�?B�QɲrY���(o&�6d�8 >H�>�� �������Y�RA��#b�V��&���`��|�����N��?���b�@���`4B�����'�0dC���%�a �H���0bR�v��H� s)I�je��FV���U�͌/%���I��B(m��!	>��q�X�eq��h�a��[0�(~~����l"`���`�n9�T,ԉj�@l?��2B��ӕ?f[��ld�	����	_ĩ�Đ���$�ԁ���?	��$a	�0�9����H	c ~��3*݀lxq$@�'?~�򆹹$� �"^C0,(�$3����gy�O��H�^'�&i���B$8 0�H��@�[B��Y��];�$$�������~ Wl�@��Blh.U��l	 �ْ��(�dDh<fIh0��,I�d�ϐ��eB0B�I�F$�r@̖�@٬�dD��#�� B(d }�O��0C/�l-�-��>X���X?B�Ѫ}$�HM�Hp.YBC�o���������R0�!J.�����$¹O��� i`E��I�­HB0��WL ���ĘlF�c�`�"@J��
@b@erG8'��c���%(��R|�2D�4�҄d���R2D��A��w$�!# ��H�����*:@���,"6�F�J�����>�L�9�9�TcUV#=���*��UUUu,���a�qt/!;OO<1�
ir�ÔzP[��wcvl�-<<.�OJ:9���qo赭��q�c����5��fY`�"�bT`��Y�	�\��l�{mMe��F���%#30������Jk��67Iٹ护]��5�9�q�玱r�ێ��k��ēU�a�]n�]���،kf����/Z�.�ۺ�V)�s7C�۔d��k��{=����Q�;��N�׏j�$�%��G鶉� m�مD�!ٰm۝.MY��<#�@"#��ۃ��l��啇m��86��r�L����jmc��jD6��f]�0�>5<���9�};��b7iZH�1��+ƺ͖�6�����IQ)�k�X�^3�@]��AX�!Ķ�2���ڐ��[��v;q�x@���4�׬�s�P��6�
kNp���;��s�l����"���ȣ�m	�v�Z:�nf�7���챃=\�<�Ƹ���s:p�"P���rp��\��ڒ�b��l0B�
�&�j�7�N�+j*񫮷y���x�:�f�{vG���j$%Sg��Ξ(�ٍ�.5�֒�P�Zࡇ�#�m�����ם)k�W3��3�Ѵr�4��E����p�Ӹ��Z�.nx=�H�9xcNu�`��.\���������������Ԍ�vث�����	���,tb^�l�Xa�B�n�����v؀����ݺ��9����v$������W�k�v��x�]s*�h��\�Rn$�W6^dIm�h�X�Vb�.�8�ˬpZ�q�[�]�= �\9��x��J۰p���7)�Y�Z]�Ň�Ve�dwlk��lH�K�V�e�N�֫8���S��ўӮ���AV�S�m���E\��k+4f����Ԙڢ�����k�w ��=Mŋ�(nz�T��V�/��6�;�\���E���t��L�cgm[��yE^�i��"��7�uٻ���v`���hs�J�rZLpNL<B oj�㣍����>T�8Sp�Q�����>8~� �I��urB1>���U
?~W�N����O���4�S��$J 5��U���} �q*L ~i���Ǌ`�����~~����B�?9D��! B8Hq��(��@��~4XiN������� 8�(qr�&��>U����)�Ţ�1QfV"G�3�u���J`��J�6��T+��2�GL�R�h�K
�)c��$���M+Z7��E�Sf҄�d1P�n�#���9Ĥ$ʠ��.�;1�v(����	r��Ns�s�i�O=���.]�؜+��W�����0���Y.�Hu�Ĺp:̨[�+m1���%���Rg�N��6�8��%J��[ ҏ�v�p���U2��y�Q9񝲇�=�۲v�nq�N���:gI#P��a`wޔ@>�}j���eXc�ڥ�����r��t_�q&�nm� �͖���ߨN�U%**��IE���Z�g��؈Q3�����ݶX��'.ptR���NEa�s����=�K�̺,7�������mC���T�I`{�0�7�Y��Q���V��KzN�~���j��[R&��9s��.���.�FX6^l+��sMƲ���
.�Y��%(DG!���E���Z�g�o��y�́��۩N%�M	���L�>�e���LĪN���xA1�B2�\ZHG5m�WFk��e������s�:�}��ԇ�2�{����n��D���T��f��ݬ�f�q���e��ݵ`��n�E*���J���&�7wm�s2Ն��nmX�ѵKiS�*;32�`j�w���6�z�����A��%8钢�Th� �eۘ��¹�ꦶ�gJ��z��;%h�΍q��*JTUH�%�ݵ`c�eX~̭_0�ݺ,�T��2EQR�R��2s��b!B�2su�����̵{Ē�gr�Q�:h�D"I%T�n��f[,������)���Z!$&�4ͅ�a�L�D�sd�d��
|o`E"o)�,�� (g�Nڰ<��V�|R�\%G
�]:v
�72���ڰ=?f;�r�u��:��Ĵ�47R�ٙj�،~�����`}��e��u}�/�Q���Z��+�����=���g�H�k�ۈ��֛���8�G5"�{�V�fU��f]�Ϙf�ڰ��YUJ�qƣ��<̫����e���j���e^��a��mR����E*�X���ٙj�I7�۵`c�ڰ>YHx��RR�ʪr2�y�'���1�v�<̫L�:�:۸�%.p]�ƴM��%�]����2��F��? 0S}!X#��k��,ԓ���uM�2EQR�R��1�2���V���nn�,fe�W9���uKSR��ⶫ�`�7,��[F��Ѡ.�#��x����<y�:�ј�w�0�*�����Ǿ���e���fZ�1粬��*�J���Ӓ���e��̵`c�eXy�W��ُU�\uQ�i��J��3wmX��VjK���ڰ7wm�a�p�؊d��tꕁ���`zs1����\y��+ �j�:�(�'j9*���ʰ5sۻ�>7vՁ�=�a)�l�5��LBI&0d�cI�T�"h1���-�3 G(B���Ƅ���% 
�x(<��Ltv9��f�c��+�$�M���:wjt{(��mv�g�MϬ�
b�4n�Y�bʼk����cg
�ISM��w]CG:���ZlWB,,!D��t������4}�O<�YMiE�*瑰�[c�jݞ�N9ڽ�V��2A���y.�WH�p�v�nN�q�Y�VTB�pm���u�"f\޻����\f�vqL�BOgv[@e�����3�ﷺ��qg���'�����X�\㶲�#����+Fګ�C8���:���v�JRcY6���R����e���fZ�2s��?Hd����>Zь	z��M9S,��W�B�6w5�;���e��q$�;탪oi�*���:��o�j���c�33-��2Ձ�<�n[�N�B$�*���q'�7]���tX��V��o}�,O'��I�䉒G`ff]�2Հgs%���`l����o������#ĺb$e�؛�':�^[�Eڮ8N)�])PDq��=Z�YM������ݵ`cﲬef=�_0�ͶX���I���PS�VO��j-�W�'�cZ�H�)�xb���:*�9��o�6��jO�3��,��6옎w���4�JD���H���|��`o��e��̵z�d0ŭ��T�2�*U��[����]j\�y���~ͫ �x6�b�PC"nB�TN�o�X������a�����`ue#hZ(r�$���fZ�5(����n֖��l�5(J3w\����lP���fLI,煙B2�5��Wu��;v�ӝ�J��N+��!��;���fL,g��ߘf�ڰ7՜ڧT�t�R9*;ٓ�ٛ�tX����������O5� �5U�*��3rm;ٙj�*�$����7囪M̛p�6xBQ$@_�����$H�4ē9ƻu��;s�j����8�)���N��fZ�>��;ٙj�^n^Ӱ7MۄUB%(�J�Xe{��f���7&Ӱ=������t?1:Cr颓��)f�r5�@�*`7/gE�lr:=��.�����E$��Q*?��ݵ`{=2���̵�K���v��ƫB�*��D�E`{=2���̵`}��v�2Ձ��'�1�IJ�)��;ٙj��+����n�7&Ӱ>�A�V�TT�Q%Ea�.>��v�vՁ���v��;�^^���ći�:�C��������1FBI!#��H$�!qj���Vz��(t�8"�rTv}�j�ԗ����ݵ`}��v<3���J\�U%:N�Qz�C���/[-���qǜ�q���f���{D�ZJT�"t�/��ɴ��2Ձ�W��K���V�n��%E(�S�;��V�^�`wٖ�g�S�I6n����j*$Vv�]��fZ�R\o7&Ӱ=���Ǔ̀�)%5)��lDD�7+7+\�{2Ն�Gvf� �ғU�8�TȇQX�L�`o^�ߗ�wk5��e�݀�95{��T�j��w�.�����Ns�3��z��9ľ_Z+�����F=���{�}.�4IB"��/����z<wp����`��!ʟG��w�=��<�Η��|>S�zG>���3�H�q�;v;-m�iƬ�
��-�a-r�����m�WV��s��y9��p/h"��Yb����@��i���$���w%�2�=��=A�S����X�z��<��V�s�B�WM&�"� fщ��Lf�͚Ab���N��=�{^L�Vod�5"JAݵ�GSGvK2[B�4�fi�щ�,W��3.B�ݥ����Vv�����W�l�d�/HC�(BY�y��Rʞva�pV3d���p�b9�4l�m*u�u�^�1�4�c��WR��Rj8%Jzw6Ձ�W���e������t��ND"IQXe{��=���ܛN��-^�ēf���ht�8H�Tv�vՁ���vooٻj���k�:�yT�rEO�'N���$����v�vՁ�W���e�<f[Rp�T�j:���2Ձ�.���ݵ`{=2������j��WQ��]ˇ3g2��p����[=��f�n���[FÂ*���r�W~�~��v}�j��ze=����vՀa���tE!Q�U���?fޗ�����0OT��ˋ�&~��`�*Y���y�̓�����X�K�q!��Y���������nBL �������Da�B5W��ɣ�!��8�$#���r��}2����-Xe{���a��&�JqUTDM�X�6���fZ�>��;�����7��**S%Jv�'���;����L,7��y�{N�����IҜ!D���W����oO��ɴ�fe��H}��k\�Ve����-ȭ�ڡ�(�Z�t�x̖��������&rU�#�Q�mn����fe��K���v��7���"���J�=��N�&���Vv�]�癕z��f�mI�QR�!��S�3wmXe{��	�QaX�+�:�R�s�mJ��
��̎�c/�]����]�jD>K�$�oַ�}{�y�R`�`��n����7�VJ֡W�Ot]s�5(�F³��w~���>e���9����U��Z(#ᡉ		��S�mOOh�1��՗j�g?}`�A���}ût0ۙ����Ph��@��z��������I�g͂��P��q��l~�A{�~��������q�}����qk����C�ޯ%���II�����P ���HL��!-��P��I����2vޛ]͇D�lg�ĤƔ��J9�T�Y����aS$�:Y�,�%���_��R�v�!*��؞�������KaV�������5�]��a���yG�w2ak��K՟,��V�⏭]�{�o�@�4F�[�~�o�>��0�H�ݦ��#ʓ�:�>����t��5u�ӵ�[X�[���v��1I\�=���CYR9HU{;>>��ϯ�NK�����U����> ��w�*�L����7�z�+�Cl�j��o�M�!u��VU���B#�J|�3��yb	BB	�D"3\>�7�g�5�G�i ���h7�|0� _����
N
����p0�����J-Q�|@�������({8��.�QM���}㫽TۤmU�C|�#�~	 �K�R�vm]`�|� �0&�Èp%8'�a�³'�r�C��8 �N?ɭ�c��H|�6<᠚�L��� �pp|�҇8m�s��
��8�S���4�2��2�����8h FI������ɑ��Q�ء�t. ���kǜ�H���BC��"��r�i���5�`�Uȯ�S���~�R|hN!��i��/��x~`#����
G��;SA�p|��,�:�w�cRN~�e;0̸ET)ESQPJ�Xj\}ٚ�{�V��)�o8�n���0��`:"���)T��<̫W�^����V|��`lB���7+�uH��c�;כ���x����=���d�%�3[��P�JHRj�N*��(�UJ�ܛN��fZ�3��z��a�wj��M�D*:*S%Jv�2��f��]��wj����v��:
�C��B�E`gk��<̫7�\ow&Ӱ7wmXu��(t�8*��Tv��{[�V�M�`ffZ�k����q���ĸŷ8~�0�=��w  ��Q�����q7�:Y�Bn��H���1�!�4
MT,[&,�2M�a	���_]�a���PRU�'NJ�3=2������n���7՚�?y�3�.����|"L$�7UIƆ�Jr�.c&Z�.V�W&::zu���/9X[ux�d�GR��ffڰ3��v<̭I/�n��v�p������:�X��M�DDL�;��ܭs`ffZ����i�{�%��'R*iө�:{����sg%�wZ�;���cB�Ni6�J��a�9�o�s`wwZ�3����ݫ�Rڦ����L�)���VB������6{����s`~�`��z B�Ҙl�4`��/@#����Ћ��P0��{���$�_�l�d�3�s�<<a뛪���<rX�^� 9�<nQ�<�.�f=��:��7G]���=�j��M�ԁ� س��#�-��w5T�1�	����Bt,v�Mpq�1]��qήvM�/]=8q;�Hw��VK������w訹k�o"R�.�ە�]�����eH��7\��oM���֚��sb�&J]H2�b����	��[m	�.���(�@$��>~�mg]y:�S�sp���0�m�����%�\��t�Z$��w��'1ӥ�y�����vg��B�a��j�;'by���hST�:�ә��t&��s`owZ�3��䣓a�N�ӢJ�d�R��M�ݵ�lfe�:#��{�`o>�=�+%U@�t�"UK�6�'7w�7�6lfVB\���s��޺*����5N�X?{��
3v���V��=���������׉�87Vn��.#^C���\������a
��%**�cd��J�`{2a`fze;�̵�q|�_�j�7Ѝ�����&�,�L�/~~^.�@�i�⠃���*M��"%��L@���}����nl�"n�o�].1l�!gߋ�6�RFK�7dd����^��I>�v�����tB�l�ssĺT��c�%:s`n�Z�2~�;9.P�o;�Ձݵ�l�<R��X��(eS�a��Vo;;�Ձ���6�!rI=���'�.Y5E
f��:vٙj���.���~w�Ձ�������~�Xȼ����b�y�(�XF�b�4el,{!b��i��mM�k���Lҫ��R��/����6��j�����.���wu�7��U@�uQ-9t����-_B�l���g�g;�Ձ���oaG$�ݳ�NjFS%��5T���vٙj��W��\ix��OP�H�_|�8��QIޱ��:���YHB\�}�Ҭ�W,������e�l�^��i�J���+��&,��y�0H�HFFB! ����~��O��S���'�#�P�(䒿���s`w�mX�NeQN�*iԊ��t�9B\����X�\����-XtD.�����`���t���@�S.�����6(�n�|��7���fZ�:�h2L�j��9K�$��&��3YX뚺t���Ylf�b^&\�3��|n�3f1]�q\��m���Ձ����{2�G(���v�9�=���8���(eS�`d��w�rJ3{�X�\���ٖ��(K�DCgk�%���P�j�ӧ`f�Z�3=X����M��Z�:sy�NӢJ�d�R��Jâ!t(���������`d��v�hԭ9K>��QD�p�e����R!cHl�	��K�%�~��=U��UD��ӛ�fZ�6��ٯ���Vg�S�?s�qn���ԧ&99R"�p�i.#d��x�x�x�t��D�ִ�hWޒB+�aL����	�@��U��fZ�3=X�.����֬M�ꢪ�Tت)��N��ٖ��!G(���s`gwZ�2s��t(M�r�!>
SUQ,�K�`v�s��̵gB�Q�Oo;w�Ձ�*��T���Ӓ�9��]
!�w|���v��jã�D>���lk�-97R�SE�+1�&��Q�[�������6ٙj������?D��
ՍR	+�i*Ȝ��>�����0��� $|���l�*́��=Rr����-��nHכ-�y�y։���.�ͳpr� [\ۃ�B�9�������FR&GcJFn�rU�4q�,q�h�3�8��M\��,]�ؙ6���=h5��N��gsy�zM��ݷk��u�v �����t&jM�5E�M7q�� J�V�!�p�Q9	�ٙ�ɇ���<}b�n��GLִ󲽥T��PqV-�[�YiI�L�eB~� �)6.��1�t�Gg�\gԽ���-�d�����h4��+n�/_�y�槉��3��:���lmvb\e?���Ł���6ٙk�(�����; ���*�P�"d��3�2����I6owZ�7���̬-�Ԓ����&�"9'*u)����e{��s�$�n�,͛N��^ʰ�B�%(Tꕇ(舄�Oz���������e;\�8����X�d�B�lU�uE����`w(P������;��X�V�/MNJ��H��L��s�r��;p��;m�B]]v{�R��u<�m�t��6�Y��ExՎ��m����fe����%Ϙk�ڰ7i�� J#��1Ʃ'������7��G(ٽf�w�W>%ڼ��<�!3ZL�,eF0RSP�%	o��N����7Т#�DD6{)hq�j��tP�Ұ7���=9����!$����6�u�<�+lln�L��U�K�B���w;w�����V�B�O{q`����SL�:rU��d�v�q%��ߗ�f�����ʰ?.f��'R�2�*�x^�q�.�<[=��i䙙f[+(��9���W{Ӻw>>xE��痍1����`{=XX��|�(��|�w����y�9(�)�(:�`{=X_BQ�%�f�w;w������a%��jBB!Ч$eHX�v�{��T�aNsO0C˂`>��%�n9���� )n@�!)O�mwFV��$q)����5�B�$`$A����!	ǩ4Ә�"�r[/J�[z��v�����o���k$0�ϊ1��S�}���`wei`�9k(%�@�T�;J"�ͽs`n�ڰ=��V�B������s��4KT��dӒ�9�+33f�m�O 8�}���m������o9�� �~��t�|���t1���e��[����2��=3n�!�jl�N�]v��I���]�
�t������76Զ�o32}�nsc��#�B_UL�ww�����mtZ����Bs�� ~���������*{�ϱq�m����{��Ϲ�:�3��{'����.GKVl+�����o �y͛��>s��w�3�m������o﹭m����Lg�=�=��E��}��>m����-���̟|�S�Ý��J����$�9����r�x��R��!}�!	"�z����6�����=���P����5�����p�w/����X0��A�r�P�� I	�a%5�1�83�@�D~���k
y7���Ŷ��ۮ�D
%���H�����Z���� �}�{?}m��3�\j�o9�l����Y|��ZmY�t�Y���&Z�WJ�k( ��t2vs\f�f1�L�iY�N�1q�j�#�]�� ߿~~| ��?q�o9�l��S�m��gV�o}|Yqo��^���~| ��?q����Ӣ��{�7�m��gV�o9�g{��U3���~�Ηh�;Q�s�����|�[g>���#�s��{���m��3�\j�|�?a����i�����������;�:��{��;ݶ��1q�o���Ͽ���|����-�CM�0Ans -���w�m� ���b����w�ٽڑ���T�P�|>o{`ݡ��1�}��Uu�ؽ�7�ܕ*�j���#�bTΈ�"s��?��H�C=���/o�[�}{���C�<p]C+��	�])������̋{��|��v��,ň���,���E�*�R?8�,��]���p����(W�'��v�$q�H�<xc�{.��?a��v_��wf���Ă
ҹ"��Ǘ~?����g�������}�L�G�D�$���B<�3�R��Ч�ER��2�V];��B�w�`�*����!C�Hc��j�o��3����u;ӕ7K!�I����}�����Y�(��|���>�t|���EDB��-��v����o�ժt�j���[u����b��@�s����������Bj�All.\lH5n�J[D1)��'��?q���	�G���'Đ\�z�Y�����C4�0{7��pw�����>3��EI�
���	�\eU��J+T�a9o��QNw��p|#	��)
!�b3������8#�q:o[����۝����V��$����;�?����GNyE 	��*�5��B�I�&ϲ:��!� `Y0S0��";ANͻ��7{�9�PP@��	�r�ᝀ��td�>H<`�@�O�h��dU@UV�UPQ�@]�UUUUUb��e�4�&�9�����b6,sk{Q���1ҙ��b���2.nVπS������=-n�Fѧ�:�:�h�zۚ3W%�vL����R��O8�P�y�l��X�2�j�Y���Wf����0۬��55`���^l�E�n�(��$,U���+Q��dus��H��0���S[�v�E����-�6ȑ��睤�H��1v��@6�V�	e3-f*D35�`����$;�8�GL��Լ$J2�Ɖ��#I[n�@.�-���W+�t�����lnܽ��Asv�8�^�s�Ya��i�v�5�����LՀT$#���lYuW�����n��k�1T^��ܛ�}�.��t�fa���h�&(�k�e�Dۥ�L�!��^$m��ʯ����3۵�3v�G�92��YK�p[F��*�:��$-�5[��C\��t��Ʈ�z z���xZ��6��A]Sj��VS�tH�H���٦ٛa��f^��x�_�ŀ����r���[j|�f^6��ی��PԊ���vx�X��^� [<��}�_c�ndŋ_=�n|\�ѭu�7��[��H̐FhǪ����5w	��8踭�y���V�5�]K3o\��-I���������39��4�<����rd
���9��`p��ڱ4�y�m�!�Z�4.l4Д5M%%뺗G�OWk�`}s^�XSWM1FdCK�Cb]^�����e��n9���ȷt��0�%��òα��4[��t�֕���Q�E<�k��
��I˷��hgO;�V�����&��0Y8�M�	/�q(���mpJ͋�-��3l�XS5��l	i��8���;W�g��by�J�b�r\�l�J�&ja�y�$\�;6-g�d��x��H�y��^��u�m�3��R��)����i��A�m8�cֵv���n*Lg��u�؃.�o�N�al&{�<)�_6�M��X��b8аpg��[.j-�: :�lfgl'v�n��_�_�q0�z���������q�Eӡ���?qx.~�ş���?|� &Ǐ���������q7���2LG�T0���B�;2'���|C��h"l�)@�h�?"��|Q~���|��	���a��\���Âq�ɑ�?!��F����U����`
2'��W��&|?��W���hD���"q�W/�|8�S3�j�f�^8��܆��Ik�qۘ���ڋk�;s
����\��r��c����رoa�3��4z��(hV�yW��;A�2CO]=��^������m�@Aɑn2�������Cm�T3ļ��q��������b�K.���� y)u5Ęa��d1���k���v��t4$m���x��v�sfz1�n���n��6E������10�3����dEEC0�@>  G�z�9��u&%-�1��B3D�qv��QCB\��I�q��f����w������.h��0���߳�7�m�f|�����Z��\\_H�{���o3nڐ	PN�:���m�f|���_�.s�=�hέ��{���m��3�\k��$T=���#5rk��> _{�:��y�s;��yA�s�c>�ƭ����ϟ �}�s��"�۳ �t��L�������}�gظն�s�ٽ�z�a�o�[m�����m�8*�:��ͷ��y��[m�����>��g��նܬ̯�m���^�|�9@7J1�"(k��C��Xsm�cDt�V׫-ؼ���4����wu������0]
�� {���> _��j�ffq�c�\�B��f{�s�s33�I����B[,H�pf$����Y�X#�p�?&ٳ�f~�0�!�����@v�<� 2�<�����$�Ǽ���H���� (T�� #�C�����ﱽ�o������s�7�wOzI>���Ck�*�Z��c��7�m�1�b�V�W�&s�{�ٽ��ϵ� ?��tX\�%Y����ޥīv^ӫm��������L�[o�9�N�}���� >����ʢL�i��[m��9�{��>U=�����������>���o ���ߥ&D��ep��<�x��0�:�-�<E�Pe����
;�������N<ϊ����FY�� ~��� ��sݶ��1q�'������7�m���{�V�1�eK���~��>{�'(Q
����9w33;�ߗ��38����K�wt�����S�.��;;��}s�ө$���b�c	h{���������|AN�usE#�����SS ��> �P3E'�TM�W��)!�X�����Ġf�0�kypd�1�Gy*��2�BP��
Q��׾�w��n�o��{ݶ�L}�g]�#`5���Ozt�ܿ�{�����﵉�m���sݷ��y@G^��D ���n�ox��s>| ���cm�\�K��3+�m���V�o���}���&�C��b�v������E��L�,U�H�(��2�[��ph�����ݶ��8��f U0�����}�> _����m��f|�����i���t[m������͂U�9�> _���|�����Eͼ���{��{>՚�����.�� ��O߽��-�\L�6�������> }����'������������> ���t{9w�Y��Ν�t��~{�m��?~|�fzcr�k��߸W	��M���x:h���7���L��@�	���qJ�[b>�)�A�Vfz3d!X��^�ă<

��R`� ȢF*$QRZ�"��_}������l����DU5!@�ɫm���9w�m�q�������w߾_|�y�v�o�\^��Д莪
JR�Y��{m1����h�Z&aa�=�m6N�V�Wޝ/��8�<�e���������-����ٽ�o9�jO+��ͷ�Ͻw�i}��L6�"�
��o �߿~O�=�g9����5m��Ͻw�m��<��t��EC���kwc{�cE3��}밹����2~��\�"��]s�s33�݃1$���ȈM���#"2BjK���f^����ܩ���m�3>_|��qr�w��m�ǭH�PN2E$������3��� �����[o��jM[m����l̴����#���s��~ �ݚo�\t���I�~/��?nc̟m��B$Z����b?��W��Ej�&NG�|*^F�h�cG����Q�uR�M���K`c����;x�z���k7%ͳ�-Uwmg��\5���c�Ԏ��gF�1L�z�|pp�GO9��A�q�X��[q��I��PX2F���X������	׬@�txq��)W>�n:�D��xjˬ),�q��\s�툚���,��b y
M�-`˙��Ak,��1��E�u�#ج��Kj�N�O���2 FC9��\d�q-��Fn&�wn����:��:��ATv
=�35�^v���珞�\�� ͳ�� �����o2e��m��1����Ľ����?S� ?~oQ�g#K^�> }��|���s���̛��ov�ӫm����}��Ī��f֕R�Tԅ�2�m�M����ϱ�b�V��)����ov��{Z�@����`���%�+���=��wt}�oظն�{�ٽ�o9�jM[|�U�{���������84L�A�7���9�{�� E{߿I��o{�z�v�ϳ��ޓ���_�~R &uf��b�w-�tr�h��#,+�-x,-`�ź�)nFm���)�����6�g3���}��| ��Y�����y�7˒Q��֬��?��TDdp$���1���g�'T�����<��8�!K�ѓ!q�sC�q 	#�!�P3���ﱍI;�wF������舅�����%TIJ�US��;^�v�̵g$�(Q	���Vk����T�T�5S4�t݇$��7��`v�Z�>�̛IB�IB}�������'*Tph�E`g������ξ��׼݁�fZ�:!B��?E\\��[k�m�x*������{��7X��8�������
��t���7�c4f��K�_�����?cv��k��(_0�޵`����7T�%:�<���B�ДCfou��zՁ��dޤ���-�-u#t��\�*�f�=�g��-y�Y;N��`+��NP�$!6si�2JC��B��D��T, �UK����`g�kv�y#��S�)m���t�:"9D$����X��l��7a�����n���O��t���I���d�	rQ�oy����`g��<��;����X�RZn���Uf*<͸�M]72�[D�V�+��V퐆���N鵭��2N2)������U��fZ�3��\�(��Ϻlޮ�
���MT�Cn��=��W˒I$�۽j��}�`g����K�BI�wf��*:�%���`v�Z�>Ǚ6t.P�7����#��u�$�{4�F�1�C	uJ�T%���}�`v���{2Յ����n�k�A��p1�<���(�������@v���D{�È��� 0!2a�-�Ive3�����+�������,H$|�c;���N����{J��6DJ���ײ����Ź�����VO�����d�&��m�1k�O��Nz�]q��N�Wl�-��``�q�A�}�$&�̠���T������|��̵`d�1����`g�������US�J��{-_(�\�CgN�;��7`g�-_B��B�͝	ޖ�H�%MU+�{���~���P�D&�{�X�֬��2*��IM*�N�;IB�P�m�7`v�q`g���:!.P��os�7z��*
�m0��[���VD.�K�{��;����<jH~1ll}���b��B)I����eI�l�(c'#��&߇�� �����ӿ�jƉ���$I�_p�l��5���\"���*bm��Yt�4�6�H��)D
�[b�t.s��q�D����n�+v�{6�K���*MBK����'!��m��\�v�N����'��b+'I��t�Ćϝ`8�6�<[h��Ŏ�@!�l�`[�&W��Ĵ��(�-1���`4iP�w=k72�������/K�e�g^	�O�x�6��Yf�\7ki���n8{�y�Z̖'-��	�B��I��|q^˩�UID�<����'َ��?c�#�Q�ޮ,����T�R1��	uJ���c�ItDCgk�n������{-_BIt%	���',�iӢ&jJ�N��{���,�\�$�n���L��U�-���ҩt���i�v�9(��߸�;w�XfeXr�Jm�7`f>c����̲��U{�j���I�wW�v���̬,���do��H�3M���j�3C:�kc�]1��SZ&9%���<+<����o�wr��1+.֥F�g��������7`fea��BK��֬CO߹"d�8�N9%���eU�b���!�<�eC�dx ��KI%��S�K�}�)	�O���{ ��(x$$b�����L�x�ǌ�3"�οM�(B�1;R�K)DtDW�����:ՀffU�B��7z����*�X���[���,��՝	rQ���`v����N]9*:�%T�K�á%Д>�wwU��~��;�I>��Ł�w>�J����0��V��V(�В������=�j��'>X�KT�jiH8�����<b�mۈ��y���B�fn��5]6h~����*t;�R��㎪O��VmU������̵ЗB��`wwU�.���ҩt�����vfV�":6v�Z���2~�K�J\�6f�uF�N���US�����`��cO1R�c�<zw�f���t��w��ןD
�igs��X���!�tBO�a��y�x_��8�����:>gk�����O���4]��uW�|e�Um��l�|��;��9醱X���>_b�n�uo��W�m������AN�Muk�tH���|丯�8�!����yw�3۞�
d>�_4L��v�TT�/�8Z���0�
�|��]��Wj��_��j���ߞ�JukR}�wNθӘ�LF��7m���s�ֳ+��z��B�q	/R ������Q!!q�h��E���NV���	pQD��	�-�+.L6�(0� Ѩ��	�Ɣғ�4�M��ω�|�m�eS�È��b�j���^b����ݺv�&f�����lXD/���Y�fn�	,�RIjK�%�%@)�()݁Ő�.��cy����g�d�>�oD�2o��wr`�Q�(H]���8�o��K��v�w��|;������ �7�f��!ǃ34a[����4P*��������+�a I�©��&�>�ͷ�|s]W\r"�R�p�|�wy�����o;�nւ��hB���W�{��&���W�����:�wp����w��^�'����F?��lߤ���V��Dh_��&�I&�!�����P2������]��dA�p6�(V@����a��?4R<6���3���:�!B�rkj`0�`x�4?N(�>Ҕ�O�"H�?/8��g����lц��D���dP���d��0��IÉjqX��"a�+�_��O�!�a�O�����Npx����'�ڟ�Hi�����6�<T��Sa��GW q�\	�#���.ƚo�����q�x�>3�'+�J�������+lkB��(�H�}�w޺�3vi`y�3��'T�F�9�(䡾��;�vfV�w7+ �f��Dʉ8�N9%���eU��swoO��ݵ`���ƺ�2�P��</i�m��Kk�2��3����x�f鳬\�b{�o���ڬ��^�/������̵`��п.���c�n���뒦�i��*��]{2���aݽVc�n���a|����͞�}5J��M:L&���ooU��?cvtD%�7��Ł��j���)�q�N�����â(}��݁��Ł��Z�_�dm�Ry*� ��W֯�bkPg��$!��InO�B{8!.k;������G,�������K���S'��cB"� ��!!"��=�}���A���9t���i�v�Յ��.�۽��{z���7`r�[�0J�ħT�2�lXj�q	ʘ�<h�mf��9::�n,�(Q}��3M5r:�*���{��C��>~������,����ji������`�e_rM�9�.���?{2���a�ͭ䉕qH�N����l�����I(���Z��&��X>�둩��Lj���K��It'����;{�X��V�VoK�7�z��Q4ʩ�Jje�`g�-X�B{���9�.��z��<��S�������ʇ�q���}�ĎM���[��Aܟ������.�χP���A �J;�0x|	 �8J_2���ڹ�Y���d� �:�5�ْ���l�#��dfZ���0˴Q`��G6�˝�r.G7��ٍ.� �V����+i�H��,l��Ԃ�t�	f�v�[���e���Cnٍ,�v�C:�0�
Q:�Z$�L*��H�9���d	s�(�1%��Y�!�3Vb�ؓ<�L�1��6y�.u#u� Uel!	b�)�,���k��j@�HP�	��
t�����j�V:j��ui�Zi�3��f<JLˌ�J�I�DrR(M��Lx9d�H��**$_�7��X��u`~�V��K��֬w�9d�N�3SN�U���d��Q��rQTe�q`v�Z�{�W�#�$�.�Co��r��%LӦ�wW}�g$�BM���`o=�v�+&�e:�d�UUUE����+ �ͫ����:DC�~��`kF�п8�H�n�V�{%��\Y�6W�wvi`g}������(����o��s#�G�:y֚�6�/3=���A��X��n��I)/����,.�^��S�?fV}���!|��ޫ'�����T�5E)�v��¿"0A�>���@8��b�$$�:�][tM׆_�Bk�c1�7Ї��q�P�%�)*`Dʙ�S	/�]�VٛV��糧޽�o����xr�0`f�iٽj�=�eY˒����;��Ł�������-0�i�yo�{������7��;����[	=�o��3�6叚uT��M9��1��9t(���>�zՀ}�eX۳0[ڙNflK̢֭�qL�m2Q�n�F��؁�s�mu������&n��8$��t��{z��3�e� ����]�a����7��SM2��ܧUN��>�Z�Q�!6��`w=��ٕ����(Y�Rr��#��wK2��Vb���5�K�B�#$��֋�`��c 
HF�uΟ8/�LR��2L�@��@ƚ�VYHZ����w{����~�V�{��2C�)*��Ԕ��kv۵���{-XrK�&�w����g655U)�QQ-�v�����Q�%ٽ��wz���n�脡{Bf����DPP���a]Llu*���\�v�9�D���"8_d�/�A����iL�>{zՀ{�ʰ=��(K�K��,k�T�RuD��ʗT���U��ٺ���=�\X�e��С��\ۖ>i�TI4��UX����eag%�7��j�7w���	m����%LӦ�9$�B~��Ł���X��1�|�6�1>��,��ғ,o3�:�F�BR�*k�|i��z�ϲ����M�J��61�UUQ`{=������|���Ձ�d����y�%IU%�S�`�ó�M�1Va 1Xd�f��Oȶs����Z���qUR#���E�fl�=�̧`~̬:�����V���T��"iU)��=���\�6{���7��X��舎I�Ӻ�ljj�S��[����V��j�����`n������*��:��i��XrK�'�����=�݇.P߻��oQ�楍U1��T��`���I%�7o����uq`{=��	V��'"�@���Z�W@�я�`Iń�?V&n�ف>�?~��T5�IƎ"c�8�$�B�>���8�[���u�4K�0��װ��3��b0!{jC]4 *l��2����1�<J�GC��۶�C�C��.
&�ږ��+�ɜހv��K�2q�$��<�qz��<{R9xF|uZۇ�d����U�#!�:X[�JL��5�
�S��-��g�`Ѵڹs��n���t�h����M�s�-�v��0�Z�Ԅ�h15�N��O%�-�JKd$�G�J&��Wd!8L������&��U����9kKCF�i�Sm�;i�TI4��Uh�}���+����K�_07w����'�ӂJ��M��+�l�޵`��`{�1��ItCf�WPRlT�6�:���,��V�{*�Q�.IUV���;�����,b�pZIH�7��B��ݫ1�`}�XXt(�����V���"	:� �%��Vd��(�Igw�>{zՀ{3*����R�����n`�q�-s��f���6c��8�R������w���ڐT��.��������Z�fetGD/�f��v����L�(��C������Z����o��K��"�\ʨPϩE"�%[��
IIe��!`~����>�v�+�脛=�A̩cULc�.�X�uXy�S��Ir���u�{zՀ{�q���N��I�M��P�;�v�u���a�%�{��`{�mԆ��%N�X��V󙹿/�3we��Vd���w���aE�n�
v-���-��`��\��]�,u�l]��RU�7����kbgS���K�7��X�2���)�tG�7��X՛ K]U(���&�+ �fU�P�fs�`owZ�3=���Ca���)*�T��U�����fe�Q{�
c��q X�?��:x�����`�I'�+5 J��[.bI�ZL	�7@5�[ގ H�Ě�i���{��� �f��=YL�9#UL�L���5q�w~V�� ���пI1	G$���N����%1�B&��R�33-X�t$�w��=ϺU��fZ�?qR�g�oT����&������n3��v���54X%�V��
�� ݩTR��"�$�xw?K��v�̵˒_0��`l�OKR�S���iӧU`~ǙN�".M���Vwu� ��ʾ��&�wi-��"�8$�i�;ݽj��̵f��3ٵ`}�v�����YI�6�)�US�a��B}��+ �ޫ�<�vy��*3�6B�|�We�/��	+��G@��B(S��a��}���E\@��h����1f�R��8�����w���=VB��p9��o���x��F��%2Ȭ�{*��I{����{���33-Yo��O��_�c�[,���5���7y��q<>�[��ib�d��!�7�����m �Bn� n��=Ϻ���=XX���.����`����j�T��)Hܕ`}��^�ٻ�j�3ٲ��++*�6f��� J*��q7P�7smX��:&�ϟ;ݵŁ����T��UEI"���{6X��ڰ>�L,6:v����О���S�Q$ӧN����;�$�ݿ����Vｕ`�Бwp������j�x��YL�]�A|�x���|7��^�Z�D���}�?ӟ�Ah�'b$��ϼ�gj�t@���v*�6��}ٽ��of�'���e����>+7N&X��Ή=�ץD�>�_@�� �(�ﳍ:��	S)Za�`ƴ͜	7�n���r�l���y�'�[���0����Z9���~|��˸��(g�����ȏ��7 ~{�
T���,�$�o]�Q歨�8���e�l�Hc&��>w�?�{��|�R�l޳�]�Y�"N��
}
�pLse�Ѓ#5��I�<�-l�G=��t�L���#���A�_Wz-���?�{� �P�����O��z�8�9mg�.����� �|����#��;vA0mڌh��g�¡N{��,?�Vl-ٟv�v�~#f��a)���O��
d�Hݒ{����pf\�,6�||��Sp�A��1-I�`�k�6b .�>p��F]Ú�c��0�^zb�V
�|,ywK�f:vp��Rg�W�������mg�T�M)�4��`�:AoI��݋Ak��J�G_�U~4v����;Ĵ� 2�E!P��!�/��'"�6"̺s|��x�����Xm��ծ�шD�"b�\pb2��f���K!��T�ׄ<���B"�P���4i1�hŵ��#x�B�b���"i�����^ �L�D�C�}��(�<V$s�O�T���p>$t�|~���.�=W���q�G���L�L�0��_�@�=�}W�@dK�$;�O��mxs<�����mU[j��)V5J����j4\�	W�m9����f����n9��b��U�6)�Lku�m�kK�45`ĺ��*��綒�����א�*s�lP�6������lv��6R)h �wwF7gc#\\1�����r�:v��v۶�9A�:[��9 g��V���`eVs�on�ɐ��s�%��s�Nbxp�(�ڴ�ҝ��;�"򂭆��i�����]0�&R�b���++Asa,z�t�VwY�ge�m�[Ab��.��L�t �%,�m�v�Z��m'`Ϟޟcq���˹qU(m��Ռ��h�=���T�b��[�����<� ���c^4���	�3��H�:0Лk�fx�����'Fw3�0�+���O[���c��iu�"��M�N�k,j�,rF�l-�
9xQ�1�S�3s�8R�"�n�����Nv�7�=��=�q�l:9.�P�H�U��Z;���-[J�����
L)��n���TХ����
��`ۨ��q+WXm��4Kq㦭(�e��r���Py�:1�v�(��Kq�݋iF�Бv{8�)�v==/q�����6��;���=�X�:���y���C�&�0Xv�:���p�z�B^ŗ��l�utаՀW�;L�!���S��q����[�)9�����ud���",�I�-��x�V'�s��F��n�+���p]�8��/a�3�hq4+k�33t���\��͸�l��Cq'ܓ�O.�1�lQ=�����xǆz�[&�y���>����*���`��u�ӌ�c6ff܄z�7$sn�q����lK��L
�X9�u����m��;��N� Y�l�hL� %G���0`Ӯ���C��v�9TؽP��ίe�!���n�mE�¯���u�	sq�qvE���x�A�m���X�Ż�i�x�ţt+�ܑ�cŬ6�&��l3Mr�n�#b��Xirhۅ���7I�ֶ)�i�om����r��,�廃3�f0̷9�qru�]���1�n8>����۳���N��ٖ/&�:O�_���:@�~ �����|��h�Ɂ�8h��:��O�	��eL�Cy����NA8#�h��������G���(@"�s�_�
���8������$C�f���A������O�"��s�����^�,B@�	M+�2�>�|�(~2@����6�ڤt|(Ȅ�x���m�r�GM1�2SM��+�Ri�a.%r�2�� ��f���hL�f ̷�]�3X�Z�%��l�m%v5lv��K��sV<Y�vk�b�u�eU�����zx��[FŰY�7�(��\��<O��Ru�7"D���]fIj�ʌ�Jꚥ�m���Md�_s������ٺv��5��������y�)n:�D�ڠ�@��LhMm�0����,)x��%�>K|.��M��a��U1)�D��ͱ!�.e�&�,,ƨ�5Ui���R�2:��n����{-X�쟸���=ڰ=��������N���=�{�a��V��s�?{2��D.M��6%>u(r�t�7z���1��GC~��Vn�� �y��H�*@�U�B��s��ou�=�a˓y��`����j�T���H�Ӱ?{2Ձк;w�_ f�U���;�B��,�NJ�$�];v)�3i.290�-�K1v������j̇fV��+wvR�D�芇�@���Հw��`}��+��;���̓z�QJJ(� �E`��_q~c1�Q���8!A�#�l�>H��4@����n�5,wu�JHR���@��X�ܿ�{�jI���V{�j���g���m�R��J�%�ݧ�V�̵`g�����K�$��SnI�E:pIDԺv�C�!?�w���͵`��Xe<ʰ;��"��R�R�$V{�j������;��j��ٖ�\�nh��E
�: 6�9e�W
��;�e�<�������F�=]���;�N4R�JCaCu���`}��*��ٖ�����6Հy����ʨ���x�ި�>��]�RB�����Mı,K��w:M�����^�������R»;Ο/B�*X�w�٤�Kı9�wf�q,}�٧�L�a+�&�1@%��[�x�OM&�<�I��i{��[�m7V�3���޶kl|��� �IYB0@�Ȟ�y��:Mı,K!}��N�~!I
HRB�m��P�rڦ&s��Mı,���N���i7ı,K�w��n%�bX����8�n%�`xFb'���Mı,K��R_�R��"��H��㉜L�g��e�}ı,<��{8�~�bX�'���i7ı,Nw�٤�Kı<����{4��*=���۲��Q��m�I�<�t�P7�����RY�F��JA�.�[	s���9�~�bX�'�Ͻ�i7ı,O�w�4��bX�';���yI�&"X�%�;��7ı,Jw�ؘ�ǲf�f�8�q��Kı?}���n�"b%��{�4��bX�%�;��7ı,O��{�i7����'{��_L��Vy���^��^���߆�q,KĿ}��I��> a����s�gMı,K�{�4��bX�%>�%)0v��Kdŷ4��bY���s�Γq,K������&�X�%�����&�X�{��:�H߉�.��K���}o��y��(�IKG)��3��B�X�|2�(Ĵ�4� �*G݉�k�&�X�B��3��И�R	uW����K�Ͻ�i7ı,?
G���O�,K���Mı,K��{�&�X�%��^���m��3&1�j��n��]���V�K�u��ɤ�ڏm6c7:�rp�1X�b�B�XW.���z�z9�{f�q,K��yݚMı,K��w: ��1ı9���Ɠq,az���|��WAዙ�O��zX�'{���n%�bX����n%�bX�w=�q��Kı?s�٤�K�&qw6�eB�RQDQ��|q1,K��w:Mı,K���4��c����w�٤�Kı=��f�s�z�zk��~�(�l�t�ĳ�9�{�Ɠq,K�����&�X�%���4��bX���ޫ���$)!I
Wl�⥔"jK�g8�n%�bX�����n%�bXy ���~4��X�%�y��:Mı,K���4��bX�$y>�4v�,n	u�b��W�0	��6F�`,�BFI��m�%���.�������xq�"m��>,�P 8J8r�$_��I�\�CYe�XO�q�.��h�bD�ʗF�&-�Ĩ�ͮ�U�"��l<�P������:�ܕ�n<�s)�f�;�U������Ȭ���0����czi35��S�)��v�@A{v�V�7r�\"���M���\]	+lD�@�X�rZ<��+ �Uہ4#ra����q��Hl�̴kAΦ4�l�2��<���Ћb�H�PDg��8y�w��J�0,jJJ��R�q�R�#�B��(�t�1X�N�cS���;��c�B۷�َ,�jn��⽲@�z��v%�bX��=�&�X�%�~�;�&�X�%��s��?D�K���~W�
HRB��ɬ���D���3��Kı/�s��n%�bX�w=�q��Kı?}���n%�bX��;�&�y�g	��%�m�=.fI��d�%�s��Kı9���Ɠq,K���{�I��4X�'y��5��ͫ�@�/�yd�4؛��m�+��D����I��%�b{�����bX�%��w:Mı,1��u;���$)!I�ֹ���rTEc&�q,K��y��7ı,< G罝'�%�bs����&�X�%�����&�X�%���㻞13��13+���)u���kL�ģ�E��0�L�v�Ɠ46uJ�Gk�k��O��^��T�罝&�X�%��s��Mı,K�ݚ�,K�﷤�K΅��_�����KG8WΟ/B�&qnMګ��[W�m��ZX҅�������Ȥ�xq�ǞȂ!"=��$�O���K�n�߶���6���!m�?@.h�t)�c��5�RD%aR5�c�Z��ț�bc|��I��%�b}�{f�q,KĿ}��I��1S,J{�����=3����g�4��bX�'9�l�n%�bX��;�I��%�b_��s��Kı;���Ɠq,K��3��Q��r骪�p���'D$$�]��+Mı,K��t��bX�'y���n%�`x���{ߍ&�X�%�yӸ�!O\ܒ�1.1�I��%�b_��s��Kİ���׽�i?D�,K���i7ı,N��٤�KĲG��g����R�:�ۚr&��؊:8��by�kRF�Ks�q�i=<5�-���qF9�d��9��D�,K���?�Ɠq,K����f�q,K��yݚMı,K��t��bX�%��÷�����2��8Ɠq,K����f�p� 1�LD�=��f�q,KĽ�}�&�X�%��g��4���T�K�ϧ�R]�ֽY��t�z�z������n%�bX��s��n%�5�^o��3f�f7���I;���%��d��#L�R���eϰ�]X`��~
�(EcIV��`3�?g>�1��Kı9�wf���^��^������@Y����e����K���D�y�gI��%�b{����&�X�%�����&�X��b'��~4��bX�'q:_[�\��P�����нн??�m�O��x�,<�~�}��~�bX�'��l�n%�bX��s��n%�bX�w�� K��4�
s*ئ`����T�m�k=���dƹy�ᨳ��ʮX�<kbe���%�bX�{�٤�Kı;��f�q,Kļ��΃�?D�K��3�n�~!I
HRB����@��9t�9�Mı,K��vi7q,K�w��n%�bX��}�cI��%�b~�5٤�O���%�N��=qsm�b[��Mı,K���t��bX�'~�{�i7��D�O��zi7ı,O{�٤�Kı/ܶ��fd��H*K���g8�ž��W����X�'��]�Mı,K��vi7�LJ���1Do�@�A�V�{��Ѓ ��x�f��� O����+I���db���Fm�����$�,����J
0Z�j�B���i���u��I��%�b_v���.��Ι�go:|�н������n%�bXx���~4��X�%�{��:Mı,K�g��4��bYн=�'�g��)3���3m�T�1�3���[�i�lʐE;����s��F�RI�K2����~�bX�'��l�n%�bX��s��n%�bX��=�1��D�K���צ�q,K�翼��[���Z�<���/B�/KϹ��7
G1��3�cMı,K�w^�Mı,K��vi7ȓ5�^���_i�X�9�_:|�bX�'��{�n%�bX���vi7��1=�{f�q,KĽ�}�t�z�z�?~6����ޢ��Mı,�>�w��Kı=�{f�q,Kļ��Γq,K�LH]�����B������1��r�L�8�s��&�X�%����4��bX�8�;��?D�,K?@�5�cO�,K���צ�q,K����\�������8�͘�I��J%�#�a��{�d$�4[�}-�I$�B�����)⚈�-Ƣ!j��Vy�tv.EL�#2�荻�i��v��mun�-��^��ȋ.�S�k��OD�� ��˙��C2��(�L���s\���RVh�Ƽ�0���l���7:�mq�����{&{�]]����-RV� �&���9 m�����p]=	g��Fc٭u�C"KW0ց�p#�w�DO�
�R��h�Rw@��t���ρ��5v�׳4�Q�K<WM�I���z�@�`2��b�ȶs���K��ř�I�n2y;ı,K���7ı,N����n%�bX���vh<O�1ı=�{f�q,K��so����MfR����нн??��i7
��LD�>�u��Kı=�{f�q,Kļ��Γq,K�����itV�;W�;y���^�����k�I��%�bw���&�X�a���{��:Mı,K�Ͻ�i7΅�^�����-�z��:|�ŞR"{���I��%�b^�Γq,K����q�&�X��&"}����O��z�z~�������eG94��bX�%���t��bX������'�%�b}���I��%�bs���&�X�%�����c��s��� #l�h��lX|:���	K�X�SF�3���D��&،������z�x�;���Ɠq,K���k�I��%�bs����	�&"X�%�;��7^��^����l{]��A˼���bX�'��]�M�����N�`�7�������)I)R�A��7�A�g��~���.����d^�b1)�J�V�B��A���OD�7Ϸ�I��%�bw�q��Kı9����nt/B�/O��kw�,0�g*�Ο"X�%����4��bX�'q�wMı�$1;�{��n%�bX��u��Kı/��HS�f�&-�ɤ�K�"@�Og��4��bX�'q�{Mı,K��4��bX d-����B�����S����UR�s�1ns�&�X�%��w�Ɠq,K�����M'�%�b{���&�X�%��w�Ɠq,K����%Ƕ�.���%t��f5�`Bv�̚��m��������q��]%e6�͒�O�,K��=�Mı,K��vi7ı,N��4��b%�b{�w�
HRB�uq=SR�neT�i7ı,N��٤�<1�LD�=����n%�bX�ǻ�i7ı,M���p��!�&B�o_:�Rt��2I��&�q,K��;�cI��%��-�ͫ���g�'�*�>�n�-[afOֈW7����i�Y���~h�AD��ɑ!U�<(�/s�3/lV}�H�o>q"z�_�!�x���y5�F�ٸH���W2�f��ɏ����y���kc>�d@Onw�v�<S�Ɍ{A����'F!H������/��6uV�)��ՠN7��������e�Ӫժ����9X�k+c��d�wu��HV�h�YY�6��7.6�ex�-�(d���@$�)a���I\�H?}l�@/h�I ��|�`H4R`�W��@���B	��tpD\ ��e��u��l��ϳ��R�1j�\Z���6`�>+���	����(B�@6o��Av�6	c��t1��
�<*�P!x��x2�Y$���:q���#u�� 9����&ya�Q�>#�Gé�PC`%޳�Iߥ*G�Ͼ��
꿟zf��H�|b�gZ��S>�I$c�������(~��g��X�!"3;���BFd������$��8x� ��һ[eA  �)���?��O<� =��jiσ f���u����@P0fP���m�%&�?ϗ�0���*�C�pA�q�`�̪`]' 8�����$D�ˈ@�C����D��!�8�� ?m?G�L��������?�4���8&h����rE�D$\��,' 4��x} f܂����
�8�G�u7Î�44��jM���t��9Pp�8��6�/�]U�6�6��9�5�NC!̈�t.��WA�Wop&X<@�D�T�X�B��Hj4�������4��bX�';���n%�bX��KN�f�#)�MӸ_�RB��HI���{Mı,K���i7ı,N��٤�K��3=����n%�bX����6��7�������/B�/N�٤�Kİ�G��O�,K��;�cI��%�bw�q��K�/O{�O^��=l0��jX�i3cWCX!l�\kb����ۋ�vw	�jc�n��r����q�g6��X�%��w�4��bX�'q��Mı,K��;���F�1,K=��i7ı,K����a=1R�<���/B�/O��{�&��H�&"X��=�i7ı,Ow�٤�Kı;�wf�q<���н?~��K�q.�:|�Щb{����Kı;��f�q,|�D�Ow�٤�Kı=�w��n!z�z߯���"�5z��t�zX�yE����}��n%�bX��}�I��%�bw�q��K��$a?F�x��[�������־\^]]�|^G�ph��X� �+A�*(T������q��Kķ���~?;��Ǯ�Y�O��z�S��vi7ı,N��4��bX�'q�{�&�X�%���4��bX�t�����
�)��F Ĳ��C1�[�ͥ�mw�Fj�u�n=I%j��p�'\ܷ&I3���~�bX�'���Mı,K��{�&�X�%���4g蘉bX�ｳI��%�b^�Z{ز�9Ht�uN�~!I
HRBכ��~	D�K��i7ı,Ow�٤�Kı;���n'�1S,K=���cok�z�&w�>^��^����Mı,K��vi7��C1��}�&�X�%��{�Ɠq,K�?߾�M�~�%�s<���/B�1���Mı,K��}�&�X�%��w�Ɠq,K��D���Ɠs�z�z[�R�zb��5ٞt�ı,N��4��bX�>Ͻ�i?D�,K���i7ı,N��٤�Kı>z��[&
c�Ʃ�;��n��Ml�cI^l��Ų]���s����v�(��f&���䛬�6����N�l�q��W���L�2Yq�]�C�8rkXH`��QҀ��.mC���Ъ�m+q��,y��s��xB��W
���$�A�t��k�)�kT��wQ(x^w�����t!��8jg��v�U�86�@��C��H9�n�k��>��û8��t�g���h[狃7e�b燖���8�`M�D��+ H2.(�>X�%�3f,3����h+��, hQ�un�S�b8�`ՒV#I��R��;Y��,K��>�q��Kı;��f�q,K��{ݚ�,K���:|�н�����h[�gƓq,K��{ݚMı,K��vi7ı,N��4��bX�&��w��(Na2��z�<�-�Ԅ���&�q,K����Mı,K��{�&�X����ǻ�i7ı,O{�٤�Kı9���s�d�Lb��%�ri7ĳ���Og��4��bX�'���Mı,K��vi7İ<�=����Kı/y�i�&%f���˼���/B�/O��;�&�X�%��#�{ߍ'�%�b{���&�X�%��w�Ɠq,Kޞ��=�-�_��is[LGgD[bb@y \�h���j���%�`c���mA�cfg�e͹��6��X�%��{�4��bX�'{���n%�bX��{�h<$�,K��}�&�X�%����b����m�y���^��^��}��y�y\��J�dԴ'����&�Q�𢼟���ɪ�^�Ig�(��
�3�c����Sd�Q�V�(���"�~�Ȗ'����&�X�%��}��I��%�bw���&�=�鎚�/C��k�'�*L�&�X�%��{�Ɠq,K��;��I��>R������I��%�b{���_�8���.�n����J�IE[��I��%�@ b'���Mı,K���i7ı,N��٤�K���Og��4��bX�%秽.	L�0��0e��q��Kı;��f�q,K��yݚMı,K��;�&�X�%��w�Ɠq,K���ܾ�E���@ݵ�C:θ�{v3�u���{u�\�8HY����0�l��ϝ?D�,K��i7ı,N��4��bX�'q�w�,K��<���/B�/O�{�j�[��Zg&�q,K��;��I�y�s1,Oc��4��bX�'��l�n%�bX��;�I��U�LD�/{ۋ�)�E&P:���p���$)!s��p�X�%���4��c|d�����ٌ���[�@�|R򐽳�ap ||H�32i�48�`�?�fL�?1��$�7��]gzZ2�\#���B@-h��*%�9�?o�٤�Kı=����n%�bX��O���voQ���н��MS��Mı,K���i7ı,N��4��bXI��Ͻ�i7ĳ�z}������nVPʢ�:|�Љbw���&�X�%��>ϻ�i?D�,K�ｍ&�X�%���4��HRB�%��)S?SA.�R*RM����]n���Mb�����l�������inQ��!�g����^��^�������q,K��;��I��%�bw������b%�b{���&�X�%���o�����]���:|�н��y��7ı,N��٤�Kı;��f�q,K��;��I��%�c��O��"��2�/�>^��^�N��٤�Kı;��f�q,|C1���t��bX�%����7ıRB�5Z'JI�3@��:W�
HRt!=�{��Kı/}�gI��%�b^��Γq,K��~����ՐW�аU���|A+�"�?�a.D�Y�*`�U���iP���'��~4��bX�'���1�$(��	R+���g8�ś���}ı,<�}�{��~�bX�'}�l�n%�bX��{�I��%�b^t�?��myF�hι����{v�`�sf�q>�(�&�d[,٣E �F�į6�>t�Kı;����n%�bX��;�I��%�bw����~���%��w���нн	��݋���7���i7ı,Nw�٤�=D�K���i7ı,N��ޓq,K��;޻���(�I�!b�$�9&e���j	 ����BH$��>�SP���=����&�X�%��w�4��b���.јM�Jq�F�܊��8��x"w���&��c���b{����Kı;��f�q,K�LD���Ɠq,K��=%�&�I����%�s��Kı/{��I��%�a�}�~4��X�%��{�4��bX�';��I��%�bo�e�O��}i� `Ɖ�����9�e7��٬�����s]Z,��D*��.�F��Г��LoQvT;�[��v-A��cA�;�Lὗkx���$��ѭ��ԕLK��@ոr׋��.��h�ĢƖb�@�T	Ke�S9�35.�KA��e\CC{8K���%W�֯\�t�.�R���`nDϵI���ݴt����3�н���v�^�۝D<X<vm��p �rvY���vi�M��vL���7�g\d�9� �xN����7��{��(�Ɖ�l�D�A��Ao��E����icqI�����6j��!Fɭ��\N��PN�'�kg��CI�Iq��9ı,N��٤�Kı;��f�q,Kļ�;���&"X�%����7ı,O��R_L�q�s$�1���n%�bX��{�I�y#���b^��Γq,KĽ���&�X�%���4���T�K�w۸���L�U���y���^��^��z����bX�%�{��7���1;��f�q,K���Mı,K�&Һ�܎�|���/B���d׌w��t��bX�'}�l�n%�bX��{�I��%�������Γq,K^�炙�_L7�������^����yݚMı,K1��Ɠ�Kı/}�gI��%�b^w�Γq,B�/O{����(R{���i	���˜��7r��VɎh��E��]#Pcmui�yɃj��@UE�:�B�/B�����t�ı,K���n%�bX���s���?D�K���Mı,K��'��Ag�>^��^��}��|_{���D@�����|H�u��1 b����y�3��~��6T��ZF���@똞�b_߽�:Mı,K��vi7ı,Nw�٤�O*b%��zOb�ے\����q��7ı,K�{��n%�bX��;�I��>�
b&"w���&�X�%�{��:Mı,K��^ۂS���q�\g:Mı,K��vi7ı,Nw�٤�Kı/;��I��%�b^w�Γq,K��κ/fC8Ź�L�ri7ı,Nw�٤�Kı/;��I��%�b^w�Γq,K��yݚMı,K����saB녮��6�qt�M�i����:�jF�0W5Ӽ�Ih��O��J.,�~{�D�,K���t��bX�%�{��7ı,Nw�٠�+?D�K���Mı,K����6�.C&3s�c9�n%�bX���s��<�q,N��٤�Kı;�{f�q,K��76��%a2��ry�r�:G�˛�c9Γq,K���Mı,K��vi7�m�q�\�G9��w:��BB0C�� �5��}�9SBǈR�����MN+�	�"�5��)ݩ����B�b��@��O��K�~�t��bX�%�9��7ı,O�r���ߥ��r�:|�о�%�D��Ɠq,KĽ�}�&�X�%�y�{�&�X��"w���I��%�/Oߟ����,F�g�>^��T�/;��I��%�a��;�{:O�,K���Mı,K��4��gB�/OzI����M��Վ4ևZToG	i�ܸ���-��{@�P�t���A�W�O��^��^������Kı9��f�q,K��������b%�b^��Γq,Kļ�o�JL��y��|���/B�/O��~�4����"b%��w�4��bX�%���7ı,Kϻ��7�&*b0�>��C����镞t�z�zX��}�I��%�b^w�Γq,}D�K�{��n%�bX����I��%�L��f�R$�I
$"#��|q3��1���&�X�%�{�{:Mı,K��vi7İ3�g7��j��Q��������
�6e!�BB_	L� D�R�vz]��M��Z��7�%5�a��X��XV��X�5^�';��4��gB�/C�����Ҍ��쯝>^�Kļ�;�&�X�%��#�{ߍ'�%�b}�{f�q,Kļ�{�&�X�%�����ظ���71m�.�CU�A��5��N:�֣��.B�LT��u2��c�cm�J�Q+���/B�/N��٤�Kı?w�٤�Kı/;��A�~���%�{��:Mı,Kz~�|�zە�6W,��н�����f�q,Kļ�{�&�X�%�y�w:Mı,K��vi7�*bt/O������,�g3Ο/B�"X������Kı/9��I��>Hb&"w���&�X�%����Mķ�z��������(�m��Љg�"c�ﳤ�Kı;�{f�q,K����f�q,K�1��_�RB���ۼ�h����R�9�n%�bX��{�I��%�a�c���Ɠ�Kı/}�gI��%�b^s�Γq,K����<��޷��c�]�?W��.�ݹ���\�G���0�����=��;38s��e������}zϑ�0��lX5�oЁh2.�2ez(6���Ȟ\6��"w�^�}��u�|��!ⷠ��DSϟ�>~xC���5_��O�|}Q�t�݄j?G@�$�ɏw����֙�=u��o�?���l�P��O�n�Q�\�?�)�0PN ��R�K��/zD�-�Y~[����y;{��p|���Ĝ�#��BLt:F�L������eԗ��|�'GqM�s���Fc���@X�A��ER��;��;�h�&
���,M«����=���܅	X
�EP����P4hLI|���un�|��d��FKw�2c��:��/�#%��PuYVh$/��=���4na o��r�k� >>+zR]��bZ�A��(�O��h\�H�υ�O�X�c�&�KQ���o?x��k^�J�l-b>¤�1���{��w����D0/���0O���w&��/K�GB{�H�������?���~��7�p!������(E��w�h�l-x�\�@KՆB~�����~�8������w6���_��7s�1 b� ���O�����rm�w�,@YS���u������S��M����[*��*�R�*�UUUUUU$�s�q��̺��OZ�.�[t"j;Z��K/���/����[��˖�q�4wm���;hy`�J�r�I%��:����n��Z�n���+�(��.�Bz^�}m��{/0�����f;�q�O\���:=�b���[�Va�S��������1�F}n"^H��O4��ӆwE7F1q�$<0u��Gj�$��R}lp�= �s�S�-���s���(�J�Q��P��@�����^y|O)�f2lmЛb�s�bmZ���Ҹ�5u��Q���x�X6����`cm�Sd����*�q	 �Y&LJM�����g�v×�0�鮲<nol���!Zkta�찶"R:Ёk[�^ ����l�܎���T�ԩ�=��h���������1� q׳�n�)��N*=���u�`B嫅�s�8���x&���"�I���ؔ9�k�o-mr�서��Ӻ���@`:��:Kn7;F�]�9x��qang]������n���1�C[ pm%������n�n�t�7!/[gu	�kq2:v�b���.]+c�#�LBB�iv�e:�Ѷ�;/+�ܺ9�x�\�s����6��*�\d;�Wi�yr�aޮ1�{��5�W��>�2G^u����`}g��ʹ�l�ׄɹv�Zm S�l[��`�j��k��)qFP4u�O6�����7&p��h�ڱ���ܻ<�X�F�hmM���n�ob<pt=6�m��e��k�&�t{c3�{��lizPM`	L%��nw�+-)�x%�sףsb�88xGc��͍������8�n����]�9;$���7
<ݧ��ց��bW:v�j|iɫ��KicspyH��;�Bޮt*��\����a�:��[����&��c�=rkבE�.�8Bm��ؤ��3���{��v�MJ��{�Aʐ��`��]�	y�=t�.@�v޷2���.{��v��9���4�@�Y�����eK,�Θ,�L��|S_���0%T����/�|������������~���pۧ�2<h����o��	!��?~8��E$X�ʧ8� �?+h�i���hb!�9�?�g�c��^U�p��O���C�vp~&�|�h�E8���&U�pW~S c�	�� |��BE$I���s�DC(pu$ �\�^�����r�����P��� �Ї�dg�tn�o��/�.�)��8h�Y����a5��M�`1�c��ƶ��Xj�e�4u�G���Y#X����g��׈��O:Om;�Bu�
iˣ���0J=<�1�w,����D�[]Ye�9܀@�m����8�L�}�� �M��jT�֣������l ��z�-�gTP��\WTxmc
ms��ƚW�L�^� u�1rKI�I1e�3�4�R+jh5
�J�P�rgY��6��ȝq�'0�X0(]0o3�Z�-q��vz'ux�M�&�Q�\ёp6ۦV{���^�������&�X�%�y��:Mı,K��t��bX�';���n%�c��߿��*�+Zł+<���/B��y��:Mı,K��t��bX�';���n%�bX���٤�O#��^��~��ن�iFFdvWΟ/B��b_w�Γq,K��{ݚMı�1=�{f�q,KĽ���&��z�����i�[�s�|���bY�"w���I��%�b{���'��S,K���t��bX����w��~!I
HRB��i�}@���[�s���n%�bX���٤�Kİ��}�gI�%�bX��ﳤ�Kı9��f�q,K���`^[�q�PA���+��S%�+Q��s8Ԙ��x����Iz���ܴ�;n�3�qK1��ı,K�{��n%�bX���s��Kı9��f�ʄ�,K���i7ı,Osږ{38�%�q.m̗9Γq,KĽ�;�&�Fn[/�
UB�����uD�)ÎXR�z���<�K��p
���{Z��,�b���i�i4Ĩ�b0�ƀ(U
�󸟢X��l�n%�bX�s�٤�Kı?c��4��bX�%��v`�)�B�� I%�|q3��L��f����ı,N����n%�����c��4��bX�%�{��7ı,Nr�w-�UT� 4�\/�)!IЄ�����Kı/}�gI��%�b^�Γq,K�$�N���i7ı,g�߽�5��)�Vy���^��T��{�&�X�%���w�Γ�Kı;�{f�q,K�����&�X�!z{���}-6��(ac0kuc��r=���+L�s�]&cF$fѤ��D�Z:�inC&3s�g9�~�bX�%�{��7ı,Nw�٤�Kı;�{�I��%�b^w�Γq,KĽ���.1���,��q�g:Mı,K��vi7(G1��=�Mı,K���t��bX�%�;��7�*b%��{|�zۜ�M��t�z�z����Mı,K��t��c�N[�J�s~��i�f�!F)�0
J!�h�B񘛉}Ϸ�&�X�%��s�4��bX�'���	���,����O��z�$�k����&�X�%�}�{:Mı,K��vi7İ<LD�{�Ɠq,Kޞ�}���L� �+�O��z��{�{�&�X�%������I�%�bX��}�I��%�b^w�Γq-�^����~��{��W��[�-�' �t�,F8�v���䪚�Xܢ��j�m�����/B�/O�����n%�bX��;�I��%�o;���|����KڍfیR����RE`g���RI&�{�V�ݖfe���$���.�䄑����V�ݫ �̖o�ݵ`n�ڰ�c��!�@��RU�����7wmX���=���:�&lѐJZa��v�N��M /1���S�=�F������J R�U�j�R�x	���I'w�a6G�EG�X���In���^�ՀffK����}��X�4�N繊nPNέX�:�Ի@qK�;h�M�H�f۩�T���j����`���!G����򧊩�Z�Lb$�r+fU�l7we���j��̵z��پ�O\r�C�C��rK �ݖ�2՛�s����V��,��Ll�BG rKٙj��̵`��a�����`{Q��q8�T|*�+32Ձ��n��wvX��V���N%A5�0]nK�bD��l��$��Iv��A�M��8p0�ܙlJ
P؏ T/�Gƭ/�m��sɺ67\U(� ��x3���5�ً�m�b�i����ď/�.������-E�]��М�l�p��7��y�E���ڵ�#��3Ur��a�<z�;���8�8}p �=C���8��%��6�bT�#CV�j�ۙ��5��(S�j,c��*�ylZz����vᙣ Wj�v��N�7��/=�F��d�tq{GTذ,��t'j% ���Hj��R��P�foV[��9�Z�t>2ڋ��mq����&�\�O��x�ON�6� ���L�a\����������̖�2Ձ��j�3�f@c�s�!%9%�f{%�l�ݵ`f�ڰ<�1��P�C=�Z�ŭ�I4�U`f�ڰ=��Vl$��%���v��V;�i��"m7r
I��)'�ٕ`�d����w~V�����Z�Lb$t�V�fU����͟��j��{-X�f�=N�ԩAMUJa��i���a�����v�7
u�k�1-m�F�<�b�qR���J��nl�;���g�֮|�nՀ{3i�*JQ@
�,��}�A4B�*������wR�ަ�|@��$���|��+��K���75�*p�Z
E�؊U �`)@ �����ÿgmX��V��K�ٚ�z��RGƩT�X��V��*�I6g�e��ݵ`{���TRGQ�'H�7�n� �nՁ�fZ؏�LD)���V�b�C�@�9*U�{����fZ�;��V��*�Թ��Yz1TAP��؎\݄) Cƹ�.��#�J<�ܢ�u���zىi�+�x���s_����w�w=��?fV�|��n�����6�uU�8�Vs�j��qq�nՀw7e��̵z���*�-j�10�ӑX�v��fK)7Ϻ�G�ī�%�M���!#�-P!�\-�1� �(qD�h�R�D(��@
TJ"��w{ѩf�=X�X�8�%UF�%J���&������ڰ;�e�\y^ݫ �f���P�TP
u%���Z�5.{3~_�۵`{2X��2�rW �ԣ	օ�7��.3۶bT�6D�$7eԎ��)cY@TN8�B	�UR+��Z�<��V��&�s���V���E$u"qԊ���e^-���n�ۛj��}�qq��y��1��*2�V�ݖs�j��I�fm��j�=�5�Me"F�ʅT�s�j��-X}̫%d��oJHV!�>�T��Մ�߷x�y懝����(�&��U\�Z��U�E�F�[
,@9�9��RO����2�uR"�8�H��2Ձ�,�n����`w=���`�n�1�����fQԘmZ��h���7\l飠[=�ϖٺ����͋g��ϖ���������-t(��!�nڰ7��tTd�UF�G`��X{�j��ٖ�������M�y��2�$�����fڰ>�e��W��}�|y�vD��T�XjI�7~Vr�]�{��a��\}�ߕ���n�N��:��8�����v������Vٙj����� ��K�lw@7j(���M �?���pm��{[�m��F5�KH:�,�X0�����su�9�Fzٜ�v��!'q�e��זи���-��tݫ[s��G���Gd�:�j��8�]�u9M2�&65$��rs��JMn�rjM���b��tɠ�7Uy`6ۤ�{k�A��ܔ!(�!	��ؙu��p�x�m��B[��Z����(Mf�J�3�t^��=nj{�҄6rh���͹2b�8�	&Iq���T�b@P��� � B���x��x����)�/7[���0��ܑ�ayus��]t���X�	�MY�؄ң��͖}�`gs-~��=ݫ ��-6�kSr:t檬{2��"d�L�`u�eX{�/R�gs#�Lڍ��ԦT���nڰ:�2��&���`fnڰ=��:lX�Jba%T��5s�绮�73j��fZ��Q�����n�J�FJ��n�X{�,fe�;�j�=����Ŵ�ݍʍ�j�ş/�G;r�:L�7,-T6
�!`��v���s/	)S��W
��J($���j���-X�2Xw�,�dUN�
R�"�3��WZ���	�ta
r�˓e��H�2�AƵ�n����c!�nIi�����%�CX�GW.&��_�� �P(H�Z� R�C�M,���u`��X��V}�2��QGFH�$����ʰ�X��Vw�j�3��C��Td)�%Xjos6X����e��I�n�X��ܭb�nGN��U��̵`lG8��w���v�=��ķM�w̜J�CV�L\�Zv�D���ru�$�&t�l�Q�n�9��f��W~�ݵ`��`�d�=���w��L5R�IU*+ �fK �{%��̵`gs-^�l׹��GQ��$����͖�2Ֆ��:�������"�d�{ZQh��}~o�	}u=��7�g��EC��B�{�3��g�U�}���Άf!�壕��k���{˯y:ʐ�k�p�6�����R�Aӄ�q��~��Q{��D���� �ބ� ��s��&
��S=nfo��BN=P�=����=���D?��u���e�մ���b�Fv0�Y����0a�}�C�$ 6�����ܨJ�7$E6�m���y�����\��;��'�1��ɠ?��3�ff���&�4?Yb�O2�e����O����S<�Ӛ
I�&�\ˋ���b5�$�a�l�B���)¹9HA����u�x����a�F�����jkoXk�L߰Ci�@bY�H..|u�[�e�@Su@��*%��a�H�_8j��Kʿ���W��Kr�D�B��5�����h	DA'~�a^�`��dO(�\P`�9�~��qկL �!�(�s��&�S�SKGo� Y �� ��gc�>�< 1f��0�E�����?-�P2
�1�x+��Mؿ%|t
?�9�@ 8Ǆ�����H�Z �"�(�O����U����%`���P1D~�#)8�<_��v?�"� !�~'�L�~^^.�X��[�p��?i@PC�Ƌ��ƃOrC�p�|"pq ���P��j��|O�K��ז�3�,�{)��J���Ia�����X��V�̖���ٲ��l����8�:������nڰ5$�V�������fZ����o��b�0��m�B��ц:�uڲ�(�áͱp�8z�Z_#M�n�m��B�g3$L�"�<�2�=��2֯�o�mX�7H�r2���8� �{%��̵`gٖ�Nf;Ԕ�o��6�k���ӧU`f�ڰ3��Vj�S8�v�s6X{�ӦeA�R�S�"�Ը��w�`c�ڰ��X����Ff�él����9[m)H�[��P*ꮑ8��Ԏ%/�N�i���Гh�� BU/� ��\k�ɺ��XY���Ѯ6aH�����>4�4��(T�RR)�PjV�V(P���k[5$��[0X�#Cd�NE`y�2�=�s2Ձ�̵`y�x��i�'J蜍ێB��m=nzZ��v.�گoFX��rXk�GB&�*2�TET��73e��̵`gs-X~̫�=��H�JQ@	$�;����K�l�nڰ1��X{2^�q&��^�$E
5I����j���eY�%����`{wmX�YO
��Өʃ%H�5q�n�X�l�=���g�Հ}�<tT���!N9*�=��`jI,�ߗ�f�ڰ<�2�
N�o�	JJ��45"��i4/0�qA0i��=�	���i� �3�g?�̎BF$5�i4B&g��џ!���`ߗSZ�f�W�v$�����Inu�����\O^� �pga�vb�)��X)	S�J��f�p�my��9����GNw u�N���,8�c4aE���`���Y�6������
u�Ii��-�e�T� 3K�����[�طP�^�;l�\=[@��˷2��&�!��b͡���m؃۫KiC/cVv���ki[<��@QR�A��jP���Pр�+F)B�� �nt���ҟ2�i\h��X�(	qwZ#�cw*@
��4�Q�m��N�V{]$����TgM����j��{-X��|�􁛛Vs#�Lڃ���r�9���Z��M��v�76X��W�l�1�T٭�F��r+�Հ{=��I&�wmX���y�iʄ��J��R�6S9��`f�ڰ=��V8�u�y��LD�T�9:���fZ�5%��ߗ�c�ڰw2X��n��mf���Y�J0�t���1��g��ŘJ�u�,�`46�GV�n35�4�-�߾��Xy�V��M\�K����x��R���q5��)'��|��{|��!���#��1�	�{D�u���L�H\gZ����CSW"c��.81$V)��DkZ+	!gB��K��`w=��y��û���ETn��8� �n�ٙj����ڰ2wu�����)�lt麒�RI�e�`{smX��V���{vX̕N�m)U��*�P�;��V�m{v� �n�=酁�K����j���DԖ��%�cQ���q�pl���<��4p��v��N4m��DR���5�v��̖{���=�����iʄ�����!ԫ �s%��l�ɥ��͵`c�e^��癮��I)NDS�,̚X��Ր[�ķ�
^A2�&/Wd���JL9LrD�������%l��nT�e1�J�#����P
�D��;�����>��;�ʧePS��D)�!a��8���+ �n� �ْ�W8�2��=�=n)29U"��d�5q>���̚X��Ձ��:UWMg�O+'�6O
Ӝ2p����s�������:ȶ��:��>�d�3ޘX��֥�/���`��[ntr�6�N����؅'�6Հo�j�?{2�TP��e6���M���*�P�;���;�,�.&��l�72i`}�=�cp��TV��n� �f�=酇�ܡ�˦�C��X�	�rR���IGA�A�-60�#8��R��8�S���ր�[�I�!&M8�&X��P�$ D� -*�H#߷=�`c�%H�����:��&�ٛ,̚X{2Հgs%��q{�kS���⎋8��+N$��2��7(��V�P`�7(��󀮩��W��4�>��Հgs&����,nk�c��QAS�B����V�̖�����za`}�oՍ�Q�(qʩ�gs%������s��̚X��Vޡ�yJ�n�G)�,5>�fՁ�������V3�ݫ ��s-���R����IV{�RK����}�)'wΒ_�>�4K�#���J,�xQ� G�H��&M�`i��M��Vaj������SUaم�Y��<�,%u �nW#���=�:3<!�=�l
;�xȁ��%Iis�z��I!�uۜ&��,M2(hg%u�.�	n`d��r5�8�����$<�$%�.I�E7"�����&��4���%����[5హ�Pwd�j��Z�2���5V8[Z[�ی�ے�H��K{Rѵ��d�g���c,���:H�u�����0�k������-�fX��'UkM�L��Ʒ�NRM�h�4h\���*�Ur��۹j�3����粬���#�m�1��9�gs%���eX�L,w�j�����H�����:���粬��~�K���m� �n��=��H$RJ����=酁��-Xw2Xj��nmX�6�:������`jI�g�u�mX�L,�;�m���Kɛ�ú�GM��y6 ݅:M��l<h��� �0Z"��.�enD�|�ݖ�=�`g�0�s�����V�!�{H�:!�$�>y���+�S���Q2�x���Ai��d�K!��9B	�$���'|	��	��O�?8�@��G��L;#G	��# �h�VR�
�b�C{�gY�ԓ��4�>̫�
&CW�̶ރ6�MS�V�M,w�j���7۲���ڰ?{��nq�e�RM6S��a)�f�V�ݖ�=�`g�0�>�0�M�1��9�gs%���ͯ��ɥ����)'��g��)��H!p��t���v��;&��`3%KT�V����Z�@a�(u%���eX�L,w�k嫜]�7v�{�)�E$�
*nJ�=�E1���Z���`|��Vs�Qcbr�1)�,}�`�ʱ��[����n [LI3�&=�;~���a��|� H7Iې��Z��L����"���b�1������A�B,)
y,�t����I9�%��ӂ0�eD�H�57�ݖ^�Ձ����^{7�`���8:!�$�>y�=酁��-Xw2Xź�]�i�#�ӻ<�`�����uΩ�Y�nMmvL<�ֳԘݤ˘�������i`{�e� ϳ*��9�v�z�m�6GR�c�D�X���8�M��vX{�V{��q6w��QM��N1�9�o�e���eY��{�4�3ٶ�[;��{	R��i�ET�.>��Ձ��K��Z�|�P��q���H��P��;�������R�Q�H�������M�]ֳ`u�R)���QSrU�������o����>y�W9���o�I=�ر���^ks��z�ez��v�� �m!&mF}X6ˉ#'9��)T~����j�3���>�d��0�ɥ��Sc�QH��nT��3���s��w6X�4�>����l=�3S�ptB89NI`��`g�0�y�7�͵`��`]x�SȊ$�eJ�T���2��=���;�,7���7e���UUOj��AJ�T,��j�I6��I�g���`g�0�<�8K�}�yw��rZ F�,�3B[-��Y�"�e��qH���;� p��H؈B�j���Cl��b_}3�����W���hh�'�����v��obU�}���V]^#��[������|��;�}��[����X	�hi�Ϸ�aޘD�	(f}���&o�I�}�ŗ�8���]�ܯ�[�����(I��h�K��Aߠ�|�'	��qi4�fΰ�BY瑭Gy��(�	�|�$ao;��ř6�) �&%ʐ�$pԵ(	W�L���e�l�o��5%K~|I�O'B�&c����j���i��p(*��Ā. M�����:��T�+��Ϡ%��&�S��FjÙA��ك��7s}F=���B�׶����m��1-�����<��A$B|�%>~���+��^{�{�4
#O�	9����������`S+������o��ۙȄ�H4W�o63F!�����m�F;t��:n�mlhHh�B@�Xc�%�H�rj, 訰����|� ��(li���|��@QJ)6�����c#�h��M&���k	���ٶ��!# a�{D�B��>P�J���ph��"�<[�n,�t<z��ts9����獉�x��]E���M�G�����k'�F0��G���I"��a�`:k����o�$�RJ�A�I%�<�J�UUUUUUAM��h��+�NwY�J�3յ	a������q�u�����Oi(�fV�e�sc�nx���Gx̡�\��gj�;/$q�����Խ���a�\u��%���.͵����=�v�ݗ\��2���4M�ųU��#fH�\����]S��Gr�a�;8�m����u�� �)vŵ.G8bp2��WS�N�kn���=� ͬ���s������.�1΁�J��De��g.�	�tҸ�t�8#�|ĝ��:�i6�($#Ю��
74Kd�%�X�Z�ƌA�#],^��,.pai�����%fta��� �j�'��	W� X+��kd��ZԵ܂��7[�U��s#���n��6���	6�$в�օ�E��j���������4���R-�6�!MI2��l�j-2�S�P�^����<�h�n(�[�۱A���!q]�e� �[���t�y0Ӷᵋ!����s��	�۞]TE�Ց��v6$(: �ԥ�2��{&�vd�S/d�� x��%z��cxς�"���g�ɞ�o
nz�l�,���u/7E�U\�Qg�����N5�r�Ɏk�C�,,&����1�bP�[Y�`����.���36[A&�G6�q�ewvL6��}�[6�%�a�z�0\��km�z�3uN���6 ��m�h�ok����iU���)�r��)l�4I�� ���l����c%�<�M:�c.#t\/��GG����<��j���qv*�-5�� �mu�`�UG=N��r���7�Şm70!([|�0�9�h�ݞ�\��9p�ֲ�����tYe[�UC�l[T���
�;��K�t�G��j쀇X��8��L�m&@�F�(5�Sf��ˉ��eP&�v#���I�<e���Տ7J����	�3��e��n�S�]��Y�k-�T
 �Sl�*��e�-�u���m����7P,�$ttK���%��3ͬ��V,y��-B�MT����C��P�E"��2qM�ʝ�x�۴L���ؒH�F@�$��B���1��0�S���?БD��`�(d8��S�c �ȟ����������~�4�����>3�W�01v�N:8\8�_� .���v0	�"q�`tN)�xq7����~W�~0(aO��??�~	�j���/4�p
�ҙ����t,�`h4~��33�����mL�^�\�9f!�La�h�A��M:��g��`�vK�C�v��Vo�K9��	uѶ8ec�= �y^���>^w��]n;y�u҂��n[���2�>;f���`U����Z�Q�3G@���$��hC�n�f^,:��c��=�)���wn��i�t���U�nUZ��z�9�F.�nC�16�EEΨil����W�s�
S�*�*UX��؈A��y�)d�\Ź�!���U9��x��R���pf��P���������%!�ԕNE����>�d�3ޘN[��j��W���Iʎ4䢪K �ْ�q�s&��6Հgs%�9��癲�H$����RX�4�;�e�7�l�n� �n���(�Щ�T!UHXo~�ߕ�o�e�}��a��e�`{��y��RGN�E`��`{2X�L,��j��Ğ����+�Mb8.�����c"紼��	.�v��%Esm�״Q��b6�0h��S�|�ݖ{���Z��|��n� ���=��J�T�UI`g�0��߂�:B�(%��P 0|P���J�H�1�:{w��ٙ,�fK������UUOj���
�D�X��V�̖��%�����������r(���Ȭ5.&�۲�;����zaa��I'���X��:�Tiʒ�$��K �ْ��za`w��V�̖����t��xL�s�۱`ö�+1՚�j���E��c	���zZ쒚�����p� �̚X{�j�3��y���,{V�d�9t�CeUQ`~����IG�
l77�`��`g�0�\M��Cz�9�Qӄ��X�vX��.��u�l�d�\�c1L�D�$�1�K�I��\�~�8�?~�y4d®(�P�b`�G��#���饁��j�;ѷ���2F�9%���ٲ��ɥ��{-Xk{��`��:��SRU2�JrK=酁�qs����}�,��Kx�M�~����Ńs9�x�r�շF�n�N��1�べ�)���*�N�W������j�3���>��oI|�s&��PP��q�NE`��{��ù�,̏]�����Wl�x�aQ�T�h���,=�,���`}��V��K����H$���*Ia��Os-�;���;�����0����0��(��΂��2�$�$0��	j��� A�D�Eq��`F$Z�0���Q�B�?����u$���jV'.��6S���?g�Ձ��ͯ���`g�;y�n�ԎQR�ų��E�U��Z�����i�&�i���dQJ�@�ԥ*�_ o�e�{��`g�=_0��ڰ���Z�
U#r���=�d��I�s#�`wsmXw�/x�^��6��eJ���G����-Xw�,7��se���UUM�8��
�D���$�ٿ+ �f� �=��S��z�n"P�z��DL�ӑXw�,���π����Oo}E$��?+��Q�e�)
-��q�����v��Yۂ.f-��߿-�?�eCaM��%F��|�<�%5,+*X���%�4vS�qL��p4Q�fKa���z�'0�חt&�[<i'Lś�u�3���ƽu��l��pQy��5�Nz�t��X�E�2�a��\i��f,��n�� ��reƇL�W[�R��oa�z�ZBpm�-LV��#ڹ�)4[\�=M���rs�>Ě���+.u���%��Je����y�;�4#SV� U�e�
����~I����X{�^�s���AѲ�n�D��f�6b��'!s\ܙ}�cR�$��M �����{��3��r\���͖�ele �IJ �*I`g�;�پɥ�o�e�g}�����G��h�Ъ�P��9Q�`}�Xw�,�.�UY������tT�Y
�*RUJU*�a�&�ٲ�7ٲ��z<vĸ��/K �z�A��FHܧ$��X��ne����/O�7ٲ��}�%��a�cJ����b�\:j�X� *4�јx�Q��=��*�v�K��)�,���`g}0��jI|��f������Ң$�T�%8��M[^f|hݤ��K;nt�+	Q��X�E��s㠑�O�	6����z^/�����G$ZT���jF��}';��RI���3ޏ�g�1mF�B&H��,}�,;�o{��}�K��&VBF�!M9(���R�o}�,̏]�����x�{��`nVV�R	$� "
�X�G���%�����l��X�^F)�|�&ԩ��̢J\:�j�4���)4A���m��AЪ����9Q�`g}0��Xw�7�|�s#�`w�D5$�J�T,;엩q��f�s#�`g}0��l3�oY�t5Q�7)�,}�,���g�_�5?��\�B,jϮ]bI	6B�Բ+V��C�,$���Y7 ��$d�j�I�JBB�
8&H��ہ̆�EH6``��b�H��A �7�q���l��=��`�uUEdM�*�R�9%��qq�e�v�&���JI?o})';�m����q���g}0�7�O}�> �f�=����)����l�6{b���j�+���-�0�+s���:��Pu�5;Eg��v�5c:u�7ٲ�3����z<z�_0�ɥ��V�l�F�"(r2�K ��K�6ndz�̚Xw�/W7++c)�I��U%����3ޘXw�,;�,�0�c�UIM	�r���x��^��͖�̖�.5)��ɲ�h�Z���p`ٓ��3?g�P�+`�%*�-�O����(op�R!£�T���}��`o8��͟���=��V�q/����1�	�r(`��
��yS��.9�ukٍ�����W��4�YtJkG��Tp�'������;�쵩%Ϙ��`��UObmIT�rRX���z�3smXw6X��/RI���QT5�"WʢS���͵`g�Y�I6f��3#�`}�DT��Q��#�"������3se��z<v����X�jel�����Ԗ��K��x�g�Հ}��`b�_��M+3i�"
��i��d��m�&#�
A&\�Z�,q��z�4�H��\���w.���h2s�t[�"Q���R��wO�y1�$�(b�u�Sg6Ѻ0��E�V�����u�M�=�ͪz���R�'d�'b�[5ɮ.7F}��NHkh$M���d8��]k�R<(��56F.��]go<��wT�7��gڻ-��4Yh�κXk,�K�9�'`�HbZ�$�;��J��oȱ9�Lh�V).�uC��;xz�\�ƀ:�nB�ڶҽv�L�	%I��rL�}���`g���{��RN�|�a�� �MGT���j�s���w6Xnl�=�G���|Sov�ȇ
�5R�V�͖��K7�q�fJ�g�o76Հg��mP����I,5q$�nl�=�+]���a�o=��=�C��Dڒ���*��;�J�`f{-X����YH>����]3�B��� ŕ�1��2�n���s��N�I�mf��)��4pi檏�32(~鹿{ޭ���+��b"�*�
�PIU*+ �=��j��G� S�g�>����xG�
�տ:>�s_ ~�x�Aw�R�lM�P
!��Lo!\h��2f�.4�)���R"��Q�@�M�N�|Τ���ֻ32��8�g}Z�[#�����Ԗ��,�ұټoۻj�;�����)��IRD"&J��y���u����ڰ��,57��,{6���UQƚn�T���e�x�}���f�;�J�{�6?f[m�T��P�<��7:�C6��s"˚l̺���qQP
Ħ�T@tTq�*E�w6X��,�ұ����6Հg���P����I,�̖���zV;��`�d�l3qJ��ڒ�:$��,nJ�d������K���k{ŉ>^ȷ>�u {��+�Q�>"������2}���1������_��9��'1}9\��ɀb��¾�8�P�� �W��*V��/� �6peʍڼOߴ�Pû�o��:џ��e��6��Yی|�n��׆ρ�w�3��J��o���#�N4i0�J� i�&�dZr�w�����$xT��v���?�oW&��u�M�K�5(�.�_�=�����������_��z�B��"���:}�Whߎߗ�e�]���ŗ��i�W�_jď�> {����o\, ј
���y�نSK*l��<��G���AW�(�_�a��hH���`�Z<5x8p��n5�<��d}52�9�-ӈ$$')�ҕ.X��R	!�L��� � ��Wh*p��O9ȟ��( L�`$0/��o|��O�'F
�݃H��'ݓ�;
~LE��/L���h\��u��#�[}��ﺗܠZ��E��a�M�T�^WF���Q<k��Ow�v
�;�z���g�� �2�0�Ϸ�7�5X����0T �0����˵�����a��"<�.�����j�t���}�'loj�s# e���_3��ߑ'�.�ˏ~Km}r݁�����Q�mXϰ`�R��_w���Vw�q ��<K9���t=�g���Xo�d�T��@"�S:{�~'E*-M��L1�0gf4S��N�����Y#�m/���Mm���������ޖq
�.g0+�޾��Oo����#�A���$a���T�q  �I�䖬��K�}5��*=�dmLY����=�r<^����ŕeϐ���x25=}u�9�w��$ A���	��n�p�l�_���Q8������/ �e@�^ ���� �8󌂒M��>x����� �>�!��o�&�~S���NA���4U~◊c'ʸ88��!��P�>"�^|@�6�W���8��;O�j�S��C�J|C������a����!�#~S��x��$ �]'�o�"$���<�������S��bq�pJ�@�@HH�B��O��{����ޕN�k$�JRUGa��s~V�͖��*�TB����́��Rr&�t�RN���=�d�w�,�%c�>�e�������6�����:�l�Y��3JhF��"��1I��F�=/#[&5p�FUI`�X�J�`}��[�s�{6X���A$�"�$�{��ޥ�6wsmX{6X��{�M�T*U �7QԨ���j�=�d�y�6g�e��l�v�)�IN�EG��V�%��ٲ�3ٲ��rV;�u�9(t����:������-M���H}přDqĂ��$0�9�o�Q"BD%jՀ#Ɵk�M^�׊�>�=�T������NI`�X�J�`}��V��%��%��]�i�"GP�&��� F3	����۟m�5���햔�ƞ�"r���UI>��Z���j�>��j\_03ٲ���uC[ ੺������=��R��a�͖�͖{�X�R�g�b��UZT�4U9�w3e�{��f����V�}�j����FH:�B�#���Ը�{��`{�+]���Z�Ը�s6X����A$��2&I%���V;W7ٿ/�;���3��`m�T������ȸZ����cFr��bO�f�A�n�LJ0���U3��I���N��t~�aμC���кnĺ�{��e�q\<%&���àc��y�ǝ�.��{YW^X����.�@�]1�9-�;"�+�Z_:7:.�{�^ź��;�U�r66klm�<�{�̦\���caIt�P/%��Zi��S�K�lLK6Ž��H�7b��Q4ӵ<�س�i�z\�8��:�x�K�a�`:X�]��
��L\ۋJ�3��YdSqh�)D�%�!%�%�i_�9#a,��u�r㩝�`��;��%��y:�m�闢8�ĪnB�R��9*>������{%�g}����������OvJeF:*8�J�X��K�ė5�6�{%k�3��W�I��3kc�NTd#��X��V{�X���q��m� �f� ϸ�_@����9$��*I�{��{%��=�fՁ��TꆶBW)��������-X�}�����V{�y6�Qq�f���Ӛ��,}�FQ�Sn�g7���[���z�n%��(ͮ�c*�U
�	9�3��X�������7ٶ�<�l���N!S��RXw�,�'I��r�/�;B�9�~�A#�i:�w�KG޴IL�7W	��P����T�X������r�����V�����6fV����Dș$�}��3��Vj�I���>K��6X�ڧeP�T�):$�;;�`{�,;��}����Ov8�#(��U*E`{�,;�,�����e�y�G�����E��x9N�+uخ$���S�R�8֮�� [״7a��:�]�D9'���`}�G���{-j\_0;���7q�=��B�蒪��>��z��ٹ�j�;���3���6wkU1��*��ԨJq�����{%�/����鸲�t1����e�n"Zs��@�)(�F֢�GG���v{���r<v�^QU
�
��GNEa��3e�o�e��};K��s7�`y�9�7M�N!S��RXw2X�e���j�>��X������Fu�M\C�`�uظl����'E�ǅ�-��u͹�WQ<��uJ��M�'�|��.��nm� �=�W���`{3j����R!R*J����Z��8�wse�f�����w�\l��c���
��T��wse�{=��M�2V�76ՀxY�"���!$��s�7��,fJ�`{=��0��P�{�Քj�O��~,HB���,�5
�8��R�|q�>"� `n�m��"B"�" ` ��@s��;Τ��}&&Ȫ�C�RX��c�7�7w��w6X�2X�1�\i�!�LAt���vNx�:ݚ5���V��Ic����n�1E���'q��'{﨤��wҐ;�ɩs�̕����U�EJ$�QX�염�l=����n�,�2��I6u��dn�%
��:��=����.j�~��V��,�r��@��T������w�X��V��U��������6�Li�!4T��,�e�y�.<����v��2�`	�*��|i�Z�]_v�R|g��)��Q5K���H��#�7�z<BcLK�m�Q>M&�@Aqv�ǒ۩i�L[bP���q���^�u���sv���lm�F� ��
(�
J��{P�(8��PDn�v���X��<������]��H/%ש�Ʊ�J�%hK�SLj�4�g�i|���4-�5�(ѧ(�Y�#f��qǷG��� zܮ��0��r<�3��!�YBo/P	�nםֻk��m�:���-�쓬�G�T��*�* .����Es0!n�\.�rk^--���ʖ����U3�T�6%@��H�]Z�U������`}�ˣ����V�n�eH��F)9%�י�`wٗ�̵`�d�\�l4�T�)EC�J�V�v�`{ٖ���6f���wj��
~eV(�*n�*�!a��y��+ �͖^fU��f\,��J)��**P	��{=���sջ���ۢ��fZ�5B����z�ԍ���74�K��5i9���W$��lX2M�331��Cue�Q2����}�ym�ٗE��̵�D/�nmX�Ƶ�
�6C��`}�ˢ����a��3;�P�,F��~�'�� ���� (��ӝ�֬���fU�8�l�cڶ�QJ�B�T��,��V��K�3*��.t�YR��F�T��W�͖=ͫ�̸XjK�y��+ �v&�TR��G$�<��V�./f�����V��KW9�04�i�R1Q/g9��[�<��ĳ�בq)H�����i[EHb�s�℃j��:n�)U+�=����`y粷�0ǹ�`wJx�F�%'N�URB��{-^���{�V=ͫ�̸^��;�QMUi!J!H�Ȭ{�V�{*ýɋR��m��:�o[���I���`HHU�ѐ��qu�Gf�������|��'#�}/��dP�Q'�b!�S�u���{�>ۻj��՜�M�d�!T�S�N�T(�ǹ���n���j�Ry[�V�e-�@��L!T���.�R�����;��c�M��#�?y�QJA-���.�ti))���;L��׳ʬ��:!�kKc;g�Z�n|����ԇ�f�ڰ<��V���R��=��|l��(d#U*E`y粯yĸٛY���n�,g����a�n֍Ȩ�Q��G%X����2�`{=��<�U�a�m�YJ:n�'*;K��+vo�X���<�U����i �E,����Kd����|<u @��=�t����� ��px�*�B̃�@7K���k��`�֐&7��i��.(X��� ��~�ʒw�G�	����[�%��j���eX�L,{2�������ldsq��v0$�<GSl�v�6cW���en�8�-=��;�(�B�ӑXy��酛��7n�76Ձ��Jn�%�$u*��raz�l�ݺ,nm��=�z�3
Z��T�B"93v�;��V�{�ﲰ�>���p�tК�t�~�ߕ��sj��raa��I�n�E��1ͧ��2��"�<��V��ϻ���Nw��̓~�F�� @U� ���Ȫ ����@_� ������ 
���� ��Q?�U��W��^� *�Uت ��pW�  *��U��W�  *��TU�� ����d�Mf *r�u�~�Ad����@�����`|��� (  (   x   >        �    t8 ���OoNOM�YԦ����=����S ��t�<��^&.�@�J�� |3S��kgW�[��^���<λ��d�{���kף�}�����I�x ��-�}z=���Ɖ��H��%�������os�Z9��;���WG�$�  �lW�lw3�� �����`� �@��t��������q_M|��>���:0�:=澞� ws�/OMz=�7;{��i�K�-�gҟ{�:}�����u�͹�|=��#os��x)TD	UPɦ�
R� #!�����0�JR�A�`&A���#L��S7��i�U=M &�� �1ت��Q��F�	�CL���`�S�"F��$̓i���4�� �Dh�M44@��??���?���M����
"�@EP�DDS��B
��Z�?�B��M *���QAEP�'����X�(�# ��������N}ў�ϜUQAEQ��*'�}��S(��{Oc��u��2��{�;O�x�����p�� ��������w�U�F�;ջs+qǢ-�Ĝ��`$�*^<I���[g-�j� "�5�3�nwi��ȴ��r�+��� *�D�x�|�7ݭkv=�|��T��U���q1�kɰg]����8H�;̼B�Ŗ�':��ك;������37Ι������lB����J�D���kJ�/Z&i��_;C�v�(ݰ0!�\B^�B�%�)H�[sl�H7�t�Ͷ�H��C����`Bb��E�s����#�۲A�����p��t����noe�1�gm��[��V����dі]#03,n��%�K�ȶLOmoZ�SAch�Z�7ul)�ʖ32��5����5�n볥�hc��oi �ֹ^j�{��pI�b��w`e���$R)���$'74h)�
<]��wg�v��Vi)�_a&>뗹7�o���.�Z�.�FYBDn�;w�6��=/�ΖVf�l�x_*�1�^��%���]���]2j^�;;8�D�:�T�/����0����v���`���Xh�⅔M������u�d,GKa<�0ڄ& ��;���lA��r]��7)c�y���c(,p71a��F�N�|Y���\4��Dh���L�ؙ��y41�`l&mw�5>�[/]�ӧ.��A��6ZV�m�!;
Yr�v"�5���ƈ&&,zV^��8��rQj������7x�,{I������w;�moQ�6H�^X;���sk ��g;62�ׯg	wf��'^����rл���JU��3#U�[����9q�R���v�v��ʙ������kRP�jީ�i�#Ʉf�p�O�&�e����Cl.��A-��7P=�����"t����6f��(�A�yi	��I=�T���;:��݋�V��؋���U�
����nY˗��j��1;��Z��K�	�mh"�s.%vb�z�x4��[�|%��uҗ��XEK7�y� hј�Y �(.$�w+z�_ToP��U����2�v��&�$ s��V���ޣƋke�B�̖�4��e�A.^�O���O�BA
Ɛ�S���ו��k3vfDC5��Wmck۱�P@&�Ejy��p2Ʋ\�l�JT��3�l/WV==���}�Oy�2�k�u�hb[���"��B�3����CAY�`��โ���;�u	�a�5��'fmep6:�vA0���F_f�h�4�������Pe��#��I�ΰ���x;��B�4�e��ʰi&�p,Z��n3y���h�G�����>Z&t NQ'��$��</,L��gx$7�·��n��+&A;7w#�d�ӭg.ju�Ay.�Ҭ��A6��,{�.�Y@�z�;���;3Y6�[�+$�3	:-W�������j�6\�8`f݋�j�(�Ʋ��h\�Mfd���v�9�V��&�c�����s.@aظ{w�[̼7��7o�L��vD�%ig;����ۂ PB��ܼ}���9�0K(mM�xJ�΃]�6��w�׳U�O1Ýh�n]��|#�F'8�Bqc9I�h��m^ۓ}�sw�u�md}qc���Fl� �v���Or�
4��-�u��J��K4g���L#F�'H<a\��0��X~=����w�n{1nr��Y�쨒�y+���k��os�磊�c.�ww/��pl��P|��n��ٗl&rys��7�7t[ &��/{���?x��%�4�sjg����;ҤI�G��Ro�s��5��1����.�w�ns�TU���T���O|� ��w���"���<Ӽ�Ê��icw�-����                                                                         ���                                                                             t                          �lK�b\��θ��sb��6Ɇ�gg�z��Ų2^�6:��1p���v7))$�8s�!�3�X(�Ll������ UԗLD�9�a5�1��<%����U��֭^;W��h� �X��]P�Sr֜Y�3��}�Si���X���|����y�+냎������p8�+�<��ˋ���ǝ�I�ֹ7h�v�㶣f�qg��g9��A�p�	Om��&ܛX�5`�A�!�ۗd��bz��Ӻ� lmӝ9�وrr�S��� �4���r%��)�2��,a3Ŏ}8�(�F�n%��v@����=H@/g�#�6ӥ<:7<�q�g����V��U4��)�	�n��l\;���gT��"紾�Bh�q��<{g��.�n���s�I���թV-qs��u\���pM�{kJ.�dǙ���7T`I#m�`Z���݌Ɠn8��c`@��ăD�*��Ԛg��c�K���l�u�׋<�s�I�Gf��,�����9u���0<:8=��s͙�M1�m[���������8�}<�(�@��>|o�V톞ӳZ���7Zqہ���]O\�R�u�v�0����[s7���,�d"lnRY�:�`�-���u��[:�'�s�tJ{cqnƷ�$����wvx�p�I�nћr��u�O�u��sse�:@���Hcx[�q�!���i�3A�W���7s$!Bn���a�ټr�\-�v��0�lS�����孋n�B�7�s{�j؈"�uUr�;�A�qv!�Y�	Dۓiz �xV��m7ȴ�e���3/Gj��m�Q��Fw�������Tf&�)kU���c��>7~�w��yv1IL9{i�$��^�6\B]m��2Ӻ�'Y�=v�\��Dv���˭���֗��m3Ì4X�v7��N��^��u��{t�7H��n��v�}�����=&[�d���g�-A��n5l���G���셲��`�p6���	g۴u�#U�<Avl�pQ͂��n�F��9��1��4������Tz�B�Zz��ǧ�����[oԦAV�v�H�m��A��k���w�É�ݭ�ѧi�����^ؔ��(��1cq!ǎ.����Ah��0[�ӗR�7f�h����^�m��6.:�n��G�x�Wz|�Ϸm
D���G�:���]��Z���nV�P�3�����׵���,�mQ�.�ݡu۵���n��Yz{S����c��qC�m�My7n�u�Mxnn��z�F�-��s`2���;m�ër��z��i 	Ƭ/U;���oe�y��rd㗭����>|����;����J�u�B�wg���q]��5�Z��=s]UCu�s�V��7e�_���~���~t��V�~0Q������Κ*~�?7�@09˒>�#�?S dK�W�Θ0V�ԛ�l�c����=Fe�gøt&������$L�rf��`gZF�&�l8��]�d������)m���L��2���it�
�a��V��<W&N�j�K7oR4�8=��2�#�Ľ����7�!J+y:�,�Y[)x�ovG���2B��zP��r�R����&�F�v����t��Gp��7	68C����ni2��˨��I
-C���(֎ �F��x
2�7�7L	�N%*v	�ٰ/���ͮ�Ha8�p� �:`hB8v,��o�f@;��w��5d$
���`i�X��n�FdCF�����"�
Sb�[8֓;	��P�3��b�)T��E���d85�D9X����X:Hz��j1�e^���CI08
#9�"@�kL�
3��ӫ��y�d��.Nl(8r���&(�:��7�stt��e��m�tu�+'�hl�6d�'tsv��e(N�6m�\𾉠,9��0��L��CK,!��*��2weޘB�(pżD�9 ��"����$�BN�$�`5T'7�}�7e���\�wl'�#���j�#AJ�e�|!A� �K�P+���@�y����	3�"�c�V�'�o�ǏV�&������젠��m�R=FL��z�n9��i��=!!0o��#+�#�3K�g@'�tS�n�Z��6$	�Bt���t�rj�8��t�b���3�dpN!���(�:-�Pe,!	�7i�ꆲ�h�+��e<�|��)Z�Fj������j�"� �e`���`              ��              m    n�q��sx��d�F�PL����oc��j�"p���9A��;�1nÇ�e�:L��N�h�8IJ��^y���;bڻ&^rgl^���ݵ[�90�F�6�e��Df�"#���b꧒���r��m�f��lmmZ�gS��-���6��7�N��ez�5oJ��n�C���1������5�X������9�8z�ͮݸ^C�]l���.�.�X9�b�ѵ�]�Ѻ秕��ڞ��\�:�t[�H��.W�̽��R�2ęI$�K�H����D @$�ūh�w�(e�CXA�e�5���`�
Q��0���@��e�ʎ�m ���* g"aW��LPt9M�^w�|��  �  %Z�-�d�8�u�5�n�gU�ѭ<��=�k�����^�����y��+gu��gv���ފU{p����+m��yp0�x}�����3�<��P�ݻF���m�ݟX$��+|�q43=Yw�wfx}ݻ$�B�LGi�I�$e�c2G�wt���7�F7߆�(�$"j�{9�x���gqx�9�z�˻/~�bl���/�؉�!�gϝϞ�ߠ7I��n��[�ca�S,-���yS�ۉ��}Yw]�M�'1��`z���Y���jB�	^ΰ����1�e�e���$�n˔����J(�C#��ܽ�Un��D1;��U�l_	���ʪ��3Ap�u�#�c�!�@����m����e�fwڪ��Emy��NI�Y���y�w]Yrԅ�wuY�B��#v�{���c�1�목���u�݃� ܈HrNr7Xl@@�1��߾�I      *p8�q�:��뫠rDc��cC��ثuη]\�&����f�e	+n��Z�3���2[h��R8���{3|������m���/�/��$P>�ݙ~��
�׳.��g6�aKpĨn !!�����@�1�{/����g�����>@*4�;���1��cv��wn�E�7��<w��3anϳ+I*勇ۘi���b0�FBL�Ĥ�����n�g[nbw^eV�+�.Z����E@ 㷽���ݯfV�qn\�]׮��7{ߠ�)��d�KLj�K-d1;����b�M���Y�w;�f�̟fW��7.'���a� "D��@9�vv6�/߾�}���g� �j�q�ɱ�r",�㉅�7s=���c�}���na+���w"��� n����p�����}��;뾼�:�>      Kr�6dLۛx^`Ư[�Z=�n��y���8���լ5��!=l{h�q�7]�!��vY6;\w�w{��'y�M���hɋ�vE������O=#����υ��������{)�"l W�<n��m�r=�U�{w~��I#q����j0��6̒4wr��vi��`���1��ۼ0�T�d,�o@@�2����cD؇��ʪ�陡<	�u�m��H�{�/;w=>��I
0\I)B�pA 1I$��;�/��q0��f]�z�ۇ#v���>�9��F��S懲�4o������'tl��,HH��L8�
�٨S$2:/ۿ��wWpA�=w�%b�]�	7L�9}��k���_��l�b|l\-R��Ac�]XЬ�v#�2�Y½���(sc�f���D��c.[�Ƶ��Ѳ�ӪFٶ��D�M1&h��T�yY���O��4-�m��S�����3QgtWX�YyS�V=� A���캡�g�ڝ�w�ř�^����ʉ�6�8 <ei�h-WfW
9���¦��67�vء�!�+�Ʉ\���3�28L���h7b���pˎ�C �td ށ��
|b�T�P� P�;�!�#G�/s1�oD>�n��̢D��m��I�\Kq1$QÁ�=T.3a�3���Cwg}36'wA���K�n\Nc��I˺��b~�A�������Q���p@�D{*V�'ka99UBت���*2 ����T��o數��I u����Sm��L'�r������L��@&�9���$ o�=��ܨ�� i ����M �g��>��$�ݙ�����p���|	̷��*����G��3* 言�4�͓��w�y���      M�m��ə�&K�w&Ŏ�q�c��D|ѷ������x�6�v�����Ϝ�|�۫t�v�E8�=;�H-���v��wwm���U$΋�L���aP�?7.'�~��������mȞ�#�ݙ�o�ۖ�,�̻�6�9I n�n�d�}�Q��Q����r�3��}��f&�b������9ӟ/(a��� v�>���UI����3�HϩǏ<��b���w�����U�ݟ|0�I��Y��s�H'W�<M���[r'w�O+�2��v���y�\j�������)|�rﾡ�������}��>�z5�*9�gA��$��}v����^�*LJ*�|R@>��޾��`���o��4��3��|{�z�����˿�$�@JpmC��`LE�Ț���~��P�s$p����sF����׌Y^�8�@Gݙ{jZ����[�F�#�"�Г>4�DU���O���>�T���9o�~�M��Ś��Mۭ}$���G�r�v������W�>�q;�(
��G�pC��� �̟�R�+�[�M�N[��\��p}Yw<<����2;�=    UUUT�q��ے=�u�ĕ�ct�n��9�����jY��v��[����+in2�*�~s��I�u{�&�5�c��n�V��~rr,��܅���� ���%�t�"�w2�#�����ݯX ����mʊ �u�$wo�t��Q s�w��U|�m���.�͵���7�昗���������}�]l��e	��"�~��'2��c�Ĝ ne���nB�p�]�fW՗-HY��eހo�m�L�se��ec�M��Ñ�^����j�[r�wH@{��N?�}-Cݯp��&q9�ȡ��Hϫ���Ї`�� @��~&�/��3�ӻ�rI#*6����1�@�LR.�r��P>�}�7s���F��A���Vܵ!g�s.���G� ���Р$�ހJǑm�Q��4e�efu|�m�,L����-�N&�Rץ�}��USQ���G�׻�d��}�wO���k>����~�u���nB���ۿ�R�eG��κì���0�?.���J��		�V���HJ��l���5�|[`u����65ͱ�0��匿������ ��m�8.铘I���Ű��c�n���I�t��@�"R� 2��B�^Y��E�dm��u��:6�M쳗�H4���j_s|;8+��yN/���|�m�        �                         Y��Su�S���z�r���Ρg�.2�m��/�����9�\lO��c��g�cW�/:ҙ�[��8�h���l�3���#�gx�p�UɃ�a �5z6v�㉫�z��b#k�y�ЛrW���w|7��� �Xݞشtf���v׋IZ��۱Ƹ��N�Z�ƯcA��f�z(\�mq�5�a�#�Fܚz�<�X=��nݹ�<=�����0��sz��6����iH6�Zr�nň�^��=�^�.�sQ���^�^t�x�ì�֎0��n���c����й��pL�� ��<�S c!�(d�~&��D�V�?:c� e�Y�����k*�X�ؙ�D�0fŵ5����ɜ��Χ�oS���     �2�.�LY����3vd�<����i�ӡ��9���Ưu��m��]kcN�4ݫ�����Яw�_*�p�����S�sg�������w�P�p�n�����o�ە��9ws�/��w�{�u5�&�;�]�d�u�ۜSU�h�;���ZXK�����u=�ڑ9�Qzy$H!(o���;��.f�ۺ쪖�Y������c��罷Cw��$�7
0aj4�fHJ�l�#G�/�1�������u�ȼk����	߀�� ��9VzrԪ��&�{)���� z����\m�U���L��y�^몖�W�^̻��n����u�ەu�`@�����=DD��e�h�:;�h[���q�}����W�<�݄�m2�,[��i���}ݻ��Z��=X�쑲����uݵ.f�̪�]T�¿;��Q�9�˓�K���$��;�      	6����nl̺���~/c�<Om�ǅ[�<a���d2�+�Ӻm�ݳ�F���d�-�p<ۥ:6�ӧ&:�ٯѕ�ͽV��%K.������ߟ���z1�*3+�USֺZ��\�����:��$]��R�-��y��s��]x�aݗr���bNe�3�7}Z6b�����Gu ȳi#!%0�!5*���<����xL/済�F��N�`�B��,� �z1�*<3�@�!����m���\Ѯ����S$Ư}jwH.ѿv%8!�!���3ܮ�Ps�^i4)�,�غP	����#e��Ux�f!}�6R��+��_Ns�<��n특yQ.ٚ[n2�nZaP>hf#T��	�H�B��b�;=��ܨ��F�dv��b�j'{C��!�<z=��,O2P��� L	�A3,�{�����j��U�U^�l(������҉p��wP>\�1>k�0*�7k�]����Guf7P�F�.����b$�Cz�ۇ$n�^G1㦔P��_<     ����ʼ���6셷Y܀�{���<�F�	��i�a.�۴sez��g�N�o�����𪪍\�Eɨm�͕�s�����{'�@�v��ؾ������B�i/݉N~|��ݣ=�Ul��:Gu?M�2�n��B��w�$�ْDѕ#E�db7�#��)W��{ߕLn����/���_���Ŷ ńHB�2F0!	�}�Dy�Ϩn#���BiÒ3�!�����&�Qᘍ�#]�qغZ���~@w!��g}� cb!.�Ͷ%�,o��S���!���/��H�i?ΑB�n��G�� Jd�xǷ��U���7�IrI,i�$��,�U�E�W��s��X_��m���g�mѠ����H��	h"�-�8���ȑ嶠��B�Waf�l�9�p��B3wW���-�5Cw�]���(E%1	���������ޫnf	�U� k1X*>R��>6M�|��X"pl�� �FP��Dqˆ�\'�3�0<�BX孫��2�.rgL��ɇ8���ٽ�p�r��Dл���&n���YF��D;$�B#�{5˙�����@�!������b�[ʷPۿ��$�Ðb��(�%2!����Z�y
�d��j<.��Z�|v��)p����r���R��4Z�X��`A��h�,��~C��9O�v��(=�> � z��@�9�Sm�"$0ۅ,(�%�KZ|����ln��@i hf!}�\�${�#u�k컖�^�a�n���}BiÐ0GrH�`����-��xn�t��C��@8���m� ��  ˈ�v/�P����nڱ=L��u��ns��Dkx�&�/baz������l[p�9$���NN�}�!�[�n��^4����ߧ��~���o�bX�����F�X�}�� w!>Cw iO��q>���5H{���J����3]߶I$���Q�$��jq0�r���zE���Cu��$w+��X�+}� �"3T�H&�����,_���G��7k`��>���.�+����^���Τf#v���� ���,��\��\T{Γ�� w!>G�d��6�O�b��v� ���r�a#��Lȴg����
�v��Zaxiy�<1v�}bmÒ7P�Eԝ����T�m���&&������?ː]�:=�[�7P��ڔ�l�s�F�ZV���!v�R7�Խ��������2�ؕ��xl�\��i��_#���
�着��t�]�u͠�e���u
�}�w-0�  W��F�\oX�p��(y�[�b<8�'-v���J\6s� �.Ѽ�I܋���ó*�8jSQ-%Y�~�������ZےI$�H    %��^:�[gNy������84'@�ۮUí�������nǴn�9��4V���3�m�8&��nI
MY�C12�9m&àg�v�T��(�b�a�;�/���|3�,�.Ю�r�a#���CH������8A�H�F�w�?�ڪ�q~�a�Ͳf�j��9#u
�;����1i�T%
.�J@�_�]�K���u
�i��a��� t�b E�/�D؀7P�U܅x
>��$�8ٍ(�i��3P�$�(^�W�Vb��l�]�Wr��ۺ�X���`dH DK A�mJ����m���@���G1��)�*<3�r��<#�?:�,�\Q�����Zh���"��bX~ :C1�g�DЀ3�!����=���_�u��D��	?�,U׈4~��!����Gu��R?ٙ��ۉ��ĵe�%4�� �i��`��w*�C�`yt3�#���b�ڕh� j��[�K����.ѧ֕��� u#1�`{��,$��a\�+�B;��:F�4%󬵓CrA$]�DQ��.���s�H��u$"�H�fR;��E�l��5VZA9Dѣ_(�:�0���+'�mI�Lk[�' �f�h�G^�g��n� �C�U�&�u#"�,������J�@���l�t�w��d�R�I�De�:R�Yos.�s="�����ݤ�zc�s�z>��                                   �	�wm�c�-��9I٤�.v�v�K�ڃt�.�k]�=�65Pn����X�������S'c���Nm�N�S�ƹ�[��Z���ڡ[������6���N�7�9��r��\�ے5�-���z�m8�)��m��҅�.3v�'Q���M��z�v}�'b�.F��XNs�W
�+XJ��(�QY��<�v�8��&�����I���ɥ(��(�'
��cb����m�.·��۶��@y��%l�����硻si��L��Ta��Q:I�Q���p��� ��x
��`��}A�D���t���y�`t�{�����me\�5�:�>Ig/#��S��~|      ܖۦf3fd�*ktZ�#&T[EҊy8�=�۱���t��P�9�%��q��W�;\�RϾ�/n� ������-Ej��܃�^��1X��"���]Df�WhWt�0��Di1���5�w-0��h`��7�M����4 E�N��7|ᛩ�+�a�.�����tl�����H0.��_jM���T.<@�#@���5��uiXa���f#v��%4 ٍ��z��@ҟ���|/U^!Y�{���@�R2�P8XM���Z�8�J��+��1��>���y�v�R� ��m�#u
h�فH`�2���f���*�d�iީ83v���I���CI�7P�Fm��jҎ��֙z4!u�������F��Jh@��:Gu� �R�N'�1R�]�\�e�	���!�@"� �A;�i�u���4.Ѫ@�}m���2Xhnl��J�RFb��� �xe8sᘍ���ؓa����cu�m�%a��g�]���E�%6 �5ԝ��	:!f��o��}    �����j�� +mY������=�pl���E�m�ۭ]����t&sB�(��=2Rw<MU^���W;/�غ������}H���B�}��bH��m1>�Q��T�o�̠>��+Q�B�& ��vC6;�p���Cw��$�	E9M��	��q)�܅w!��>��0����p2P�
DT�W
.OA#G���7kܔ؀7P�#���Ӊ��H̓V��C�Ӓ��G1��R:MUv6�n�6ܹ��!p�!f)$P<q�Y�{�$N�rw!^�6ጛ����p$C%�pQ�����
��dd�$l��$
"u嘓a��7�;�x�7�žDu9�<�g�y��:��x�.HɌ�pI�4��Aگ{����6�O�b�h�+�l��#���B�u]��O� W��B�2A|�+����� ��C��jH�C�_��ݜ���{��ɨ��.*f���ۇ13�@`�v���I���Z���6����3�Fb7h��SB �B|�b˯ͩ�b���>$�͑7=�ٹ����'���      ����,-t'���;�a�61��8��\�v��o[���E��m����Z�@���5�/I99o]t"��U���uQq��rEL���!�����&��Qhf#v��	�ԑ��44#u��yØ�
 �'-� ��7jM���A�CuU��wI$� �"0dh�X��ZjH�J&
v�r�7UO|��a�j�f��H��Q�F����:�R'�uR�#��;�c_t��!��F��@�I��q�"|v�n�n�0bT۪G�7��[<6�k]T���B���7���p�#�1�r���U����}�b��((BQ���l�t�^�,�)A.o�x9����$���m-�n����u0�eJ
�$��>���y�р�P���� �=�Gu�B���*@\����u���4��ĊD(+�!"�H��;u����w&�w�g6�z�B�01t����؝����tsF��^�2��<|OPh	��cth+�m^�p����������=�u����ۓ�Ll��5���7�8C.��L�S��E\v��GG+O���}hn�����)�b ���G ��V��nZ��q.ZA�!Q�څ(ܑ0�{ʯx���-8H�. �u�P/�q�"|vyX��sΡM��0,�cu�wP��c��ɵ�O(<�k{7�L\�=�|'>^}�y����c�=l�)3M�X�BSR�0�{ʬ׽�c�W_�ˡ3�]!���� >Ԧ�8;�:Gu�S�M�ᘏ��v�5�-8H�!�*���'x:.^���m��nfe�   %�qo7q�Fz��9ny��ۚ�v��6�.����΋m�$U����S2�Ԏtm���j���,0���EbBDԑ����Yhw�n����F�5܅y�n:m�b<7Q�G`ݡ��)#���A�C1}��O�A�둻��͟$�;��	����mb��$��I�a�y	���Zkݒ&��U�N��pឰL��9��\��o���GuA�B��˖�/�^C1�/j���Ps�n�h y��m�X!.�l�\����i���_Hؤv�1z1HRs D
���b�!��v�����5Z�!$	 �1,��[�N����T�9Uz&!����wQ�5=���O�b>�r�3wͶ��=[Vo6x4�e�I�p{����q"Fb7�{.d/�^C1���si�b`�^Bȍ�ro�Ӈ1��#�(���" �G��܇k�%��:��y�]��od����Ӊ6˂H؈�̄��51�[��ܓ�a��#���  �nR�7Q~V��oP�Ӳ��B���A�C1U��B��5�3�C�ۼ�Ey�	|H�鹿     q�rV� ��gJ&G�l�ͭ�B8�q�n�F�]�-���N�:�l��n|��[���.f��$��뮀�ݱ�QC$Q$,����n���ﾧ]��ۇ1�I�����TDv���gu@��C1}��O�ֆ�f"�R�����n�k:�m����v�̓D�K��}}��ΰ�(�kݼV%S��e	��d� �c�F��B�h�̫�nB��5�d��!�SI�b`Y��H{<2�9���F��v�����m�0��n�g,ܼ�'U�o}}����]��=�j�g�c� z��G1�R�&#�Q�P��g��$'�T&".=�P�;�H�v:�γUx�=�m���*����^�ʞ���I$)��F�I$.$,�#��uƲ��^#��^�剃���Gu�����G�b7H�V�r���w*�]�)�a%0���E,q�{�#u�,>���lhlV��ƞnh�A�[�_@t��7�������GԎA�B�ܖ�$s��.ѭ�d�!x���p�b�6��
�u'u�G�0M���M�������k�����"�K*$W^�	b*w`*L��;_V A��1�Q*���!����#gA�>�y}kFm<�Mg'a��lHгO�yBFj��������t�X����FF��0QZD\�wWB] ˔˶f��l�� b�>ZkuWeo;��{��=l��w=�Y<to��Ǐǉck!4I;�޼������{��z�k��                                 UUU"�۝��`Vy��1�3n�T�؍^����vxR�t[.�sh�n�v�,�q5�n�z���by����U�Ț zw=pq��9m���n�{]��83��x�uLzݠ�w<���p-��8���O=�,��ϓ��n
�,tqr:'y'^�`}0�#�(� ��ld��(����8D��3m�@(�S����W�q���1/<ON϶��]�4�v�/mms�ɲ��I���j����5�� �>Ǌ��qvb62:�z@ի��W���8��w'\Wl���'v����ÎC'r��.CY����4���h0��c�8q�v�N�4�L�Cf��ÛxwI��Ӊ�/���h4{��m2���4�4�0L�Mi��G�ߠ     
�vsfxî�t=&�v�1�\�͞���������W`ts��.�ۃ:hE�Wabۅrrj�������&�Z(9�;}���{���7hn!��g1|`T�3�Ѫ�D��KLn�����4!��n��Gu����.�r�Vk��C7瞒I!
'���PE�Y����|���� ��F��e̅㱃,ى� 3�{��-�w
e�u
�@��ro�Ӈ17d声s�C)��b>����?yǿ~�ݕr,��b�[t8Z����S��n�Of���ު��q� ���oAv=�W��a�G6 ���c`���]rӄ��>����7�{.d/��]H�G1 �[v�m�qt�,g���c�j��o}}���{ԗ�I�BH$��twx��2��H'{v��H��%�$zP�	"w��q*	���10^2$�H��%�$jP�	"{ԗ�Nr�I�9��k���I��+҄�I\��$�{�bH��k��ֱ������On���	9���Ĺ�$D��K�H&wv$�H��%�@�@�B�"�47��I$���8���)`�[������۽�_K� �&�IpI��$�H��%�$���x�J�� �'�IpI��$�H��%�$�����7����YYMA$vP�	"oT� ���ĐI���$�w��U�J�A�
��R\A9��$D��.	 ����I���qX�2��H'{v$�HyB=�& �	=(I�;�K�H$�@��)�j���L�2g$�333&I�M�:      �Z��M��Yᮧ�,ѵ����{G����{�9��ۧ�>=Wn�N�n��=W77�Iɮ���ݩktF9����y�P�Gol�҅(v�$D�.	 ��ؒ	"s>��bK�j	 �����D�).	 ��ؒ	"w���J�L�=W�\Ȓ	"{ԗ�L��IZ��R\A'e	 �'1ߪ�d����r!�bĐI|��$�OJD6ʉ��\A9��׊ĪȒ	"{ԗ�|�kr��Iޤ�$�w�bm��ߧ�����Ue���r+3%�̼�MQ��J�P�G�\A;۰�j	"w���q��J��S"H$��R\5͆m%J$�7��9��X�	"o�K�H$�P�	"o�5�+&SPI�nĐI���$�N�A$Nr���	�l��0^2$���{ԗ�I�BH$��R\A;۱$D៞�8��6�)C�
�h��JN��I�9�K�H$��1�cĆq"��!4�27g|�v��;�K�H&wv$�H��%�$rP�	"o�]암�A;۵�5�7�K�H$��$D�i.	 �����bUdI�;�K�H$ԡ$`:@�q���;֤���/V�}�K�H'}v$�H����b�����v!�В	"st��Oz�I�J���\A;�9*�52$�H��%�$_	o$�H��%�$�Eh=���~I$�8-�Z,6�[�\��>d�̜��l� �'7IpI�Rv%A$N����	���10^2$�H��%�/�B�>� ��&�t$��}=]ė��A=T$�H��%�9
�{�bH$���\A&>���u�$0*'�IpI�.ĐIޤ�$�E@:���� 05�BH$���Uw�VSPI�nĐIw�LA$v0�J���ZP��]�����1��OcKv]h)���m����%�$jP�	"w���H'{v$�H�vs��*��j	 �җ�F��'7IpI��ĐI�����PN��J��S"H$��R\A7��$xE���%�$vP�	"}�j{��)�$����A$N���	=(I�*'{IpI��{��/A$Oz���/���	 �'�IpI�nĐI�"@��ܓ6j�G�K�]      .�pI�2f��㡹UY1��\�0��s�3����nå��\SֻT��=�[r�p��6���UUV�S*=b\�R�hɌI{M�$nP�	"gt��N��I�9�K�H$�ӵ{%̉ �'{Ip�A5˱$D��.	 ����-P�'3ߪ���	�]� �&�Ip�*	=(I�;�K�H'3�=x��YA�
��R\A&�	 �'�IpI�nĐIo��*��j	 ����Iz��$�w�bH$��R\A<���^�-�b3+�,]1��˃6�
�A$Oz���	�]� �'�A�b	 ����I�osؼ\�MA$޻\>�)l=&56Q*L��$�~��$�M�A$Oz��|Ĩ'~��b`�dI�=�K�H$ԡ$D��.	 ��ؒ	"s?N�1%�5��!^�$�H��%�$޻A$N����	1�j�d�Ȓ	"w���|,u�X�	"{�E�
P�(Z8κ��331V�$�fwps$�4-��{�-������I�5�K�H$��$D�).	 �����UdI�;�K�H$ԡ$D�i.	"s�����q���|k-+0u� S�~b�A�`�!�B�* 2B/1�[����6��Ӥ�5�����As�=�ڢ-yg���u��� �k�e���@쓶Q�4U�`��f�4M�Y!w5��PˍLDa�nYM�Y�v~�����%&+�:\*��xI�-�K�=v���K���y׶ �j٦�����B6�D��d1�I�J�Ѥ�d0�6hr�v��d���;.���A�:6�Wii��P�&\�M��Ñs�&"�A�.�{��۷��sF��Cf�'5NwF���c����]#���# ��F�sẍ�9��=���fm�qW5-T�V��$09]ʬ�r��q�K��S�U���%4!��A�����3B��>�\�t�����h������"-HFM�d��*ٙ�@�g���e*�Y��7UeߺI$�!rD����drDú�Yhw*�B���r���\D]#��E v�F�sẍ��1��n�2;��=�f#�ro^^G�wg{O9F2vH�'$��~ϟ^�      ��n��7�d٩�u���X�۱S�ǵ�g�����z���n��n�c�I�.�c.T\�W���j��OVlV�Ս<Φ��o~p:Gy�Sz��B��]�����;������V�jD�`��t��9�_T�nX�9�W��F���Sm��['Lv.��V�P:u3�����]#�Đ f!ڶ-�����	F�������p�!���p��M����O��t��7h�bSB��+��b2��6���:*���h魪�Z��c����C0�GuA��D��o�q�"|vy�nׁ����{�e��D��-*F� 
V>"�P�˳��&�{λQ�9�v,�p�g1"*���n�m�3�{3�g����g��3��_jSbդ���� ���{	V=�W��P#ƻ���󉔎�>��n����/|u�cjD������7�{vI$�2���K�E��p�fd�G5��e���Zk��GG��r��9�v,�p�g1A�B�~���O�����Cw�'u��6!��C����i�{�|�Y˦ͫ������{�     U�%��]�=V����K�[���ALq��Җ�D��/��ZVn-@�����	y��C�]UTܵ�)Dbp6X��Ӑ��ڪ�W�n��ϜL�[ʬ�r����"l�q���n���uM)r`�X�wP�Dd�Tk�1����7hi&g6�i�"��r�R��VC�~�:�}�Fb7��ܯ��j�$@F��w#ܰ@{�M�pwPt���9�r�axn�"*��e!~�r�a#������U�{vI$���n)��M2��H��$��uƲ��Y�8��^�׼�Z��5�K=d��Uz��kH� +��\����^9W���s�F���7+� �C1�:2��mշM�xV��V��"����#����|��B��\�vbk�3	�}Dn����m��O���!��Q:э$���:��&��s�=���=mB[�d�a�I���n\�P�F�����jط6wV�@�PwP�T g�3�q>;ҰI��s��R�8b�B��,��6��6�����o����V=O����"Kk��<`����\K��!c��ؼ���&���kE�j�դ6�^Qb\���{N�":�N ��.�>; �^fƄ����$��<p�h2�5J�"-#B�@�@KnI����[GO ��$q[ֱBZ�8��-�����N�{����>go�                                   �cїq�1�<�F3/1UnlF��!tn��z�C�X�|�N�N�vC��L��-ۓ��ܺ������Z�ݧ��#��tkn
���=��Cf,����<�;�O���vH�0��7\<3���g�{ k���/]�mXOF��Z5vg����+=�XĨrtݴec�Dv��+9�5Q^����6մv���6�`θ]��4�p�Y�[�ώ�����5����ۣ�][Z��۰r�]y�+����̽s��0��=1��)��N�+�ܝ�7�f�������}������v&7�2hْ�F��v�����Cn��p����c8I��xd�&k�\{#�s�8�4���$�	)�$"�	���m��    [u4��q��P��!����+�q۷\<ڹ��4�;:-aۆigr\��W6<<��6��v�|�UN��������q�q2�o�Y�yҫ=��&�A�!����3�b�LL�+�X��A�~�r�#�uZ9�őNl�#�>y����<����hۻY5m�,�j��r��Hn�����W-C���AP� ���{���`o�Tۈ^��#�nЧӒ��C�1��A�B�d���H�7^5��r��$���H�m�	.QF�1$$,�$�k��]ʴ׹���<3����Gjط6wQ�0�^@�{i�0��	@�(��@	R�q��J��.��F��T��1 z�i�u��q���[�89����}������ƀ`f!~]�ӄ�����;sNc�`ו��G1�T�b`X�hީ�h��``�焙�vꓖ�<7Q����s�I��s3-�T��K��W,�Z��߻Π��23���<v4�7Q�V��C���#֏r9�|�hB��F��v�5�-8H�!�����b2��5F����0B,�8]���)I$�I     r[f���w'�z6e���^Uhۍ�g���޽�Î�۱֋:'d7N�[����0B��%���aJ�xu5"ą���Fv��Z�[�o�d�k�
�9����N[���Gֺ��C�lS�cu���b4��s9H�~�<�1���n��f��*n,�92�5�!1W��Md����w"!���.h���",7�n�+���k6Zp��G�>��3�۶Ә��5�3�f!����+��#pn��ڪ�m�g�Z�*��
N\�xf#�G#�f!چۆ%�ՠ Q�y�[}��n��Ĩ`�A��!%8��> ��>�do�5�܇��,�A�g)��7Q�ܝ���|�]Ui��)��.�U�)�$wQ��.Ѿ˶Ә���Hn���r���Ps�#����~�r�#Á;�k)�9�A9J��PO�8���&�܏��!v�~��m��KD�&BĒ0�RÐ��W�LC�^�@��Xθj&���F�@�9L؅ẍR�3����s	�}u9�s�wH�7^5�7��o!�"�U�.�߽�     ���v�յ�z�*�m�����pt�cv�v6v��HCW�݋v�aI�n7�-ʺn%�n�Nu�޺v�����6I�$e�c2G�|�Z=���z1ˑᘾ�h���-�`�n���T�1]�O�F���ݣ"����ZC�[����n�$�Gq��M�F9E��M9
��N�x�d
{�[�H�&xzM�.����kD7���1�\�j����jB�ē��b{�����GA���n
���F���z%: �W5��7h��!�k���ǎ����-�z5�;C��>A%>�e��� B�� z9�4EZ[C�{O)��I}j�%��Z,�%��S�,�U���;4f��x�,b��bV����0���,����{���P�CWJJ#T"4)J/t��-Sn�N<�̰�m��՜��e�Kõ������4�w��ϿB ��мv=�{H���2�݀��i2Pw���6���x `rA���f����M���<����kq���:7�����4�<h�$+*�W-�)M8^���9h����N��s	�}�U#�}m�ݕh�ט��E��Q;���ʳ�c�֑qV�5ޖz8Ŏ�W����BlJ�ܫq�F'��@$�C1Ԣż��zL\����{ʷP�V��I$��0�p����q�ws�5���U��k����r��F�A�H���j3c�(�=�.�����\L#\E�[��Ҭv�Đ����_A�7      ^v�<�S�m;��Klݜ���vl:��G����m^�BVƅ��l��{tj��i��S�n�i�wɲ�JHd�G��*�U�Yh}�̏&��yCY7�2�:����3q�hC�f2�s�4��Ӆ�ܫ-W�g�I$eF܍7)��H��ܴ�m�J7h��h�gci�y��~|��b��	�C�;Uڴ�k��q=ʴ׾�}c�uZ9�u���C7h} ]��7�? 3*�C4ɺ��m��k���5uh*�b�b&FC�s���}��VN��j�{���B�����s�m��GqA�n���ci�{�s��y�ｇ��-���2la��28�a�.*����5���X����;Ux֛�Vz8ɕܪ�q�u�Ox�1�ӱ�;�S����FT���Cw�
�iѝ��\y��[�S�׼��%�4d�ɻ*ꚦ�
�ܪb�5�[Ϥ���u|F�7Q"�:�LO�Aq�F�7hM�7-HP,�d
�9���z1ˑᘎ��;�x�B����!D�e�I}��}ff      9%}�naطh��1f�L���r=�O'n�6��n-;�����Vj�\/>ާ����ܭ�|�ʪ�/V�y ���ّ�L��5�3d��	�y<�7����{%ǐ�ѡ�����4�x^�Z;�zk�nbQ�G�nR8H���m�J�,6�)ķ$E��I+ơ��3�x�aq���9i D],F����eTs�#�u�v@�Ӌr�!�"3�9��M�_|�ư��Y�?��H�F�R����.�(����U�����*�r�z�ƴ�97�$e��Udp������3�sr�g~�1X/'������/�nZ���4nѨ8Og]��n��e16�c
�aVw>�U�����#�Vz8ɕܺ�k��WUTFޟ�T��;@�۱��<��p�#���[��Y�``�N���]{����W��vxV}w�I$1��Ra�Wi.��x����ߞ�j_<��ݻ��T�!_��V�����ۭ��n-�Z���������"��UV������DO���:�X��")���X���$�?ﺨ�8,P @j"�B(�����?�
��uPqX%���f�Ub�@E/�����Z%;�������h�(��r~���~]ݟ����Ο�W㯉-=U����i�����4l�� ���w�~���?c�q� ("�ć����TS��h�_�߯��?��ߕ���������#���z��TP"������A���	B�k=�n	�h�W��d>ߞ���5W����y���2�$��~o�?<����R��U[��������!�(")��)	��n~�����lp%�~�QS����k��^>�v��Exou<z⻃��g�II����[�<A������L>����&����>/e`�>�8*UJ5U_O��Hw��0=�O����������E?O�FD�-������?�����O���~�K �DO؟�QS�g�?ڏ����?�5(`g���0C�,�=@�"�'�$!�����Q��?�#�vܲ��2.Ckn��eF���Y�.�6(�)�?_�п�~�D��}�����󾂿?���>�#�]��U�������(��y{C�EG�(����IH�)�����������?_�����k�����K�ִ��HW������to��}��-���lQS�>
�2Q���� W�G�w4_xh� |�|CUG^���4W���G��)����@�伂���
U'��%���J5�;�zp�*��(p':�����)��R