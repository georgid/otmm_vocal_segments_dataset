BZh91AY&SYZ����_�pp���f� ����at�� )@��� BQ Q@%(���$ )TI@	�p�*�     H%%(J�R!*�
��� �  (UT!@   P	)J%E N   2 � @ (2���S$�eX��s�+��]y��ʹ�{g}wf\���l�Ef��*��y��Ю']i�� K�գq��V�j���n�mN����  �z�i�݃ZӉ��Ӊ���r�Ҵ*AE��    Q�`G=uK\����c��9����V� �L^�MD�ܗ��4��������O��\����J���7]=w�
��<}��>�9��U��R�[q��k;� 7K��gbs����y�.�nMp`�� A@
 �@�M��=�^C�k�]�s�Z�s'�@���}���{y/��rj�8�U|� ΃Jbk�� ��d�=��}
��R�n���ꥌ׷�=����@�&&�>�^#%�Tp  {�
H   ����<�g�!��MWN@����ǡ��t9�3�|��=�2b13� ���yy4-� s��厍rb��_|� p	>����F��5p��P  PP� �>�Z���3{�x=�y��� <y��S�o�9����@)Ǒ�ӓ��^� A���j�� �g˃��Z��:^3������}�rV]>� �g'�^=(     ��m*T� 2h    �I�R��h��2h�F&�~��=U*�4�      ��U*F�J� 2h    ����M�T�P h@   B��*Bd�B��OSiCF����zG����/���?�_��p���G^���h  �j�$  Ҁ  ?�P  ?��@  �����`�   /�9b�  u�_�!@  ���@  ��P����&���?�O*?��Ç�O�RG�xX� F��#��0q *��2��C�Rq2L� 4r:��<�hp:��Eۭ����c�Kb�h0{�˻��k��T���s�{)@�L�� a��o����oJ�"��6{��bE�NMy	O��ê�cdi�ݧ����4�ȠH"��F\�x�D/}�H�+�1b� ]�!�4�%O�=���,�%BI�T�f��fg�㼭xfpFe���tC,^,�`�����
YP�yh�x����1�Q��8 �W�o�)".0��4����yy���>�Qn:�!�H�hjx� �u�g��xxa��ٸ�������h����sr�:2`! �e��+̿o�i
�S/�n� 2LL�(J2\�P;�zǚýu�1�^^g��x���\�0dہ�aAu�X�Ūi4.غ�x���p!��^�dN��2o*������<�m�b�8g��V�bf�}���A�ꉟtr�W�^ R���`v�W��������Ǭ]qs[:�瞜��U���䚃'e�K1��6�&f^F�@�a�x�{��t`&!CK�rwO^::�\�\�i�DA�'S��Z�ԴQ��f��,�e08�GBH|k�n��^ !��l[w�'�L� :6p:B0�6fk|ZI��gP�a=vw������ �I`-&U�\�i;�bװz��}�����s���N���r�ΰN��EE�BR�NA�zMǠu�D�6tn4G��J=�٠�&`wv[7��2�"�Ftw����5N�Լ�NZC'cw�΃PzDd��C�����ԍ�V=�B�0[��MSv���a)��k�YH
�Y�_����~���o`9�xE�ǘ�"Q �=�����	�Z��o��B�ܞ�f'�Շc��MO{�iA�Ey�j�f�p��6\ѧ�z� G2c�kj���7|�ܪ� �U � j��Z�oI�v΍\C!*hJ4BP2x=���of'}`h�p�&T��-V�`hS��i�`�( i���#2��hb�d ��`��8r�D*tC��<F���T�B��7�Yb�Br�]u���2�a��K�{ Ԛ�'']Bs0J0�r:��5ivj��0��X����r�4m��:�����y��%	BFA��P���(J;�~���}���ކ�X%	�a�2�z�齙ٛ:�38F�IC.9C����y���A�5����5	f&�5:]Bfa�:�%	BP�%	BP��	BP�%	BP�%	JP�%	BQ@�@�V{�y�x]��7d��X5mD�lx^zzf�Ǎ*`2��0A|C��<������g+���.Q|�87�'�P�xv�ƣ@��	33�b!	�p(MA�tw����^��Òt�!7vZ�7��sf��gK��h�
����h�%�@w	�{K���Y>�^oӸ�޷^�;#v��bm�'%���zrj=��q�i��#w�m,�h:����1^�&�'<cܻ�+��h!.�<	xI��c�2_0v��u&<(�b=������P_��0��u�p� ���̅T�@X��R^�ǥ�~> �����, E�)�OA�'��{V�T�Ao���	�k+�]P�CE")S���Ҥݲ��,��5�H	���g�e'�Jw�o;���<4-#�5N�0WI\X�4THBy.>�Ǫ���EP��s���za��x��ǳ�:�ͭ"�ŏ5����-Ed��`��pO7ɏ,1���w^s���<����#��;�F���]��p��ǃ���S�9�!@� Tu�Uw�	~��۱w�� ��`�-_��B�q��҉�@��
���iQy-4!��Ai�wۓ2�ۆ�ӣ)#$��\�tI�B<��������~S�1θ��Z��� x�c+�����@�%;�]����Q���h��5!R�偡�%�(<���=�MBY�!~�L�Ȫ)�T@�"x���0��-�x�u	�%)�N�=��(N�2P��g�P��|��d1�e����vf�%m�C`4��ByӮ�Ow���	�&v8FC�큔�1F�(�{ �{�X��0�<��b�:�h�,Plzm�O�P�C@�aFN&̃
 5	���xn*�}@*z�k�!���*�i�PbGm�0mfܧWb�s�,�z
�}�����6z�X����=X;.��h���X�;�����'���z�����C�x��n��S
�t�H8�7���_��[��:-{�|���0�C;����� ���%	�%	BP�'��M�<A^}`��QA��%�\�B�Q븖 ��}��<��X���F�c���`�{���Y>�
��х��xU��K�i�[������9� �20��%	�ݚ�k�0<��0��:P�J.c�:A�e4%�G�/���`�F�˺��Y޶Z�rѳ�=�O!<��%)�%!�'pZѣP��*+p`�9C��6�I�8ڸ���M΍l-�C��"�Q���ܦ@GP��I���!(vBP���AD]����;���٨
B%:5��y�{�[s��y1=Η%�!(J0#�w��pߝ�v��,�4դ�,a�J���8'ѳ�ݫUD�ޣ�NI�d�5�܂���LAPA!F:6s�I���g���(�22&" ��P����s1��C.	뱛nc@0ò�� f	'���
�!�G���Ə�]oY��}r�={�_��@%�d$���(J�jX������͙p�t��#	BD�g{Nh�
�ڱ�(Ҫt	�,{3Ҳ�Q��ѳ��1hJ��(J��J��(I0i�\zŊ�[���4�`��dT�C��d��:N�A����ݽ��̣V:*�x�pB4�@Hj21(�i���$�0t&tGAA��V�����jp7ٸ��۸J�C�di��sF�.��:+�����4�t�b�3�A�,�5�^��w.��u��P���<wt����i�u�����&��̍tvan��F�2��>�Bv|=CD :4�pX����݁�A�T��+4����,��+�����d_��s8ֿh�@�/�:���0�0�c��N�B#�P����lA�za� �W
���a;�0�hu�)]�\,[��v���==�����Z����t�=��"Pd���'��WgQ��F�@*����s7=21�)4�3B������Ţ;�Ϩ���� ��U@h�'�����כ%�7��j_������8bX���3Ǹ.
��K ��b���Ұ4�����ڨd7cA�{�Ae=zM�ʱ�@ heE �,eZ�wVB����v_�h5,�1ĳPy��'v��v�^�xaܕ�,�C���!B3{ە߇���8�Xiu	d�K"OZ( ��7�ó۾�h0��E�|w�d���KhS�j�#A�F jÞ,f��}7��3޿ѭ�;��X�� E�{���P��NC`�^��^�p��}������`!٢�#���%�H�&�7�!�''R��&����j0�!)a	B\H���=��2�:,�n8Ǝ���va����y9I��iup�va�;vj}{6n�ួ�������J��`��l��� Թ�[�����\�'��F�ۙ�u�c�&����3}2�h�=6��� X��H�
b��M�W��1XA�J$��w��\��S�i�8��r���0$.�(&ǰyXYD&���{✒���l��]֘�Cѣo5��ln�x�aI�P���}��V+hYA�w�s|����Ո �( 2=��~���w���S�.weND�{����	���'����ᨺUc��h�n��4�0��c�÷*�S,�t=�LХg���T��}��x�
$�p_�,x*�,��[9�|9}�0Os�u	BP�%	Bu	BR�%	BP�A��I���Lj&� �������H���$x�����#��Ʌ����6���8eǉy&'3(*�f"�x#�3 ѓ�F��RJ��	�fY�4�Ր��(#4ጆ�āT�	B{��3�@�"�:�,��1xZV��7�{�2g�����S�=��'���b8P�ׅ�c���z��M�����v�PT����㞆����¿���T�lF%�+1׽�45lZ�c�����d��`�*Kك/&�Oz�qt���*��(_ ���s3hd�:9�x%��d��èJQ�Qy	�0N�=��8�bJ�0� B�"ǰA,wQ�=���A�G*�)�=����� K�,y�BŁ�;�D�c"�H6(i� �08Χ0|�f�=�s¸&�&�:�I��I�������Q��e]��	�7n��⽡�Q�%f1��z�z&�$�{�n�~�t ��=�d߫HL�*ǲE�83H6d]z�j�Ii<�É$�2���4��(��&j��j���tś��7 �5\(�؞ٷ�=ʗDR�����y�0�D)�yxFW!+$ĳ̀�1ɞBPa��!�������`�Bd:
)"��y�4���t��N:���9�)�^E���������O�RN�g�bg���Np���&BP��Д%	@I!Bd%��΍���룰�5�v9���3�DK����������'�I$�I$�I    6�                  m�   m   \�m�6�6�[G��� �a$�m�i	ٴ�2�m�+t�UP�V  8�V�f�6�ӡ����m�v��z�۬�ٸ�`  �hjF�  !���6����ƽSJ����n[@��m/Y( E�   �շ    kn� UʠuJ�
��UUUJ�I�#��s�H�)u�E�p�����AUUT��� ���v��mm N����@��NP�쪫�\�AH2�      8   m�3 �T� �[FA�       � �-� ���m�.��v�   A� u��u� mp          
P                   �  A��`��    8     �6���   B5ٵl�I��ж�m���m�  ���8 p (0 8�� �G 2� �p\�2 R���� )@A��8�d$� 2 R����  �J� H�: d ��(0 8�)I            �    m�   H
�������K�B�ڧ���e�� �p �@
P`8 x��  �J �   � H (J�Cm��t� -��   �` ۷` ��  �b۶�N�����m��m��oPp �`[WMm�p6�I���I 6�m� *�S0U�U ��N�gj�=UR�ʲ��+���I��m� � @-�E�   �`�l�� 5�3m���$�`   �k��u���彭��79��jv�\[4q�[c��QRPF6��e���sm� �OԀ�UU�ss�ThV�Nm��ê��.u���e��<�7c�
^d5X�;�|�Z}���[�\$���Z�d��Q��U�Ŵ'K�h�k���$�X���2rY�Mw@T�����z��gc���%�IUΩjS��r�	&�t�l�v�K/B�hSA5R��3�T�K�]�@9���i��u�PH]7n�q�������i�mH��a����';�\v�U*�*����k���5���X�i�&�&��W]j���t�C\�-��@�^\�� �wm�iMy��-� �ArA̵J�d��Ik^Η	f�%�Y�����7B�R��\	��$�5*�KKUUed������6 6�	�%�	�m����l5�n�.k�@�v �`�-��$� �m��[��K� ���`  H�[�I��ڶ >���  ����n��ISl�l�`m�  :�mT���㵝��{��ej���¬x5��rn�;��],�f��#T���f�)+�L�q��i�yf;r&�FYzW&jQ�2�[TON�N2��i�<�e�啪T�Xg����KX��f����2�#��Z�Q�C�҈����K�� ��ڻN�н$�ΰ۸�-V��@Wmn0�q+�@� )j��JM�^M��$�[U/8�TJ���2:^�$���U�+i�I��h�0 q��I����[`A�͖�lv�%�`*ԫ;5�U���Ն�;#Ut%j�	em�|۷���'Y�:H@�ȋЃ��Pu<��m�m�v[��p KK���)5��/nZ�T�m6�t�p�mUUPC�z����h�I=sT$6C���U�MP�P *�����`sn�p}���݀���S�yj��P����l.P�ݥ�UU*3�UWS����lh{l ��c��v�Kx_K�Z-�Ŵ�^����薨��5V��5�9h  m&�9Z.rY�U��UT���a��v7SUN�tͬ����<��pK�R��I�0K{Kt�  ��L.m�n���i67��&���gg4c�[Gn�m�rYv�l� �� �ީ/im�u$uӫ��  m� 6�[R6�t�Ӗ�� �cm�� �nUV�����쨛fI�� �an�o[���8�p�C��S��5+*.�C��*�M<󽚠*��U��ճ�j��T�p�J��s��G���ʶ��4��(�WO=�f�U���N1 �;`ݮ�m9ɛm[m�m֛ kI$���׉.n�	$����EMJ
��Tl�T�N���k�&z��� F��R��xH;p/e	j�!���j{P,��}���R���ѷUŘ��y�V�i�W��D��'PU˲�\�-�Vԝ��PR��k��Sk�R�UW/�6����[���$�� m <$$$�U��K���Z��/[֤c��� �E��ĥU�` դn�� �  [d ��#^h�I$��6� ��m6�m����� ź���m��y���-쭀]6���L   ��m���[���x m�k��  I�-��6�i�&�Zm�i��`$ ֻt���Mc��`ݶ ۰pݼ(;t���[�D�f�d�:�d��/u�  m�8��[<ԯ*�c��_���ò��KO$�,T���]�MUU*������V�t��m�����mp[$��21��h ܡ�ʙ�Q�����5V1T�j�7Yݐ����:m�t�<�N9Q��m[V�:�YV�s4�&V��J:i���xwc��\�3��:��YV�Xh	�8(S�����rʵUTr�,�^�DݷT�z���u[t�O �Z���`6�.L��䠳��8h�fm�e�`�UUZ���Cf���KQ>�� ��W��$�l��� H���TO����+�j�U�e�n�nFט��\��mj��6d'U9T3d *��35mUѡN��]�%�eZ�P2�ε06�R��	���J��O��H�N��-�]6N���m����[� ݶW��|����n^�Ҹ  9��/5J��,��մ���R�Tڪ���'K���mղ�*�ԃꪠ�[�i �[/-+��&)\6�[Qɥְ-�.M]}q�	Qm���m�="@    H�n��Hr�mD��lŎ�۶�����l $��m����     u��-�J�ߤ��:Ͷp��m jGnͶ�����knl�� жKm����		   6�ͶH��Æ� �6�W]�m�%8
mc[CI���@A�	$ps�M1����*۶ �v� [D��rRmp ��� ��H      kX  �� 7m�ֻrD�K�0�t���-� mU�&��& �tqo9� �f� � 6� l6�O���t��M��   6� �  ��mͤ�-�M� �X`R��l ? }��� $-�䲭���> m����S��$�%p iX N�L�^�U��K@-�9��  A��g�ks`��@m�l@��ڝ� N����(�����U������Ʊ��t ��m�m �n�޸6٢Ȑ ڶ�8 �ݭ�m��&��xm&� ���a�u��v��kX E�v�^���J��   ~��~����9B��[@I�am��ONӺ*�]X�A�gB�յUQ�h�=�� �`6ۍ�m���$��( m���v��cT�6㦗F9��z��%���j�ۤ8�X'+jٶ���_ZO;-[TV�>V��(��*�z��0!7��#<U@����B[��Li4����   =Wz7iej�� ��X杮���[Ӯط�w`@8딷	�:�꓾�.3/]�V�+k�S��KQcţ��^�v�6�=��4q�ɇl��mWS�3�ڸ�*�N���"�S<���
(�m���욪���.�"�-ײ�W.���N�6������6�����G�Ù����������[\[�B�$NR�ite���d`�Pmʙj���dk����|�σb+�*�.���K@Y�˷mQ��h�؇h����sN5�%���M�:�K-���0��κzxy�i��x����,b��\��I%�m�8��� �v�]�m�Yv�v�J�Б��BD����f��ô"Uz�	�SZM�\��J�*�'+�j�ujg�[�Z&��-]��=�� .�����Ӈ[`!{uUV�mm�r�;/$f�RZ�n
��F����se��GM��lwU�.�h	���Jʖ3Q�7kl�V�u�Ɣc�	��j���8�f�#�؛a^S��m��Cy�p%��%�����Z@م�9ڧ�ؽr��y����v8�7���!�MY�ԣ�z��Fcm��<���n��9�y���m6��+��[E�4�	��.KW��E��uvb��{��w��w���D@���ˊ"��P��A+���?��~�W� �
���*�"�������D%�S�^�%�W��@��|E^ ����U� `�6��j.
��"��&* �	)�`��b &i�)*�D�"�'��v���<�HJHB4��Rt
�(����&��:�BJ�h�B��"f�a"H$ i�f(���F�LL ���FA���.����(���dD�(����� ���� T�:i�d�$���M*u�^�� �}�A�@�D4 =��B@Db �Q4(H'�0��"<D<A�q@4�.�<v���=�l� v� Q�dD=A
�`=���@��F%�f�|�\TQ�{����!�Z;@==A] �B'�	�dT�D�@:S�8����PaDЋ��B����� S]�'��m]��v.�~��   �?���������?�;?� ��`@Re&�a"F"�)A�eJ�ZU@sfm�`  � �!��B���m���f�]+F�V��k��J�N����l����Ԧ�
�v�VM#d�3E� �ò :��m�i�k	��d      m� �t�ۮ�Ŧ�P`8�aJ8 �����	 Q̀  ��RYxT�0)@A��
QC�%ݧ(�W���L���͙
t�l0[\�2�������kR�dg���堛�n1��q�XMq���qv�' u�q����\n�zSK������NsN�e�����뷉'�����[��s�H[���)㋧��ym�qR��k���Z2�^��*�a��z-l6���أs7$v^����큨�E���$������wm*�ג�[V�����s	�R�����΃�z�EU�c0:0]v�6&u�����0�m���7k��1���i�\����d�j���4�QӥU�8(��f�(��a��N��ym����a���ր�'��m�/udj�p�o �>����	ǵ�n�'#W(9���Olm��V�� �b��I�l�,�2d��r���u�8��9��L1��.P�q���&M���҂�!՞7:y0�N��X�k�t�ȳ9�;.��Cs���ahcuv<�b���㶝��Џ#�r�N�ۭ�[n���VںѸ�,�7\����{s=���U��g�|κ�Z�����
��ʂ�t���n��g2tL��� ���gz�-UC�Z�ٻ3���(檫lU�DTx&��T�D��Y�p�&���IJhT�U��U���ɳuu��2nƢQU��ڎP��n9t]RF��ɰn�.b��Fj�s�:®W�vneɲV6���WZHq�ݐӷK��ocN�ݶ�6p�����;H�IJ�q�kNz4�m�[�j�a�.w��%4aے}���v.����s�Uۜ�)����s�C�Z�s�ܺ�{Z�b(��k��Ş�ն����;E�UO�@S�PS�C�.x�v���M��hQ4��ٖ߻8�6|V�����f�^�fVa&�v�s��Wl��$+�c�@�x�&-X�Fm��7]9���s]�KZ�^1�.��
]����^�㍯h�R<I5�E�|u�c��]��K�ʐiwQ��.�s�v�M/*�C8mF���̽/m��n�
=і8����sY�'n^ִ87)�إrK�����\͸|6yb�4�;@P�UB��$��HE�]����^ۇ�2y8˃y��W��9&����w�P���d�f�	7�4�'ٳ��H�Z9*�t�%�HVـ}�|`�>0�Ӎ�}��,��c�`l�E)I���>0�ό}���>�>0{��$m5P��)8l��Ӎ�}��,��ό}���{��HIݴ�T&`�vV���o���>�>0}]t�߾")��(6����õ�=vp��yɦڰTd`�mv͎Wm�6�l�1���N��ό}�����o��X�ZGS|چ2�n76I���v((U8J�8�$�wAd�ޜl���8��Q�X��\��9�8�'۽b��P��~��}��}u��9;���Bl�7���s� �y�}�|`��G6���4�N$���d�n�6I����>��I� !�M�DSQp�v'9�T�(F��s�� q���g�e��ݷݼ�BI��!��V�L�7�|`{��ݕ�}�|`�h�2ջ-�����s� �{���ό}���֘r#����$�n�I���Ϫ����q�NoN6I�o���wmջi4�~��}��}��n�X�O�zŒ|���6���ۊ)��� �we`�vV�����:�|-����+���e�θ�s�N�lcǮ�l4�� r���만�9�v������:f����7���/u��ό�a��JP�SM��I�oX�Nk�VI���d�ou�$�'��l%#-:m��I�{��>ݜl�U@%���,���X�OVh����	*2I�d�n��&��}�ʺ��xr�_��h�(	!�) �]y�߹ʼ���ՙq5B�)H,���d�n�6I�}��>��I�ir�e�����F���w;6�X:�w��s�h�����Yܜ��ݮ�ڤݍZj��i��ό�.��7w�Y'7�$��C���
(�1F����`�ό�s� ��� ۯ���6��Dل��w6q�NoN6I�l�d�[��F�Ĩ�P0�cf���o���>�w,}�� xӬФ����-Hl�����?
�6���f[8��Àz">
Y�)���`nא]���=F�V�Z��e:�َ���pG$�Z��m�b���n�q[��3I	�Oa]h��ga���]�{b�pΣŃ�WFΰ�a�7�Ӹ���2�\�=�eG� mW���N��b�㰶�R����v�^8(�v��㑹�y\rb��gv%ܤ�:���gKvf2M��u�t��OK����U�kHaCs�����D	e3L'#�+��,0CL*+�G�wi�E�O�s��B	���m�;�kW'k6鎡�`�`z^
r�ʥo�m�����폷g$���d�n�6I��r00�Bn�2M�p�ׇ5$�L��l�f[8���{�u���V�C@+L�>�>0����� �y�w������Q&p�'۳��qws�N��0{���u�I�vӡ�I�`_w,�y�{���7���;�WX��|��n[��6���9��kv�pq�[�8.����>!�"k���w>X�Z��b��y�{���7���>��X_�x�J0�$��;�8ހ(I���G���[����r�]�쓹���N:�}
JDbI��f��e`_w,����s� 8:��T��$�%bN�����s�wzq�On��$�f��p T��m`�>0	_��C@��+ ���`Н$���p�K�"D���1��Gm�Ռ�p��5��#��p;��:1˵b�L�=�|`�vV�.��;�|l���98�Q(I�6I�ޱ��Ix�p�=�|`wU�I:MG�)I�}��=�8��P�E
(P�B��l����e|/EQ��Xؐ˶� ��{���;���}��&��&6R�0�dI!�N�N6I�ޱd��ܬ��Ӎ�sa��~�td���<�n`�n�s�������-�K��NE�	�n��{5�*�
o�߿����]׀w����l;�� J!�L5#i0�h��s�r�OgN6I����=��,�՛6���AR���d�Μl��Ӎ�{w�Y'9�+$����F�QM���;�8�'�zŒs�r�n�x
�T9t�d�h:��R5L�V�0��+ ���w���=�|Y$�h-�A"��	$ ��$�D���;�X�5�2�]������re�u�ظsena��m:�>�|`�>0{�{ݕ�|W�$u'm۴�[L�7��{���=�vV�s� ?x����]�J�%lm��ό��e`w>0��I�4��!)���R'� ��鵀{���ݕ�*���!�D:+T�i]�)+u�}�|`��X7�$��X�Nq,wR�
�#�c��ƺŝ��P��\� �e�H�Ym`�!pv�Qطa�B�ѻg��׬ٸp�� j�c����1�N�;�=��&��ܖ`�\(�5���8y�w�Ν�{iç��,���!豮'��ɮ���+�U�S�୞���_�8�*W:b��m�J�HtCX���\����e�N8.c����@DA@ �Pn4�E�8Q5u%�^���N`.�i�^�kN����"�՝�ę3D��j((�8I߷�I����{���ό���]�jݖ���Sv���Û�ə���{��w;�Y'�rq��(�*8l���c ���X�vV���{����I�v�wt�i��I��>�2�{�szŒO����̑�ن9�}�8�>�>0}���>�vV��Ԃ�y�73��ku:�xS�n�Kr���Խv��V�[t���n�j�������k������|`�ό����7���>���B�BR3m��6I���� 4(@T�!}ޱd�v�6I����'A�ܛ��H���� �����>0{���� ���]j�6:bH-4�`�|`�>0}���we`Z6�i'a6I����;�8�';�+ ��� >���T�mR:`���.�f��s��۳�O���a68�T��{���G\`2'q�������;�8�';�Ł����s� �W���I�v�wtԒ$�wX�O��+#w�X����B�#�4�����"��
�Xϗ|�w��P�4zA�K/��9��f�AoN��Ɲ��#��h�kdf�M�#��m�c�&I13BP����,��`˄lCa��$b�X�Lj�:M�3M��Z#0���Q9PY���k4Y��T�0�D�f�c��;0���`ֵkD��s��tX��]�ﳧ ��%���5��2���v�#`I���Fv�Nk�oy�yܺ���V�A@m8�j1�,&�b��@�^Ą��0F�3�M�
 
��6j�*�P6QV;�f����m�X���Wb,P�~�;д�b�wD&H��I��pݫSaElK1NF<u�D�s���:+��X`�E�AJ�i�e�sz]�&ְК�"&a��(xlz��	�;EЇ� x":~D\ػ���b/����ߎD �A	�⎑"�̑��	F��q]P&�$�q��+ƨ��{��)JRy��}��S��<�_s8���MV����!G��V���T��{��)JRy��}��R���{�qPD ��cv��B�ٖ�s6LY@����OΔ�Z#�˳k��r��9�f7��Uۖ�!���6�l��\��5@��o�:D �_:�<�A���-�>"D'���B��<c���We�*V�����z��;�^��R����߾��)J{��┥'}����Ò��l�2rj�eM]R�Sw<�A����)O|�\R������ԥ(ϟ|��T	�����RF��([6�9��R���w��)JN���=JR���~�)BHm|&!��H���)��I�ɓ%3BH+�I:��>��޶=JR��{�f�nl��]P&�C>ﾱ^4�����mG��~�`�w�Q�]�{�m�7S����p���{P1����ƭ�3��O�9�7^]s�ac����JS�����)JO}�~�Cԥ)����IrR��߿~��)JO�kB椛��SE�U�"D ��8�(�R���~��);����)Jw���]P&�+4q����RQ)r���)���)JRw��}��R���}��!BY��Ҏ�"��MU]�iֲַ�)JN���=JR�����)JR{�{���)O}��qJR��~&���A���x�j�|��Z���g��ߴ=�R�}��qJR�����R��g@��y���1�Haf8`�4E�82���27{n��۸�?{~Y܍�z�x�Kk��ᵩ�nܻ�qM�s�Slu�iqJ��R�m�y2X�j۟,lr��k'g���"��k���k9��~����p Z�DC�nfێ��=:;�vcb�cE�����t�;oj���k�Zf�1��/��󁸹Gu<#�x�G<t�%��l�camvݶ� �Kr�َ6��I���ۂa$���۱��܊6�a��P AUW�摌3%A��d��z7;M��o�{Ho����NM��ޙ�,��q���quP&�C�o��ԥ)���R�����pz��;�_|��T	�����RF��(�F��R������)JRw��}��R���ny�!,���GH��ɪ�5oz޳�{��)JRw��}��R���sȄ!fN7J:D �Y�l�B�Mp�:�?d�&�	Ib�j�5C7<�A�d�t��B����D �A��⎑"f&5$�Ղ�.��y�!,���GH�	/�B!�͸�)I��߿pz��;�_}�R������{�߃c�;t�gi��k&f�c���6�U�ZI�q��un��s�<������f�3s7��)GH�3-��A�ͷ��R���}�qJR��s߾��)J�8�j��iJ�����D �A����~=11�!LclC�����ls3�p �H��b���	�)(#1̜IȱS$IdHg%\fH�2�$�l��hd�����┥'��߿hz��f[9�DD�B[͝��Ww%�*�ky��z��<���)JR{�{���)O}�\R������ԥ)���L����	���n�T	�ܻ)O}�\R������ԥ)��o�u@��M�|��r$�nFZ6�دJR������)I��}��JS���9�!,���GH�=C�@571N�!ص)�ϱ+�z#���紗
�T֌�N�n�{k���nuS�����ԥ'}���)N��\R������Q�!B��g"D ��^EP���zַ����=JR������VrP!fN�Ҏ�"n��B����u)JO���V�Yf�[�5o[��)JRy�}���)O}�\R�� ���{����ԥ)߾��R����ވ��E��	D�˶+ƨ�Bm�ND �A3wx��B��v�D P�BD��'wiGH�a������YZ5j���R���Ͼ��ԥ)��o�R��y�}���JS�}���6�=����nD�6���G�iE;e7�ݹ,��Kp�v��<rV\v{��h�N�HK�4R���⎑"��9�!/z[z�)O=�\R���Ͻ��ԥ)���
̌��m�ۆ�5@�����)Jy��┥'�}���)W�휈A�4塗v��l���g��hz��<���qJR��>��R���)��B�����GH���m�˒"��Hn�T	���}b�j�*w��8�)I���}��R��O귯���hgÈ�l��8ێo|�)N���g�):���=JR�{����)I����JSϾ>3Z�_Y�����:�5���Kl�_�9i2�X��t�vS��/[Bb�-R�����=JR�{����)J��>(��!}���!BL�xˡ�H�!(��v�x�j��O��?R�������)O>����)JO;Ͼt��-�(�!6^��U�ԕ%�ow�)=��߸=JR�����)O�$������)O~��)JR}Y��MA$F�	9%������ԥ)<���=JR�{����	�H�HO7w�:D �M�QE)�WB.ꪵ��qJR���~�cԥ)߾��R�����pz��;�^��R���_�������rXX��gGY�^���*�	�nĮXj�t�	����]�n������=q�������ϴ�ݞ��F��8�͇��ݞ��;z6��ta�*�v0���m�Ӌ�f��m�ѯI��\��r����_���FRܘ�]h�ldG��q�s��.xպǫ���Dyv�ظ���蓅 ��i]�9�uV����.���r��������ԇ�)�ݑm�%ۧ�^�i��l�v:�C�=��R�Uɳ�B�6�4�G3f��7��g��sc�)����┥'�}���)N�׿g�)<���=JT;�?&m6�e�	BI$7T	���6���B��V9�B��<n�t�����h{F����3$q��k|�)N�׿g�)<���=H�d��}���)>�����)Q�L.jI��A4]U\�!B^}�ǩJS�}���)=����)M��+��h|ti��� ��@�J��scԥ)߾��R�����pz��;�^��R������=JR�xk�F�On?"r��4��Ɵ6qh{0/����\l�v�n�G���ȭ	��[�)JO<��=JR���~�)JRy�mҎ�"ٖ�D �A	��n���Ȍ-q��T	�ϾV U�6�.`���I2���T3�b	#�ӂ�0��3��d�5�"��o%)>�o��R��}���)<����)J{�ūFr���]Ԅ���!B^���GH���g��I￿~��)Jy����R��4=�� ㉱�$�ݱ^5@�N��\R���Ͼ��ԥ)ߺ�����-�Q�!Bo%����%U�a��{��)JO<��=JR���~�)JRy}��lz��;���qJR��|�����ޢ�-�nZzN)��\�l���un�f����P��`^�;�.��4��Z��JS�u���)JO/���R��~���)JR{��}��R���}]T��ՠ�WSW<�A���ڎ��Jy���qJR��~���R�g>�]P&�C�K�q"��V��lz��;���qJR��>��R��R��^��R����Ͼ��)�r�MU]�TE"��D �A=��pz��;�^��R����߾��)����u@��M��n�0�K[��=JR���~�)JQ�F}�}��ǹJSϾ��R�����pz��<����*6���2"�7;r�FI�iƗ��k���V�Le�:���ͩ=�����R��_{���)N��\R���Ͼ��ԥ)ߺ��┥'^�|���-M�N�
����)JO|��=JR���~�)JRy}�ڎ�"y.h��ՠ��D�������'�}���)N�׿g�)<�[t��B��e��"B�/"�j�q�p�,W�P&�g>�]P&�Cw>��R��~���)Bv-� b1)�8.:�<��}��R���}�i�%�q]P&�Cu}��W�����߳�R��y��pz��;�_|��T	��o��c�0DZM�N����i�!v��<��#q���[kn�L�����[���.د�MP�}�J��y��pz��;�_}�R������MP<��nH�,6Yq�u@�)<����)Jw���8�)I���R��"ec�D �A	�Ǜ���urn�35�o�ԥ)����┥'�g�}��R���{�qJR��>��R����QA�Wu0U�5sȄ!{����)O|��g�)<����)J7��+��h{�&>A�q9i[�4=JR�����)JQ�@��~���R������R������=JR�#��p��;��m�e��iNG��Z�
3.sEo��<eȀ��P
��C(��oΠ/�e޼�p.��f�fnNt��X	Jc���R��P�th@�@I��m ���4l(M0��dLZ],%�g\;�v!����sd��z��%�;M���w��λmh���c� �a�k ���Yf��v�4>3P��!�ۚ0M�dN��ݛ�x��6r6���!%���@h�%DKa��D����s]g]$ƻ,���AO�è�ߘ�f$: Ї^p<����6,w��kD- 4�@���"Ȯ�;�$�� � -� �g�g�d:t�Y�>��(
�^��vU��v*�j�U�]����g��F��nu-֫ij� ���n i�G[��	��n       Kx�����K�H��ă� 2l���)@�[*�@E��q�v�  z�z�Kl�\ٱ�r�� ���e����	M�I#)�RW�ـO�Sm�0�7�GQ�3,�s�ݚ	�Y�Ŗ,�sT�;'�m��ǭh��g�nhu�22�mYɌ�˞�#���{)���h˘v�DK�n9�:�k��IΥܽJ]Q������49x�͊Ȑ��q�1�y"�n9�h�h�Uh�N^L\U��ۑ+�m��$(���ڌ��l�:0����S�^k������s�e���OMP��h�m�k`��� �c�=�$'u;u�vY�X��q�ٺe^�*�:�Nn��i^���� *�D:���N��w�J���z�4b�8�F���f�g/OlݎɶN�9ڞ#1��{u��2ml�%�=��'X�g&��v�U��eyN^Ã9����9�蝜aݶ�O����~Zƫ�&ۭ���Y�R�'������پ~�|��wI*ʖk��hI s���L&�^-	��P��t�6��Y麗�O&���Km&{;�6+���c����Y����!3���5�M��Ǣ�����g�G�yB�
�ocK�)zWgt*�N�ʷ��Z�am��(my%ڧ��5U��g�g�9�e�);�@Ҡ!irҼ�[�2�ܪ�f�Z(�^�Vy^�we��c����fΠ�(�V�\%j㣦旁$8춸q�к4�m���d�0��ݖw���bM�p8Pʲd��Z݀���ck$���<ގ�IGL|;}�g��tvT��*�ϝ����r���{cnN��]ƎJ�d���\D���$g��V�{f 6�iծ�fɜ)��k�'�$=���1Y;6nn����1��a�n�5�3f�]v�z"(���� J��@��� ��qU6"�֫��kY���e�f�4���,K��Ȗ�̀q�`��j���VH�n��]���Uطn��s^�M�g��n��b����l�;���z%ǲs\u�F���n�:߇_w�yO��`���7:gyۈnc!�5δ�$����q9;v�r	X�ۃCn�k��A��-�u���-è� +�Bb��p�]H��(����8������{N�q���N:z�i&Pr2�UR�*
,���p)/9������ٺ�nʻ�9�On���\b�/���m���羵g|m��z���Ҕ�{�߸=JR�}�~�)JRy�}��^�)O|��g�):��=u��V�7wwueU�GH�α�"D ��Khz��=�_}�R���Ͼ��ԥ(5��|bm�c��jEu@��M���hz��=�_}�R���Ͼ��ԥ47��+��h|ti|��$C����s|懩JG�5���)JO<��=JR�}�~�)J�y�}���)K�����܅6Zi�$WT	�����W�PP���!B^���GH�=M��j�4;;��Z�8Q5$j�u�h'۱qp'�� ݥ�;�u�T��ч}�������e4�rK�T	����bB���J:D �Y�ny�!/y��"D'���94��`��&j���_}���8�K�Y�����șE(J�T����J9�=M� ��}�u�y�!D�>z�NQ�jn��ML�f-r���ޒn�UA�^�)"�$$�v�	7EӴ���T{�M�=K�=�$ZUWyIx�x���)	[m�����t��RE�w���{�M�>�JAj������Nu���n�4�<�p�R��L�pf�m�꽹���|k+i
�@�5m��)"�;�K�=��v!B�!DG�f�Ӏf�L��ڻ�]����-�������=�&�����- �!�I$�i
ա6�y��}�Uy���9vv�v"��(�?��P�� IBH]|�o��k�����2�U�%M]_z�B�Q�og�fV��@�Ss��BJs� x�S4rn%'�qws�MP�}��;��۠z.��}$�(��Ct��7v�����]nט���ظL��B�n5�<�5�ȥ؋�iշj햮�f-���ޒn��^~�T���@��F]�`ZL;I;�=�&�U�=9� ���h�%����������m�cOtNp�=�m�M�
�y[��37w� ���˚��n�*�����(�$�2�v��_�g*�Ͼ��������Bh������͆�z����؆���X���.����ޒf�����)"�Oq�@�ɉe�L�`I�#Ƃ�j��ͮ��#��Y,u���-m�}��k�a!Z�&����t�0yIW��=���	_K�6�$:h�j�6�@���ȈHz�u�=��<�m��B@�A]�-���n�V�0yI��.��{�M�>�p�7������J�]L����l%�B̷��37w��;g�W��RE�w˻lMЩ�I��6��!B���pz�u�=��<�~w��o�N��礳��N�R%,j�:iX�	f�l�F�sU\��A.v�Ý���\�]�^:�q����5���^8ꛀ��:�װ�������Ǹun�S���2��c/��u[�i���Ͱ9�ӷ�f����	�g��Hm�˸N�]��K�nù�N��2����N���tqڵt���57h\[R���������۾����|�׶�Z��n�d)�C�k����&�Rg�����������v;%ζ�8�yu�Q���x�qpz�u�=��?�(�BR����\q1%v4�$�u�z�$z~����x�$��I��z.�Vը��t�6�7��yt�ޒn����""Of� ̭ݮ�x2p�U7w3TUT�7w<��m��}����ͻ��]/ ����i�C��V+M=�>��X���@��K�=�&��\���6��#�C����#m��Ǘ<v�l�96u86:�G�]�{�� ���Pdk��{�H�yt�ޒm~��I��l�g$��B�^woĝ��+ڡU\((���/_z�� ���]�P�)�R6n�rfn���U%�U\����@���p؈IL(�������xqxYD�%hmݱ��ޓ+ ���h��x�~�ޒn�W��1%v�:��n�yI������^�I7@��e`�������ՠ�I�"�b�4��6�;6��l%�Gf%pn��5����v���$��ۇIRm�<Š{˥���t�&V~����- �_��j��]�� ��}�S
�ٻ��3+wk�{Վx���N�4Z�v�{�}�2�yF뤨P�B]�U
"��}�����<l�����WP]̕5v��D@�D�V��@̧��=��z�IO�w��}�dsu��ML�w�1h��xU���&hzL��RE�{��J;T�[n��=�J�9�L�n'��	��m]zX'X76���=���Ѹ]�Tڈ��qY'w�����e`�-�]/ ޯߒ%!T���4]_z�o���!
R����3)��y���	)�������®�m3 �_���@��K�=�&�z8`����j2��)6b�Z�ߒ���y�ށ����iJ6�P�F�31rɊ�q�#�D:RX�q%깻] h=,����&�IJ�x�$��G�RE�{˥��ߟ�~v���ߑH��UOl�����9ܥ���S���6��wڗy?^��t�ڛ�\�I]�m�����)"�=�����߀����{��k.�_���i3 ��n��DəOg�fn�z�v�%���"hn��;J�f-�]/ ����}��{�H��Ae�n�+T�Z����%{;���ަ�tJ=�����]�"R���COt�0z�u�=��<�m��TT"PAIE�� !LD�H��p�D��p�0	��")k\�Y\���{���v�7ky�j`z�1y5�Y㫠Z��I��Ng8PZ��6-"YWW��w�J���Ս��a�tnq;Tn{��c�\� /8�轮^6�m�]��s��L�`����e���q��ӞE���]1zs�6�A�M�f����/[��<ltsv:7�Nq�̷:q,v�4�fs����Q���c�ӣ�<�.�ɹ��=vmzX�l\�5n��d!�N2�p�p���sj��^xK���Dێ5�7��m�[�r]vW����VU�j����
�I���_���@��K�=�&�z8`���HQ�T�K���W@�������37w�ٷ� ���]P��,�UUU�Ԕ�Xۼޒn�����)"�=���'�.���L�m����'�A
���8en�tz��T(P��DNf���k�*f�3WW5u2T�Y�=�m�@��K�=�&�z8`�EJ]]��6ݡ���/n��$0j{q���x�sW<t���q�������ɾ|�c�>~Š{˥���t�0yI��H,�-ӥi�V�w�{�M�S��� ��#@kZY$].��Q&���L���JY�ԸZK �-h�4,���5C�֐ҿ"!�����v����W�kϾ�Uy��]UP ���u&~��n�s�$���=�m�M����̧��37w� ���l�ۉ ���d��@[��OwՎx���CTB��o4��ӻ�'l�����1f-�]/ *����$��G��#�:R���j�q�BI���?��wçY���:��cu��l�
��cAV��I1RV�mށ�����ގ�񻄔tz�� k�e]Z�-]	+�M��>�p�߫��#�=�����t	� ��]������I3 ��n��X�'�ش���]IB�q:�����Yo5���
̫W�,< :m� �:�bPhW�ZP9T:��>G��m{.�s7�4�l@��b�*a!�_�~�I�chq�vw���2L2р�4�5��p,�Y�i�5�B��"��Ay�|P�`@�)`�1��LQߞ�ރ��4b���5�0;�������d:��4�}@��x�>�]NӤi�EA�x��00�sY[�Ѿ�v�'p�{� Ц��Z�4�tl�&:��tx���k�@<}Rq�HkYΒ;,N�2�]�>,J�UD
 ܰS�ܢ��Y�(ɕY(�}�N.�=��iO,�N���*wf�N��t h0|�]k�~B0.�U��iay��1Q�0����4��s����6l��5��P:tRe?p=P��� �E���D�E�C�C�D= �L(P�CP�[������:ם3#��U�sUٮr��)̷��n�z�v�Q��n��6W&I�j���-ZI�ޒn�����#�=����o���*Si�"8 !��5댭��;v58s�.�d�pW�2���w���þ�"�V�����G�:G�{˥�B���Q �w{�'+T�L��]L�i���:G�{˥��&�zL��TIߟ����
,%ۻ�$�����t�&V�#�p_$�b��Xۼ
�ߎ��t�&V����IF�� ������9WǞ��iաӡ%wi��ޓ+ *�W���@����o�b$�cSJPO���U�>$U�ۭ�t�ۨ#C�q�7���h�a�Ë������� ���|�w�d�ݾ��V9���z�o��u�:.�ȭ�T�v���z��^W��$��I��z�H��Ae�n�!!�դ���&�zL�
�UG�t�@��K�>��]��)����4�@��e`���@������o� ��SR�lI����n�\���.��w�����Ͼ�ʶ!�G@�T�n�� J�*-�'e��鴪��I�^�l�%�6m�q:$����j�H�u����=e���+b��88��H�y�NY6�W6K��l�#n�w@�g��l���vh�5��DR���J��yq�K���Uer]�;nڒ��g���\)�s����e9�Zg�I�jŖ2V;Sͫ6��ݹv;=����@[�;n�d��U����*N��F�C���ݭ�t+ۜ���u���ܽ��k� �C�N����7b]ڞz��ݵ��Z'�4G1�{���[VbmU�b��ƞ8�_����t�&V�#�Pp_$�jĭYws�3;�P�}�����w�=��<���(R�K��M�TL����{7x���w�{��o��l����ю�r&�� ����x�w{�w���}�2��苻�+�2���|����| J_�D$���π�e`��= ��R�7j�4�
��V��F��[8.�&⼛��S�j��l[,��$$'v[��Hh�ZM��&�zL\��I(�B����Ƿ�=�I�Ѫ������@�|�r�IE��Q ��F
�~P�@�/s�?~�UX�o�{1��b"aD~!B�(�P`Ų�)�YwtJ����d��߯��;��(S8��z�7k�}��eԎ��I2U���|�U��M -"$	����{��w�}9�`v}��� ��������j�n�{1���

?$e�߫�d��߯��;��%ȉ��Xm��.���F-����S�hZ�V��'����� ��n�4�`�=�N-��d�N6��;ℵ
@�R��z����4�~v�!&����@=� �c}�O��Y!D~"" (=���&fO�7dUپr� ������ӝQ	
����|�p�������J�WB�.��j��
j""��ow�ӯk ��H����{���h��U�:�]_z��� �"(��A����t�xzI�ӉJ��V&�um�:�5�8Nts����҇z�-בۍ�m��6b�n����ЛX�t�@;�/�g�}��!(�(J|�^� ��)F��M��դ��i�h{��;;��� y�|�A"(B�@�Y;557RUM]M����ށ�΋ =:L��G�J����N��3F����I��T�YF�~{\ �{��{�&�"!� !�e%��C~�������]��M4�����N�4
��*��B�HP�/� y���K�\�����ɮ�s�.�X����͵�^K���H;N9��i:"��w;�v��u8Iy~t5��fh{��;�M�>��e~�_�R
IU��~�U{�������4*V�"�o �I7@��E�}��s��|����*B�����"j�l����5E�����2o���7� �txzI���R�J�i�*ޭoz� ~�$�		���~��:<�$��,�usi7Q2��f�wW�t3�!%��"I����=;�\��w�-D(^��n��v��]'��$9�nFuf�9��f8�-bF*�h�u�.�t�:Z-t�˺�\�wL���A��h5ø�E/&[F�M�4uŔ�G�gx7<Bm�l���ks˄�ͣœf:�i��g��6��UK�c���07i���C4jy�y6nbۈS-��'W8n��S�ٲ��AK���瑩���� ���k����]��u�`�����Νp<��1s�0�r�����I6�J6���Q�Ϸ=��bd���~?���~��ۮ�m��I~H��Q�	'��?����M�S��T�&��\�������f6��"� BA
"Mkt���5st�&�E]� 3ww� ����&�\�`+�wdV�i�o]k9�s��H����, B��~�����߻�>��p?$������@��ٮ���J�TMU� �m��B��"�J�G�wk���� ��|�a��6�p�S����n�:xᘳ����:�#��#�![��ֶ덎�îs�].��m� ����3�!-�BDH7����4�U7D�WhT����U�}��o��~6�2)C6#"�9�+%(��'�*�]W_s�򮽒n����\�Dm���![�o2����co�?(D$�	D*2~�\��߿_@0�p�553s5SWSw|1�ށ���z[n�B�HD%-�x�x��4ؓ�T�&��\�`�$z����M�=ʹ4m�]dp��\J�N��W[��l�<�ql�7a�u�DM�� U,]�Ĥ)�d���������w�3}��o �W�.�ȭ�T��ۼy�;���HP�D% �������6�4�\K�um�t�i7�wN��_y����Rz,#��l33�B�D�W&���	r�f�(�J�	��Ĉ*��{G�?�X�N^����7v���&��TMQrT�_z ���I�4wG�wN��!+jf��R�5W| �x��Q�(P
"u�� ������ lŊf�PQP���6W�����m��t��we���w���WD����P�Uci���� L���N����z�r!%�I( �	Hd�� �
����ի�v�M&��$���8���1�""�(��D�����*�.��4U���nm��=2H�wG�wI7@�)�;li�T�7f��ܯ�Ad�aVX�BJ�������������<�� ��08	���}\�Ϗ>ՙ�}��R�Y]��� y���IJJ#�ID�ȁʲ�����U�}�o��U�3@��T�HV��`�v��[IRsƵ]����]���;fס�Z.3k�EGh��\ұ]:�V�xt�t	���L�	��z��Z%"�ݪv;m�=7���
H0!+��~���� �����M�����v�&��UY�=-�} y��	B�BB�DKz��soN�X��wr��T�]�]����u�� ޽�@~v��K�!������)٩�����.��f<}��(Q��Ӡd��1�`z��xD�6�m9a���)d���2Ha����,Y1\#�^�p̵��Ė*bH��Η2�c�DD1���-{��%�ad��i*�%�@Xڒ�"o�m;p֬( ���]	��Ib�ؑC��DE:KW�dמ9fi�%��0�0d<<\<I6�̢d�ZL�)j!�̢`���{$�D��I 	  �� ���d\ۡ`����u;[R��V�y�R9e�U�[ �@r/N,�]6M��*mv�&���(v����[I�e$-�n�      	e�
Q�ל�l�kv�� �@
u6����A�^��ā���  �/Z	$�+]3l�@
P -�۶۵�8$$:-�8�;D3F��J�v����KQf��k����lh�P%ņM����a�r�l�Ύ�=��y�&d:���u��+�>���p�[�AƮh�hVxX�]�^�u��\��y�l�%��8���[Y�w[	3�H���:���[n.�1[�!&8�9Ԫ\/X�t	��m�=�XW�1��A�᧚��[L�e갲���n9��Li݇rd�B�p�ص�=L�L;йpl彤�ơ�],��S�Ϯ�	n�"-v�eٱY ؇�0R��� ��%�֚����A�C'$�fˋ�v�譛y�}p^��7�NΜ�8�۞]��Q�m������kl���v�FLYy�j[[OI�e�5�$Gf�t\ʽ�I�X]�����V8���fѭ<�;��km��ꎳ�����n{nCGQ�qq�um�2����X�Y{U���e��R���]4�;������]�˗�Fթ�֮s�%��v���+��m\D�Sm����
֐B��c��j1{Rs�ڛ�����]C�������l�lY����vZ�k`�!�iPwvm�5U��9��=�h��W��eڪz�W�/+̨M�x1uJ�"�c����G�L��Dq�Q�@�/;m�{j�>4�=���v�ڠ��;�v6w[�LlcY�׍�8z�n�\p�"J��<�����ILs�eg�ls��X���/h@5Ȼ��I�#Av͗�^���Bwj�-Y�>�Ƿ:���ݵ��zwN����ct.9c��Ňjw-Xɭ�3h;��S� �=@H�(t��v��WD=�`m����umq�\�]Ac,U]mrd�Z�jbM��]n�e���dSVΡv���j�i4�ש�C�Gl�+�9nɞ���hMl�6�B;��1�5�$��7Ǯwnq8��%c9���z�C���3�e�͇��\nݝb�r���^;����A#��w=�k�ۻB�gɫg �;tٻ��2xT�����r��x�c��c#f����"{H��=X_]���wQ��m۫�C�s��;�<�Ol���v�\����~��8��w��:�B�$�B�o^�?�����cNڤ�M3 ��#��:�����l��H���B�������?T�U�e�s��?N������'���G�}%�X][bT�MIUu��(��BQ[��~�@��_�z\�����=��w��)���S��Ot	��z�H�	}�`�&��R�{�Z򍹢��/<<�1s�^-�l��^�;I��N��ƭf�ֵ�8��ZD:ݻ��Ʈݤ;I3 �����@��ޒn�<���us��7t�
�coU}�����I@=��pѱ �w�{P7
8.�0���1���Z����(�B�!��K���ࣹG�@��G�%�(J8��}�oz�ݞ�x��Urզ�ݫHi��w���?Ss���H��)�׻}e�� ��4؛�ҵI	����\��/�,�$�����ݫ�;VMM��K��$�4P�i�� �w{�'���wq*(�;�P5WMQrq^�� 0�g����7���^`*����P� �kS�Lտɔ;F��z����t	�%�U~��z�H��]ł�lJ�!իk �I7@�R^�#�%�E�}�Z%2�ݪv;i�<���:M�t?3B��A�o%0�ĥ��!�&�	%#Z޶x�x��D@(�^>�=������T�L��+�W55s��
r���@�ok�g�}�
#�!%��<6�w7S�wLV�Su�<z����t	�%�K��~�T�SS�7%�UTwa�ȟ�?�ū,���ɬ�!�)x&��=n�pm���'v��i6�����7@�R^�xݥ��:�a�e��Wh�SUhM=�'���z�H�	}�`�&��"���T_���޿�y��v��5$��� s�~���1� �6�����~tUUH�n*�\�پr�J#H�!DB�ok�<����nxQ�%_�R�>z�J�VحP�V�I�<��@~��z^7}�c��D%������Msb�[��l�مh�NF�6�v�0�;͞Mou�f�ѽe�n�����L���	*��&��I4������~u�����=_tXzI���R��nj�+�������J��B�%$R�H0�����?~�5�5��������X���]ܫEUe�6�����;�M�'���z�H����-ěi��r;$P ~T B`dQ���JB����%eT>����uW�u��r\��/�,W�6ݦ�V�К{�O)/ �Α����;�M�:^Ǌ����`�c�$$Դ��8�؍)��u���8�3��]A�
:ɓ�:�ͫ ��v%r��VӤM$��.�%�)�]���a���M���j�Wv9.77E���@܏<�v�Pm��v��)��N���;i:@���T�z�)����kd�ێnI�e�8!��v��-����n3�x�N���.��<�g���؉�MЪO;q\�c��� $��p�����ȑ���J��?(I�BP�%	JP�%	BR�4@*J�J�	H����C�ILL�#$@R�J�3JQHU4P"U%ED�P!�J-0T��EJRTBRIHP�2E,ԅ	 E$�BS-(�I%	R�PQA��B�AD(�AKAJ�4!E P� �41AE@G}�4a÷m\Y�";u��',�u�9�<�y��RY��p���+��U�s �~���n�9�u�3;�I$��nm��>��*��ڛUb.k�7�s�9�uĔ/�0R$�JJ�
���PD�B�
e}��ߺ��zp��@~M:�R]�Қ�%X�XzI��p�~�vwH�	}�r���l�,3E��9P��BV@�����r���~�΀�1��B����@<a�ҫ�&����ֵ��W�{���C�BT`YHH�"BKi�� �w{�����>vȟ�2]ctr\�q�������{[Pۜ�gu�Y9�#��׷��$���+�_j�4	}�`�&��K�N�4	�_ȧ
m��1�����{�PU� S�E�x ~HD�	E������	������	\{��bn�uj������nxg��Q��IB���e���o{�1�t˛��7eUJM3 ����	}�`��n�=0��J��V�7�v�Rx�	}�`���!	$��{π��Ӏv[�}�S�|�G4<R𚺮��v;1N-����Ml=�4i�b���u��݂�<�H�<0Z�&�	:n�=0�:=_tX�W�L�e��I��@���U�""?D�Pz~���?N������ ���4�v�;�i�ܝ��{���C�1	1�"�U&R�J<�qDB\�����[8u�.n��ʴUM]U�&���~�	D�7��ǽ�x��
S�n�����	��M2�m`��~�_�z8`rtz���\��\La�����ɣ�OƼu�(��0�8�I�y=2�@��9�ء��*un�U�m=�'���t��K� ����������Չ+M� ���IDD(����������@�R^���%aE7�iio34v;��}�
?Ss��t��X+v�I0�V�x�&��K�/����i;D^�U�^s���W~{�Պ��Sj�������J��@�-׻π5�� �7ށ���D�o��kG�n�\OZ�ŉ��މ;��F܅7>Wݷ�k:y��g@�}�ߏ�@c� �7�Т#��ݞ�M;��ڹV���&�O/���w�Q
���BD(�߷���ο~� 7��?+��R�L������'I���N�4wG�J����V��M\�_zB�Z��n^��u���<N�t����ӫ���HM� 7��~�
	/�
�ۿ��~������K�;��"�C.�:��v?i,�MΊl��1����$
�+�I!V%G�IN	�ڎ�{:y�!t��I�������{�=�4�r��h�Ú��镺���{/�s����n���W�kԀ��us�9W�������{�@��&���Ʃ�s�.0P�� N
�K�V�
9�����3�뛈�x� ����=�X�]XJ�۔|�3>�%θ^uz��E�������f���a
^S�E� [� �Ð�qr�NSj����Z[�� ���t��O)/ $�3@��Q`�۲�$�I&�	1���IJ��I�[��׻΀<�|����L�U�&��yIx'I�;��$�7@><B*M"ݧN�����߿UPI�f�N��	:M�'���H��m+��E[t��y��wG�I�n�<��\���%:�ޓ�;y��zx��,uT�u��6�ֶ9��K�k]��o����;w���Ј��6�	:M�'���K�#�	�+�tlJ�[�Ui�Ot	�%��_���P�B_BWc�m�@r�� o�H��A�SPv�uo�ؐ��\��N��	:M�'���o{��"�le��R��9}�	B��:�� �{���K�%Α��*�X���R�E�I7�I�n�<��\��N������6���E9Qs\m����xgA��ru�J��9���5��������a�u�Ub�I��@�R^.t�@'tx�&�yT**N�[�t�[v�w�Kx���;��}����D$u�ҹLtSM;U���@'tx��t�����;(�}�z������2N����!����hvr�|w�y��h�:�`�f	�5��1�t.�)�wln���Ȏ��u�]/Af����,ѳ , ,X1S�\�Z���afh�c�d�	��d
6؊�4~a-a���:�LΫZִM�޸�]�u$E uP<z\�Q����8��L�mu��u�(��s^/m�c�'W���J��Gg9�q0�v��E�����x�������4&fNsaaZK9��h�=5ke�Nb��M��$.�f�5�Eav��A��`,�0�,5Q��tv�a���f����-����0�2#��э�c�zt��괸�ͺSZ��?�����)���{7�J1(�HI�/H�v >(.����� �~P��W�<�_E ��Y�{��<������R��,&��MR�n�o ��n�<��\�@�_��<W�4�%N�ժI���'���K���� ��7@�s�pi6�.�pܢ�7`�8��q�Lon=�^^'����I'-��חF\����~zG��<�t�����<����BSC��$���]��/�1�?�"&G��z�n� �~n��j_$�.fj��U$�xN���*���=#�'.��}��w���T����K�:��@yX��P�*I+JD�W�<�Pz�B���U�hv��I;�:�=���x?c�@~��<1b���g>��T�l�;Y�g��9-l7�bɭ�/[m;�ѷ�]��0��1e�Ոa&!B�˞$��^��7@�R^�=�����aT�jiUPU�� ��}��0�I�[���=���� xa���U*�ڪ*���z�7<%����Dκ{<�=�@���.n�个.J��灩$��	L$�g����?mo���������^�%b�݌�ލ��r�x�q���[��2_��@���� �LW$�1�~��;��7��.��8׮3pXk�T���3l�rlU�+T��qҽ2;O`C\��l�c����=��]uÈ2�v�q�m�����1���x�sn���{=>���擜��vM�tu�slJ���Ξz:ު.p+����&�R'�֤L�n�3�q�0�]�V��������ًk��qT��ۓ�t���V�C��c=N���d��	Hl
�T(!��e�k�,J��������i�a9�s�������wVW����w~���q��͠.U��������l�/��<�s�7�~��j!�/��6�@����3�<�s�1�zD%��R�Zm*��.���զ`����������p�:/W�r���&����h+�~�ހ���jI
G����Ȣ�_�%N�BHn����p��������(�j�.푄��XDO�Yú읯,���kZ8�S�{u�{3�WtLi;WN��BT�{�OG ��|�+���v~�{��~W_�R8���I�$6I=�����T
*��P�]��|� ���?;g �W�	X�[C�w�o3@��^��7J��=0��f�=R�e���$[���N����p�������߻�ڈe�N�M��'���(�J��|�{<���g�jh~a��8�uS���x����tu��^�3�^I\O�:��S�Zy��.���� ��|�+�~��P�K�ͽ0	����W�Lc���x^<�r�x� ��}����~�΁�8�M+Uim���7@��z����/(��(�y��@ݭs�c.����$%M���ߧ�� t�L�'s���7@�|Km;䝗hf c�|�2��1����l��B�y���ݿ�ќ�v��ObN+ѹ��t���|�c<���_��̹A������)�}:ϭ�<π���OI��p���4	�2��v�-Ҵ���t���?;g 1�>t�l�D�z2&i�bv�'M����K��t�w8`�{�x�sP��É��(�-����P�_�w�[�8�����$l@#b����A��X���c�0���-8�;p�	I�2qO@ �������>�z�����U��V��X�4	��U_Ot�yIx�zL�>�)QJ���$bE�l9y������,�6�$�v���jf�"�D�Ȉ���U6�MPU]�ۏ{����}���(��5�Ӏk4z]'j�[��Ci�<���߀;�I��p�>���U]��Th�eڲ�g�o�3-Y�����z�ݞ�^�%b�41~�zZy�T�p�>��������O@��&;Wc�����}=�t	�%�}�3@�����!%�!K��Xv�
�(=Y�z���.�5g�y��,$�]9���T�I�i�R�K�z�Z��n�"� [cv���ӹJB=�����N{(�������L�n��ם���=����]��a��u:�d��O9��h�v��vO@��!̜��l;n��9�tr�q��W��c�����nȎ�c�=B��=%b=9��2�y���g�֞ʳ!>{#5�^q�GU�ٙ��М�^�۷m]\�������ea8��x~��]�Co��m4�@�R^ wޓ4	��}=�t�\ �;un�I�i;���f�;�0��n�<��Aup�R�j���<�w8`Oc�MI(�D���< ~��t��l��Sj��U���I)��ߺ�n� ;�I��p�'�4��an�-�����wޓ4	��}=�t?����,;v�dω���ܥ�m��	��Q��wT�r����Y�tS�VjՖ��}�3@����7@�R^���J�dhb�n���4	�Ꮏ(�(��I$���>��nx�y��'�\��$�ժHI���7@�R^ wޓ4	˥����]��P���i����%�}�3@��^��M��p���ջhM'E�� ���=r�x��7@�R^>�R���`�Ѧ�:'*y��+JCv�C����-	2<F�S(�K) }.7u`��V]˿^V9�?c�@~��c� ?f�:��~���%J�
�m���M�'������@yX�&�G��\��3j��.���7+vx�y�t�Sp�D)D	X�'?`��'��hriL3�q��KA(�N���a)B;�蠠j1�J�Q�Og�}�7�1T���KT:�t��� ;�I������7@�R^�+�$�A���WZ�ǠN]/�l{���ܭ�������햍�hx��5u]ng9����f��`띗j�Yq�i�Ͷ�O$�1����.X����@~��z~�w�V9�̌��tX�VU������ny�	L�>������>���O�DA!�4�W6���4�m;��f�;�0��7@�R^!)ʃ��˴�WX�c�'e��{珽����P�(�)Ee{^�@�Ј��j�U�L�*���>�	�%���@����Q`+��ީ,�<�:���b{q���P�v�n�P�]��^���c]I)d�0�o��m��������	��wӦ�ԯ�m�e�.J�n�z_��H�$��N ���t	�%�Һ�J��C�wZ�Ǡ<�g Ϟ>���w+vxN�����̱�bT��ZBL��wӦ��K�=N�@�������V�V1:M��@�R^��tz�p�=�����ö����
��`�i�
f������lfPh�X!(b*��
�:1����ږ�	b�����ÀK���1QA�DQ	RuR�N���i��e�����,��$�bF2-c�O��ݘo56i��iх��`�#��)���U�X&Ն�YF�(4^ ��0L���0�0��.f��0Ҏ���S���B��!���+�`$$ (`��I`H� px�LAC�PM=٢	c.u8���h���0�(2gmw���atXk#T���2,46$ņ�\Rsf7y�L��� QD�!A&�P�D9Օ��t� �V)h	�5bK$L��h@Q �(�B6��$�$��I H m��8 �ukT ��º��Cu��KT��ܘ�v8��ڣ"�Usv�̜��U=jP�B�� ���۶�l�k�L��HIl���    �i m�����4k�����"@�g [@BE(m&�  ���`5MXP`8 p��)�u]]U7�	�v��Vb�UKɣe�9]-S��H�].5n����C��R"�b�I�칺�z���kƸ��;�����k%������a:ڱsxphā�-��L[s�-�s�U�s
�1�����6��"��,��0I�,����VU^]n�,�����b\�\��Ցg�vq���N���j�6��nu.�S�K�j�졶��y}v��O��6t�X�۲�\-�b�Ƚ����;���͎��9�b�gi��^|=�Z6[�.1s�΢ܛdyZ�IcR�R[J	݇�7Z7��;8Ӟ�ػf�g[���6�-<�!�K����˓GXk��M��3��t���u��R�j�nڄ;Sc�m7R<&��g�%�
�26�g��� �����{;[�aU�KY;�*���q�(���Y�)7A�n_d>�O@�[�l��q�[9��2�Y88t��c�3k<ƜY)�񞮻`�����.�nvR77v$�����6�94�2#�ʵ�{j��V���l�\���B�¶�r�@;USp7[<�v��W�ۚ���/0�h�)a��୶�(StZ��`5���$�lHHڥ���h�VuF�v��3�e1�,�V��<��k�ѡ�m�x��"w(���l���d�Ɨ�ˮ�y�uj�^g�e8�Ky���Ş+�nt�ݣt�,�`�X�٭��ۭ�n��{Z6�m�ƞ`�l3�8pȋ&㸶�8�y"\yõX�7q��Y��[pN6k<���87�D�ܚ�s�T�"'!R�C��q����jv�8��� Ȟ�=�h��� �O
(U&O�`�Hq�*dm$�n����jJ��m���pl�m$�^�gMo�p��`��B���{5�p�&�M��Ch�7<�������]� n�u�8y�Ӽ�;Gb�ܯWE�,�sYq��Z�\X6� 6�by�>�OXKI�V��Y�^�i����bŢSi��s[[��e�w>]s�蜜�uv�5v��q\���s��h�6��T+!qm
�YB�pߢ&"���AD�<��Bs��u�z$�9}v��ׅ���rhu�]����4�v��:�=r�x��7��=&V$�ʃ��˴QM�b���+��x���������������B"wI�UWJeR*��{����L��z��@��^8�Tj�V�:H�&���2�_�#�'�K�>�I�r/�i�V��	��=~�@�]/ ��&��2��R#t���u��l�i���u�e�F��r9C�����p�q��q���t��
����� ���Վx�6����l.�d�n�@ֵN�K�R�6�j����;�R�������Â� 2�8�&)��bN�	�x"0���vL�����˥�P��Qw�
���4��{�V���=yt�~�n�}�'n�e�M&ZN�_���˥���t	�X���w��h��
ř�@�]/ ?o�L�'�e`�{��=	N�Zn�V���y�Ʋh���[�u��77Z�nK��M���v�}�����-*Mҫ@�6`��t��X����Np�'z�5m+bhV$�{�w���=~�G�zs��I7@�W�hiպAn�HM����=Ͻ��.�����8ÈN.N�$. ŀ���ߺ몾�����k&����H���ڮr��%9��p�������
��Ƿ�5�S���RT&
դ��o�M�;�e`�{��=9� �W]JU�v��i�e\oX���w�Z�^1�F��FdSu���m�b�j�I����2�_�����o�M��®�\�)��;N�� ���ﺡDɚ�N��w�<�+ �X�����SaX�1���w��zl(P����.��������T��b�Zl�7�&��2�_����Z�m<A_{��*��ﰍ[J؝%wi&���X�����8`��t	��E�Wv&Z�'���݂���;�r�:��{vL�/[;�Um���CN��vZCn�_���Np�7�&��X�+�$�����jY�@�s��I7@�t��=~�G�O@��m���V�f�I7@�t��=~�G�}9� �����i1Yl�I����X�����8`~����n�� ���UsjK.�&�j� ������~�n�����UDfX�U1�@Kf9�X�&%��bS�!��FcU���`L�-I��&f��%H���4�UM]�Z�j��s�$mf�$��@9����lHf�
�C\�Q�[��IS�tF�+�{ur�q�����;�s���<�8��[\[����ۓ�3��;Y�Lt=�;��5åW[�5p��1�ܝo2sruk��Bt9���mx�%����:(Pt����$��E��ώyq���b�)���+��9M�7�=|F��v(b,j�+00���JP�I-���e˺5s�(�-���g�u����-��c��ם`���SaX�1���p�7�&��p�=~�G�O+��R�*M����M��:n�����tzӜ3�(�Jd�7d۩�*�MI5Uu}��z��G�}9� ߧM�=�un�[�I[l�=~�G�}9� ߤ��w�� ޝiZ�P���c�=��o�M�=��z��@����o�"��C�x����u]�G:���/��3u����t�prv+ztX9���I7@����z��@���wQE��b��n�M=�;�K���:�PQMЅ�~���#X�V��6c�)	 ��6@iK�MA�[�͚�
���{�߷�^��~�n�}��t�;ucm���z}�w�<���T)�����+vx��*���e�Vc�z�8`��t��_�������J�j�Պ�f�I7@�)/ ��������R�W��ݖ�v��whV�1n�;%�;^R�c�-���V\ڞwl����ub�I4�@�)/ �������$�r�#CN���$��x����E���I�yIx��J�GM��lU����^�I7K����"`�"D�YD1B�T�b!����"V(���@�0pH\
U, B�(IB�BK�̧�������L�&��軥2�����BS��w��g�z��@�]/ ���q;N�V�i����%��{��=K�7�&�ӿ8G�yּ��N��g��q�]��v�{+<ֱ�Ht�S��s��@Q�1q�9�]U�� ����y�9����I(���{<t�z���M�WD�r���E���v}�3 �.��}{��x�ܺ�*N�جVۼ~�7@�.��z��G�}K�$$�5m	�1U��{�g��O��}�X灊�!$�D%���h�����V�N�%iZw�z��G�}K�7��t�8`Ӯ�**m�v;rYrny��On�&�w�=�b�\koqgqI�K
;W7=�n{�?}~�}K�7��t��_���	��v��n�E��x�:n��R^�����^���*�v�����4���0_���E���t� ��]-Rv��4R��I��������:n�ޓ+ ����+�VЫ1�=Ӝ0�t��&V�������o�9�my���+������U�א��j���[-@�Sn��P:�k&�0�K����K&s�i�NԞJ�>��E�t6K�=����I�-�7m#��f7k�nzИSi�;z��F�cts��mv#Y��<���33�/Ӻ���g�[����V��c�%�'��n�{lU֊@��)O56��<�c����i&��(��R�����P.�{r'��#NA���?�~'w�VFypkֳ�=v��su�N�7nw㎜c��C˪����~��������c����!%��hN�,V%m��;�e`������oӦ��_GcN�����I�X��tz�8`��zL��i%Dt�*�V��z�8`��zL����=z�[���Vҫ�$��oӦ��2�_���Np�$���n���"�;��(V��4r#�۶6�f�����펴��;*m#�7����Umݶ*&�{�w���={��=9� ߧM�>���'n�e���i'X��c��D%�$��G��8�m��g���𒈈�7MVց|\�V�榗9�r�k�8~x��3��pO��}��b)v�'N�ZJ�f�N��I�+ ���@��0		,�[Bv�b�hm�'L����=Np�7��t	~�;c�Xv�qŬ���ɹ��b�(z��.�4tF���[�h�v���I�� ���@��0�t�N�X�:Ҵ�t�ݪ�y�@��0�s�@o ���ﺒ���joI������UUg �5�zx��ZbW$Kټ�� �)�5Ӵ0�z��nc�F����'%�ZM��k,�]K%�oFef���9͆�p�zI�tKk0,:6f4!|.8�u���FG`�7:(df"f���5��a�F�' ��k��� �B��BV��#�m�Z3��ܫI����ᢂ��ֺ-!�x
� z�	�",pG��W��� 
��W�D6�'��}0O@U�PzQ��h�6׷�zG�upU��e�j��i��{�V�]"�>��}����Z��Ռ��ZmZu�o�H��[8��}��|\TF�l��5D�#����N�ʜy��j
����r^D���̗�=$���AX�I�-�15�o	;���0��7@�t��7ˤZ����J��j�%i� ���t�L��)"�>��H{��[Bv�ݫV����2�|��@��ޝ7@���;`�B���Ӭ�)"�=9� ��>�;
D���~ɪ�j�T\�T�r��[8�BQ��~���\�RE�K�%�n�[iU���5tмsc�=��rjv��;.N�n3��^9��B���lƓJ�V�f�wM�;�� �.�h��{��m��V�M��;���J&O���t�zp����>�%���S��j�f�]"�=9� ���t�p�$%>���t�ղ�����}��z8`��-Y��E.Ҥ�ګIZl�>�t��8��n��[8$��g�And���0��g�|Y2|rl��n���m:@���x�t�mU,�.�z0�p%nMl��풫��%v=�v�[c8<��A���Ɂ�k����88�듷!:�_N��Iځ��v	��@��v�y��;�r��C��]=�Vk�N���N��6T��ѵչ�y5f�α��:[�Wa�'���dؙ��*��t����BCs��{���ޣ�v6��koT�xH:̛����)�9B�.�P����^7m]ew>ٍI:���t߼���]"�=9� �Ӧ��_Gcn��V�$�n�|�E�zs���M�;�K�>�֕������ǋ@���N��w���o�H��*�U�tƕ�P�$��wM�;�K�=�������(��m�ڰt�m��R^�H�	�����>�`;�)4;�m*tƇwa{�һJ8�������%�<��y1�l���Ź��n��U������t<�p�1��B���+vx���/�(We�Uw<�O@��w��*�H ����^r���yt�~��z+��\�MӶZ������w�c�@�Ss�TD�{-���zp��wSt]ͫ����������g�g���@��g ��zYS��m��Jƕ����y��Ӝ0�t����I\(��7Huv��n���C��^�&\�W�vr�y�x��;��(��B���S-��ne���oӦ��nu$�!����@���x�j�.��3UVp��}Q#�ݞ����@��g5BS'��
j�lSwJU�����/����ʻ����ub�R�!D����P���峀wُ����J��W7B������IO���t�zp������R�y� �5M��9|(�E�7��=Ӝ0����0����IB����f��sA2]��U%̖&��M�79�;�6�8l����=�qۛ=��s�䁮��iUUM]��=���|\�����Q�k�8�uN���w6�n�����ޓ+ ���@��~�7@��TX;Um�ڻI�X��tz�8`�I�zL�zu�j���*cV*ھr��[8~���3��p*">�J���=uJ��v��hM]���o�&��X��tzӜ0z�Ԡ%\Th�6��q��Gˮ�&wZe}�:���b#c8��u�ûp��i�fo��m�镀}~�G�}9� ߻��_��
��S��Zm[u�m���9Ix��7@�&Vҥ[�,�CN�'��=r����n�:L�o���W_�r�7N�j�E�� ߻�����;>�w�Ԣu�����;s7E��.�$������6���9t�}�7ĝ~%	�a(�)A��H�	��G]L�6�Kħl��V�8r-�t�-��W��i5laN7��n�Ӈ'[�v�Ixn,����m�v��ϭݜ��c.��nx붭pXc\f�Rj����cs�H�%���\�l��<��8�u�ܛ�rumy��!�z�Dvwb�2l`�L%�E`+e.˰6\�ӎx�zv���l�zۍJc��v�m�F�[�v�˲S��wb�ɼ�Y���!��s�Xƴ�9����y7oc���׍⛷��i&s[�[Wi[u�}}'��'.��o����e`t�J�պTƬU�=r�x�OI��m��z�s*�Sv�'e]�Ӽ�wM�'���6��=r�x�ҠU�M��WN�M��'���6��=r�x�}}. ��7HV�V�`~��9Ix�N�+ ��껨ҫ������sθ����n��jv���bݎ��������� Y����Cř�@����wM�'I��m��z+���v���Z��{��w���_S�+�U�GG]]jL�oӣ�')/ �zTL���Н�ot	�e`~��9Ix�}���ҹI��[Wi[u����r���:n�:L��iZ�:�J��KU���')/ �Ӧ��� {�4	�w�J]]�ݶ��n���I��������¾�=��sZXcc������7����uv�n��:n�:8`��2W�r[�ҠU�I�mUӤ�ot_u�>���K���M�=|pPl)�B��I��H�	}"ª���\Q�IE�>���7X�65o� �-[�U��ŠK���M�Ss�����[ݮ�k��٪�E�T�V6��>���%��t�@��?m����{�#Ǳ��J)���ȝ���	ѹJ=�c�ں��Ո�U�O��^���Z�����{��-_H��:n���Gr��I���I$���.�h�E�}��t	�K�>�֕�#�t��R�;��t8�p����RQ3�oL�]?���w2��7m���v��;���@x����Q���D �B���
"��ͮ���SsWe]ҕj���tp�>�{��%��zM�?���~q��]k�:��lg�3��v\��ohݶ8H��N�΍)F��N�s�"�<�۫�[m$�-\�`���I2�uu[�,�CV�Uo31h� ߽&�I��}��E����i7C)Z�Hv��>��n�$�X�/H�	rE�HzTL��텴$���H���W��O�%3������B�c���������V��V�`|��h� ��7ހ�|\���]Q�IG�HA)(�I����m`�&f���`X��!��KL�#��$!l��0t��B�*aK00�� ��.FBZ�K�`XR`aa��6�3gS!a v�X�l��j�S%�8�A��B0�QN�����f���X�NC$Ã���7f�٫f�ʈ���RҸ�b�1�8o�Ã$�LP��'���Y�wo��/� [@ H ��aR�ҵ�X��Kp�l����n.�7N�5uF5�A���Ԉi+v���Mn]�� �M�Z �i6���$�$:ޠ    �� ��0��J+5��8�8 �8��B�@CZ'@�   l,�q,�ͧ$�� )@m��-i��[WS�cb��#	�����N҃mul�l�o��O��H�dK�孢�������>��8	�� �î��8W�Ѽ��b%���Ix'�oYw$��)�kp���Lb"�(��˷a�BRR�<ck�v�B�6��X���z�Pb*�W�8���Os�%cu�RC���4T��5^�ђl��V�ܹ��nx�7`�0]��r��j�N3���wdk��&�i�����8LubTk�;n*޺��]��c���Cqؗ`�n]�L�&$M�6�q�r��l���!T����RQ��k���dd'�s��m��כ�tm���V��]��s�6�[و�4.���;9�O5y簻i';�sJnn���y9�����9@˂�vu��%�X��LlP� ���EɲR�p4�2�X����r%c7Fx`�d���ɇ6mꋦX�,c<nx��W\��Ĺ8�&����mppy���
�u:r�z�E2��a֢�m����cv���ɧ� ��u�9N��Q�m���\��*�WL\l�ur�L�YF�c�j1�k������Z��.�͇�e�^��͹�I���V�l�	�iV���B��ζ��SB��G5,ԩ�E�&��Aڪ�Zŝ"�t�<v�*�d�`�v��� ��
��Dׄ��eYa�'vcP�Ά��$hVsv�(�{	�n-����3�l�Y����n^[���Mu�m֖��n�9����;�1$��ul��w/�;1�B������s����7/lpFų���x�{d��JI�ۓ;��#���4������d�����O����`@ڋ*t'�P=D6
��*�(�*'U�ޙf]c���N5뤐! �2�п|��L�[2RM�75jJOg�]����u��ӻg^�j�u��8�\!��������Lsv���=��]��<a�mq״���vT�gv����p�z��!{e-K�rm�X}j��|֤q�ݳ�E��@�3[-t�6�@`w4�@r��=]9���|�`��1�.�v9�#�v�a�˺y�"���L9H�j���P���L9�ȶ݁��,�Y7;;<qڷk�+��I��q��)h2��������<��c����,~���I&V�����w2��7m����w�}���I2��^�h�� ��n�bmUӤ�7�t�X��"�=#�����K�*C���B��M��/H�H�}��n��&V�]V��2�v��W|�9]�p�{���x���E�{��E+W���cB�Wm���,�.s.�ޡ݇��=�WN�s{c����Y�ʴ�I]�h�۠N�+ ߔ�B�K�{zp�۲n�������ot	�e`��:8`��7�U\��ݞM��]�sUUSv���}�p�>��n�:L��u�j���ue;�Z�ǠN���M�'I��m��=�.�eZCvӶ���ـ}�t�t�X��#�'G��҉�l�竪�l��+��A�wn�ssd瀜g���k�#��v�kv�*x�k���~~���7��Z��}�����'c��![m&� ��H�	�� ��Ͻ�|\ԔDɚ��k@�rh�E�W������8��}���J9+�!(A�`:bGLhtڒb(�0�%B@s~��U�}�o�	��\����i$��l�>�t�t�X�zG�N��N��m	�:�EQSwހ�.��!}O7o�5�������N-��H����f��ր����כ��V6�Z�ŕo��ͷu��؂ƕ�m��ޑ�����M�'I��N�iZ�lue+�Z�ǠN�{�7@�&V�=#�=���U�7m;iYhm�{�7@�&V�=#�'GzqEZ�M&���!�}������<v���%��Ĕ�������򡯽��h�J'c��![m&� ۓ��'G��7@�&V���Ab�gAMn�H"<y��jUFz{�/]�u]g���olSLEբ�^�`2�n����c�'G��7@�&V�$�@'_�r�n����V+l�;������6�����mI��j���Wm��.�m��!B��[��o{�>��v�bV��Xܒ=r�����2�	ӭ+U-�n��t�R�z�%���t	�e`�x��+_�|L��[��R�b0�P3�Q�<s�-Utj�'Y�5Lt�d��`��R�>���@�j7M�<r��B�
��Xqq�X84��dE�ta>]��q�9K��S�f1ٸ��N#Q=<��	h�gj{΄$�n��sGud�k�Zڑ�v��)]Y��}����� ��ێz�r\ɺG��sm��F�ݹ�{n[���8ݹ
ke��P��f�y����M��t�r�چC����'S�`���쥫g=t\��7�	�vn\�1uRMw=����|\��u�D$���vx��5�U�M�,(���@x�6!L�mn�tu�<31��ƪ
��e7HM7i��6)"�')/ �N�+ �WU��̴[��Vr��Ss�33z����O�{�] �1��UvT�jjJ������a(��w��}����Ss�rb$�4[zJ��I�̜bwi�,<g���ݷ��:�^6�7��ݛ�	ti��_���X�:-yIxw�n���Tq�nB�Q�q�d�|�*��P��DD�.���8>Ss�;�����֕����wt����-z8`��ޚ���n������,`��U]�����6�{�7@���zE��%;��8۬B��&軋�Quwހ�� �	o�7k�76����ށ���붘�s:8��z�p	������s��}��5��a�ǘ�y4�g����f���O��Z�p�'��t	˥���� �-N�+����	��}=�t	˥���@'��շCV+Wv+�8����V9�Ԣ(�B��H!� �Z�Z���_w8`��Q���1�۱*V���K�;�:-z8`��߽Q�v�b�%�EU]� ϩ㮁�!(��i�3q�z��<TB��������Qh���xl�N�[qѻ����ܮ�7��=���Q�#,�(DɌD�L����'�'�O�t�r�x|��@���T�m�v�U��X�t�r�x|��@��+ �HQID[C�Н��@��^�)"�'���=;���/�V�YMի���n��I�=&V��7C�
�N�8p5�s��ɩ�ժ�x�-zL�Ӻn�;�0�I���?����5x4ɉ���ݼ�)����Vώ��m5�nzx�ۀ�&k�.��X�t�w8`�-zL�k�Tl��1�ڱ*V���� ��%��e`;��~�wm6R��l�:y�z��XN��p�;�u���j��+E����OI��tN�����}R1P�NӶ��Ӭ�t�w8`<�����$���Z\>��q��-Fb�c�����zGV�X��$�Z:����H�d�Y� �n�˫���!��Y�	%��@DY.t[o]�Sp��x�&��n�:��a{7��9��G���\�#Vq�^;'bu�T�r� ��=�����:ݫ�pv[��nZ�V�O	͘3��맀�N�÷\i�-�;q�h;�<���\f`8�Hq{{ArSz�w��w���NuU4��B�G�X���������g�"��=�����F��ݹՅ�
I��e]Zv������:y�z��XN��Uի�1Ю�n�f��K�'���:wM�'u���(��55/��\�ԫV�T�/��77x�<�ހ� ��nz �1��7C+Wv+N���t	�2��r^�=&V���*���P�+ot	�2��r^�=&VӺn����v��M�"0��!؜�h��uҽ�^�n@��ܻXy������y;�Z��s�]h9� ﻲ�w�0��+ ��ɠ~b6A�Q^�^$��}b� PH�I&V'���}R1P�NӷJ�:�$N镀I�%���p�T蛢��	����CTB��[ޮ���t���~�ހ{%��Ւ��]�7m��$�d4	�2�	=�t	�2�	Į���*�����C΁:�/(5���8룮�1-�Ocs\H�<���Z� Y����]��a�OI��IN�+ �ݐ�%����t�Yt�:�$���N�+ ��!�N�+ ���Q���1Yh�i�:L�}����A�|w�~��q�Rq;���s�nw���[�]{�n�XU��n0�9�Ųo9��w�{2��yC(U��UU<��2��K(:�6��BLŃ0�,)�(�t�]uѥf�m�H2�6`�F
�q$Ԗ:�w���L�Y���#feS�aCj��;Kqu��!���$ڗ��耍NEtɭS�f�HA�p.�ծa�p1d�w(�	\�
jDѰ�Ŝ5���!�an3��eX���dDv�$��Zw�}��gǥ;#A(BH]s�Z��\��f��Z�[�o�rj�0���3[&'j�w�&�AN�n�#sV���b٬v6�;m"�sz�"!��(i^�y� Ȇ��T^��<؂� ��]�~�b�;��{Ĝ�>�'(!�	[u�Iݐ�=$��$���wI��t��]\UmP�E]��@��+ ��n��+ ��K�;�ﮔ�.�)۴]��^�k��Wqn`9�w�x2�h���p�;����6��1�n��n�m�=&��2�	9���&V��(��e���@�I��Iϥ��2�	=&��®�Y)����n�	9���&V'���&V+����2�T�u`�2�t�X��t�=���G`2��%4UB,�J$�C� �
�8UP�T(r_|�I�u�6��:V��[f'���&V'>��{��~Jjz�
����\�UAuv���O���YN��i�{b��������z��ĨJ����t����$���tl�	%����@�bw��V��%Ъi7X��^����tt�Y�Wc�6h�;Jn�r��S=�O@Ƿ� �Λ�{���;������Zv[i��M� �N��{���;���0��Wm+l(I�ott�X~�s�=����>�	�����U�"N�s���Ό'F�{A�V�;�t���pl��b@�$`���G]6Cm��Ӛ�S�-��nA�Onzً�Z-t۳���g:k!������ٞA웞D�����e���+�f�.$����[���5�̽!Cc����:��c3s���s�su�vlu��9ym�hGJ�
���GVF.�-�V�mb3�]��[�mm��]�ӷ�s5&;F�؝��&s3ε�n[��m�&Pn9Q���m��G+e�-C�7`a��xѭ�	���,ګ����[���l��z��. זg
�ĭ�V����{��'�n��+ �ϥ�ʸ����B��m����L�O>��{���{��e��ĨJ����L�O>��{��'�n��x9��黺�h��L�$��z�8`{���ၿ�������E����3��&�g V��u��r5�ɺ�-��u��(j8��jUU
g����l��z��?B���[������*��&��U]���{�]m� ����H$hJHF�(P�(JT(��������c�`�
)(��V��v���0	<�^�������VJcE�'m�`y���0	=�ttp�%z��X
�1]Щ�<̽�0	=�ttp�$��z�����w�F����8y������NI��m�����xsd#����ۯX�Hv����m��{�=����㞁�v����+-��P�+ottp�$��z�8`'M�>�8;7wWm�I�3���c�p�T  	H$)"!�b!�b*	��
�v!DB�<��z�[8��4]�Rj�t�*�s/@�G�:n����B���1=yJ�������M� �N��{���wy�z�8`op$/��H�2ĂI%��j@�ӄ�wof;6�K�g���6�����ݹ�ۖB3u�ݴ���%��r^���t��Uի%1�Ɠ�m���%��~JJdǷ� ����e7<��9Y�+�:�/@�G�:n��R^��%�ʸ���0n�
�E�p�o��M� �c�:� �"�����`�!�!$&ae(�Y	���VP���iS�߿~ﻕxO\�����P�$�@�)/ �t�h��}:M��KX����RY���n�m��@u`��S�L��E�ˢwKۉ���`�������IZw�w�d4tp�>�&��%��KE��V�2�E��0�I��Ix{�C@�Q1RI�m�t]&ـ}:M�=�K�;�2�8`{�E%ے�\suWކ�Q��g�<{�:��`N�t\!WV��ƋNݷx{�mh��l�7@�)/ �����o�9]��\��]%t���Kn�rG��lppZ��Z#�M�U'g�iS��l�����ƾ۰f�t@>��t�'mv�F1x�� ������ɛƉ��;s�t�>��t��2;�0�V���x[�8s���]Z>wO6�v��ϴ+�v�҆���砭��+�te���y�f3�FǌHA�=�8���á���stu켺mܖY�E��qf�ݭ�_ ��k���`O���t��t�ʞ(�U5ݮ^ۺs�H�7Q��:����'x�a�o��3�������gI��Ix{�mhʸ�.�CWuv�ـl�7@�G�{�ց�+ �t���]�b�*����}��mh�2����x�����#���!��6O�
w��=�8~�}��l��d�*b��C)$+I�h��o�&���}�t��wR���M*�m�m�97k]u�^v�۰�wn5�˓�e�e���vI����n T�e�v�I�`�I��8`}�6�tp�7��IEv���@ڶ������ڪ��M�>鵠zs�����z�
��d�4[�����}wG�{������{����z�L�
��(��ڮr���j�����i�>����+ ���@�U�Ahv*"좮��y����{�]������0U�t�����c
�����*j�fN��k����Z�=���k�^C���;��^�����w���>����=�� �w��NV�_(�"��ېY'wG�{������{���;�֋���t2�B��=�0���;�~�U$ӱ��>�}p�]�~�������I'wi����0����&V�������)(��[j��M��=�e`�wL�=�� �zM�����_�v�Lq��B��\oA��gN7\��Oq���[�6�/�Z��8�uᐴ�U�۬ ����ό}�7@�I��z�S�݂�.�U�̶ށ���n��+ ��믎]v�.��v!6`�I��L�{�0�όWK�Uۦ�/�B��@�I��o���w���g�D	�&�+51^����Ȱv���+[s0��m��֡��ktj��� ��(�w�����E�00�"���n��p�>�>0����0��J� ��ۦ+E�B�2ޔ�]����y���97��ùޙ�h�hqœ]l��]��8`�I��8`��{�u��N�&�
m3 �zM݄�S&=�8�ޜ�e�ƔB��O�@���۫v7V������0�p�>�>0����\T��J��m$ꮬ�̶p��� ��z�'�L���?�.̻t
��3@�GuDGٛ���Ձ�z�������_Є�  3�   �7�(�+�K����0ب;�D@�DP7��� �9
�*�*�/R�����?�Z�B(
�*������w��{�������?���o_��6>���_���������������4�  ��?���?����   :APA����z��)�������?���    ���?p����%� ?����?�?n���?�h��G�k8��� ڈ���T �Q&JP ��Q �I@H`$���� %d	BEa!X$ d$	H�����  %��!	B !BA  @�$ BY`!$I		�$ ��BE��dBQ�!@%P��d	RB�%BQ��d	P�%BT$	��Xa	$!P$	B B `!@�IQ$	B� YBQ� I	�@!	@�!P�BBI@� � @ 	Ae	d	Td	$T!	�!P�%�%D�$� A� PaU	XB@BDBd� Q�YPd	 !	 A%E$	Qa@I@�P�e@$@aQ!�$�	B` % 	PeQ`	D`YE`BUA�U� YFE$ED��2C PdE�A�a@!	DXFYE	FDHFdQ$E YdTa	$ aP%E�aB�Y!�`XFE�eIF�`F@�`I�dHF��e YA��ae �da�f!�`�d�bP"Q�E��	�b"� �fP&E G?����S��  ?����=���N��<�?��   ��y������������  �*?������g��  ~�h  ������   ���xm@  <?ㆿ���c[:3�k��g�7~ލ�@  ��_������  ����?����|������1   ?����   ��p�d��p$|�?��W����̆�w�   ��������Z����ߏ�@  �7g�y�   ���������/�?���?������
�2��C�/��:�����9�>��| �@�(�@ ��4 ��U ��N�T9   �   x �Q@�   � @U	�
J��U���J�*%�P @���EB����z��T�   C    d� ��[�ԦM}7�[�)�� �O��O}�zoz�/[�����C��)b�Z\X� ��Wm�����z z��[�j�W�^YU[��: ���y��x��94��6T�� ||���@� �n: ���&�  }0 ��  h�`�@ g@� [  {    f �0  #@ m`1  "(  @� 6` 	�
$ �M  �@@*� ( L V( ����}�uu���ݞ} b9��uy�{�v�;����j��{�m\ �]95֜�x  �szW�ǹ�{� 3�{�ꥋU,f����V} �z�'���ݼZ�>�����]� �� )@P �@>�����\���]�νw�+�ǃ�-��R����������֝�zU� :U�����׀�{�7���y����,}޽O�֜��.,�� YK޽/z�'N�x�� �      d}{��ũL�|�����'�0 б޼�,��^O*�d�>��ܩml���� ��,�/y��� ���{�O�^^��5�rt�� ��O[�n�ɯ�����ד�M�    OQ4m)JH�  ���2�U=@#@O��I�S &F "{RG���  S�	)J�  D�5%"� x��Wߋ��J?�������SP��~��Q	D+�]��U]"����_�_�TPUb(����^���ĸ�����?��SӰ��X��Q�B.�ԅ`�"CA��Ӻ��R�|���f�q�[Z�>}�E(�G���-ti%0���7������#�	��#B�rI3oq
A��R�$�x|37�X��p���f������K����sEMN&�HH��s�8��^K#���r^y��~�H��k|6zp��k|%����\#���,���)�'W��q"(J�$	!��`�Ԧo�s<�Fxa��)e��[��54x���"H4��_���H�: �#�@$`H�� P�g������>փ߷�R�g�Ъ9�)|�O��H�.�)e�n���_dd������#�pI %XC	Ձ�i�Mi�Lcr!\̗C$$6�eBr��B�5���p=�O
羞�!d8I@���kA{!��{�^yw�4jm�ae�Ò$��썚6�L�/��E_tՕ�R�Թ��p�k!a3Q,�
�$ $u(��7�5�.���pt�$��ċ��Fd���s	�|���]��r1��������3 y�X�9�M�-ќuM�����44$�$,b�[��N>��'��T�+��ܸ��E���J�W9J�ԣ�Q>�����>�k�K��ea�N Y)R����u.�u��B����'�<߳�!�
W`l!H���B,v���Sp֡|8B���]<��\8{�$q����`@�l��ݼ=0��kg54�!.�ߔ���*�)x��|�7! ��Y~6I4�K�5��`l��Ĳ9����Swt�-z�e��x���GW1yzѫ��r�W�tB�LŒY��7�7�<#~�v���_ГC���������$<���F��+�`D���
AbD��#�<�U.(�B��5�?:P�&�^]l�
j�j�A��qb�]B��)���<�K9 ]�T�*]��^�i<��Tٕ�A����$`�	d�4�ֆ�K&�D!
d5�2HC&#��D�D,"Dg��<)�"FH�! h��p�@<b��2
Vs�W�ؕ8���$*`F�dhd$!��0��M����H�#� �C����!CÎ���aK���'8g��e޸�U�,,`� HR�r��7_}��e6( ��i H�$R51`W&���O3|�h��� �H�r-I W�|YxS�Je��s��ԊP$��5�5&�L�5�����dE�w��r�1��x���1����ֵf�|~����f�V4�&�]$�6���Ħ��W*��Օ2��_���}�2R��U
T�ugL����R�U)��w��'{�*R�ʑ4�R��\aV��V^�^M�r���r�}4M�
���� D��8��a!�B/�;.�f���aH��tH���D�M��Mb`Rr��������J��;Ve:�/���} ?
�5����s�י���:Hߵ�7~8�$�� �E�$�T�	\�P�9�T�Du"6p�fxG�o� <�b��F' ��:6�3�͒'�g����!��o���BA�}_6D���{9O9�"�
��՜#	�#��G)x�Å�w��Ӑ�C� 6X\�0��1�D
��Ǟ\4,F��ɢ�4J9)�o~��	�F�v�W�y��a��ˣ͞�!�ě�I��<!�s�H\7�p���8x�榳����y7�<4�sWz�.�=5ˣ�c�4�6!��ﺗ�!0�d&osP��Ɇ�Hy�B�y%ד�����)T�[W��I���}wv���R���n�W,�K�R;Vr���>���ߜ��z���F0�LtiѱH@#V�7���k�	�|Y 404@�y���8��p P1�G.�}��7�y�u�霺9��<��.44�M&��}�p�oz�;�I7���'�|�/U�[{^��\/ Qò��Pʋ;1U#��1���/)��y_0���j�z�msīHR�k�k��3�F�QHP�#F��*b, �Wq�B�٭߮�O��5�N�������� �����j��vŐ��R��NO\�2<�0R���p�4~X4�n�>�ѿo���Ҹ����
iqw�SĹ %*�8��� ���2B �2$��G�}������!33���吅|AH� ��H�I>�C�`�-��du
b�	��8�˲w$���(Hm_7揦�[���<�L���g|i�h��-L#HL�@��Ԅ�@���:�|�����]���_N*q�p"X�GP�Ĩ`�FHJg9�j�˜��<��� ��,,�H���t�=�$dVB|���G���2�	o�����kG$�f��Jx��B��>&����sz��߽9��\��ĉ|�K�Jb�.W<���%vzU��i�6��P����^�~�.�l�8�ry��<���2�۬W��
S����L��]Q�8�>��Y�QJ�C�u�`�Z�p��Nv�"��T��X���7;eb��.)\��]�����8G*yIWV�HI��5 ��F;&0l��p�����S�VBA�1)	r�Wmt�1I_o��.{H���x�&0��K����nA"�Wܛ�s�I�1e��_<�o�������޼+W�����罋6�v{�_���w¬��Ͻ��W�i�>M���#H��Л� ��̑$����<��"Qpf'��}�a1dO^,0N'�'d `�5�"I'�p����<_vJ�2]o\+�Zz&k*�s=��k�È�B��b#�����Ȕ�b�<�W�xz�^Ϊ�v�k��^�}��B��^�HR��c.�e�t�aL�.��|�
�HY�0�P�5w540��J������!p�|�Kœ���y禮1�0цl��t��ᡣ�4b
᧞��v�����ˮ�]�[�{Ҳ��'�C˴s��	�J�1��t�����g�����y��ׄfkfk��>H�55�5����[+�������|���ɭ�*#��H�8I�}�Z������D�� �,B�sf{�x��a�j`�t�as{�%�<���ƏuN� W
i��`�1bc�y��y5��0Ü�uA1Q~���'��O�����}M"��fyyp��9Kx_n�O�����)�l
j�7�w�a��>|�H\4;����! X0M"��8���:��0��tŮ5��M>�?
a�|���񭌮7�e�t�|1�:7�/����h�
a���N]����<<���b\]D�#�1(F*$Jh�NWA�SZ܁E�I���#���P�I1P��:H	@�J��̮� �#��O)RXYe��(�Z��mӿK�^8���"0!�Ssg���ּ	����о�crn�|0vE"��
�i
8��hF�6H3,@�H�,xs3F�����'��u���|���i�5"K����	����ъk������/��O'�9���}�_Ff__��݆	 �IG�=3�i�Gr$��@�2D���\!���>c�Fkxj����$��"���EqLJ�ޥ��Ԅ!8Qi7J�;i�*�T�ML�*+�p��|�|t� dߜ�%����$$��P���K!	�Ⱦ�a.�Oy$|��NrM�|D�� �d�a,_b��A�`c��߁��9�O�k,�z����Ԥ��Ƙ_\�5]��{xFN\4F�4���w,�!!
�泓D�X��!=6�|����,!H��!�c�$!0����Cn�$B�XS��Oe�)���ڑ���i��RH��}׹�8��R\��{�� GJR���q�t�LKo�᳙}%��%�_p��.D"$_!!w�y�֙�	M��g���ka��F%"X!D��$5�]8W,�A�N@�p�3.�̰���͓y��
��S�y��"HH��E<��A�����a�4��Q��4l�3z)�,8�`±�c"{!�m�`�@�2��0%�I#Mi��nA�2�(B�
{d8@�3ɶ��ar��$��
�)"H1B��@�C5�kɔ�7�f:����g{����4�m���4J��ѭ>H��˚���N0��.0�2I�&;�/	Hf��V@�!d�S!bd�/'$`�/#/"]��`P�t�c$J��Y�}6  �m4P I#j�m�?`�m��         �	            h�         �`    �`  p                          iJd�sPm�v�kX6�m�� 6�j�t�iVBA������m�$�m�   	 H�5�� ��	  ��#� 8   �h��� �[p ��i����md����KuK��]@R��z�3l��u��	 [Z�P� �`$|}o�k�m� 5�ګ�� O ��UQ��P��-A�l  �i1��m�[m���j�$���m�,�    ���m�6ض�۱ �iZ��-� &�_]���r ��� *�UR�Uԇ\��1�m؝��[�['3�$��,k֒q�l 8	v��mpm�l��&�  `ݱ!f`�@ �    �� 8    6�PH  �6��  �Z�M��}wπ��        	                           @  �>     �         p         ?h|    m���     [@�    �               � -� 6�     $                             6�    �   H   6��o 	ՁfC�f����cC:�U$�q%�$u�[� �[@ �j�қHY�z�]� �  6,���1�Y`�M�U�R��+l�
���|�R��-l��PxK�%uz.�ŕ��Lb��~|� 9�Z��r�� U7j�j�r�@Q�]Qm����I{iV�H����v��S�Ω����`�# �%ڻXQ�UW��n��d�^�vzF�'����=�j�(Rb㮡�d���@C��� �)�W2��λ8P��e�[���w`6j�2յ�k&�)uT��V�*�#Ɓ�S%U;0mHR�����ڪ�k�c0���ԸgWVwd����6>?>]����m�ʎ�ǣv쐚�K����7N��@M�켆����U�w*�)Bs�-�=٬:�� �۵,���y����i gsq�;�Sl�yp 9ǉc$#u�oZ��#!%(9ô9���6:iy��mg6� -6R�%m���ڰ�[�Pᳶ]�mz� �[p�������"e  m�m��i6���|���QT�ppƱ` ��( kn�-:�n�#*�U�@R��Q�ѶĆ�\�` [D���^Lf�vt�д��> 6�5�&���6��	����]��r�U ���U*����5Q���@[@�[k���h 6ͱa��8�kZŴl -�i��a��a���W���<��.L�UUl H�� ��)��-��pm�f� F�s�A�my�mNn��kn�  �� 5���nE��#P�m3�UPqN�XZ��e��VU�1Wn��\��g\Ny�PM�U�K��lJ���YE�\h�a�I�����ҧM�h�q�A����� �s��tA�@�uhkۮ428Zi���H���%@N�v��Q�0Ƚ+���T�l��ٻv-÷2���ݫ�b��f�9�����v9���鰝6��[n�
�"�Q�+T]�{��ú�Z�mU�����Ͷv� ���`�N�dv� 8 6ӳ&�6�B>����)DM����     �B�	�Z��
BR�[zt���� 6�e�K�[G }�Yo�z�mK��h�Wm:i��KjD�"n���jUUj��l���@PP � 5�  ֛��Ԡ���l�      �6H� m� �l�������m�P#	��%*U��nV����MT�ֶ�    m��b�qHi��W%�@��jN`�` �l K�j��X]�R�ny�eeJ*U�D %^B���ջo�A6���%��	]Wd�y��Z����S���'$a(z���Yr��[*z�T�v�3M��$�f�f'D����5Q�Y�5�
x��` Ii���6$q#�� 6�&�$�-�ܽ�2-�ȑ�m���I&H��ݖہpMj��0�����O`mu�e�����ͷ	�`Bt걷[��ӕ:�vʭi� �����X -�#'@�U�tH�E ���N�2Mְ ��,�S�Sga���-���ygF'*�3KMζ��km��l�!"�M�l ��Y!�l�ݬ��lR��@j�*������O<ܭG	̵�)��kԪ�5 UuR�m���P/[��fZ�Sm��{s�u[@�&� <?}��v���9,�˧Ip m�O#]��r�[UJKZ�-ݻH�VŤ��4Pv��ZǢ�I �bh������D�+U@�l ��	$%�m�K�i3P7$�+Z��n÷jX
�pXci)M�m���e,�94���-4R�g'NJ��*k\{Jd�m�u�>w�q�c�gg��i�W[t�v���U�u�"�T~>@|�����F�pk:5�P�z��6݅�(J�UWT��宊�ڱ#-֣L&����d������$݇6ض�/�ζ�7����vЂ�����jP&a᧗n ��9�L�Q�l ^�Q��v�6�,b����&uAtv�j�W���sʎ�'�:����R����E��UW�yͫv$:R�"�(�����Uʻ*�V�Gݮ�
�Cm۶��R��UM����s�$�f�t����h8��%[cu*�Pkn�A�[P֬C��`8�)%�m�Z�Y)�b� 6�i���-r%� UR�&7-`�f�e � $��`n�p��  �6��N��  �Κ��m�3N���	'M�a�[�	6�ocn��kmm��wv]�k�Y��}��I�   kn�j��*�J�T�!J��=jRB��@�d`�n�\�J**Ռ|��ў��UT��Քj9�)����[�m&�m6�A�l�t��-�  �[�3n�M�m�k��ni�؋h�I��`  $_�6ػr�9�kX[N�̒I4��j T���.���ŵ*�l�^�̘�+A�
����.Y�j�a���&�=h�`:3�ձs��A;)�c��[z�6�a=2ܭS��I��J3�K��I��U�I�nL�L�ݚ.�[ݳ�ppP�<T�5��(,��»pP�eR���#� �m�ѻl6�e���a�it��b �I�\KT���hh���`�`�% �I3�m�mЄ��,#���F�V��4�I^x"��2�!6
.�@� [Nn�& �Vp�\���XSAƨM�6�KMrSrާ6��J�	 ����t�Œ� $#j��a[lm�2�E� 8[f���sp�U�P j�:UWj�j�&ڶ��khX�	Ö���ݎ:��b�  -� 7m��h�C^d�U�TԻ6� !�e�� h �`rJ��mn��nٶi$���   n����� ֲ�*�)%�z�7bZ�Àl�vl���nZš�vm��@ m�6ͲCܒٱ6�n���&��a� $�XHld��U"@���J��.�i��I�[@ n�	��n-��Ԁ  �Ž��l��{:�V���h,H�T�6��H�:rZ dt��۔�FŶ@mI@��,mP���U� 5@ �@ l׮�-��OY��-� P'1r��ԫl��V�U�(�W��)�&5�WY/��[�/���$����iP�e���U���A�����W����(�F@j�W���Q�#��;-Ӵ�UʛPt�XAtGQV6����ui�[Gh��6�����Vv@]UUUX�u�һ 5J�@ؚ�����F�����S4@�������Ʈ�s!f;!�kT�0���0w�[K^ͮ͏h\O;e9P{v��G��Z��&ճU�K]��<I�T����P� ��wiZl�UIӊ�%Nғ!�:��F��y%Έ���[u]�cq,���o+ Ӏ��gX쩧|��|���DD��U��q�U�0WR�ɴ��+���0�ҭT�H*�5��չ@-��1�j^y���;n80�Wey�jƽk:�[s���8-�-�Q��|V4�ͼ⛧g\���n�T���O	��ڃ�c�8�H�]�^���cm� J�[|�
�U/7(��P��R���&x��,UCY��e�0d���t	F���:��t��HB&P�����8j�%���Fѥ�fA��8T����K<�۷[G4�2��Wno���}\t����j���/`��ڕ��F�pȋ���;�S�):_e�ki�i���EM�ԚԺ�u��ֿҀ�*���@8�����
��D�B�D8 �x*EW�h��P�'AH'O�.A�&�4"�a$ H,�aċ #B IB@""1�X�"F!�BBH��@� E D�A���x���A��#G��z��!��D��Qz,HH�� EH��	@ ��DȒB$"X	@H�@ddQ�p@6(x A=JA@B�|���Q� �	U��)D��C��� /(z��=PP0E<�"B)UD6	����B�"*�P"Q*A�D���O�a�=�#Ev
���  B*�"���b�0h"����@�H !��/��>���C�T� # ���4�TC
&	��J�D�G�E�P�%���� �:AZ? �h]"�P�t+�������A �� ��;��w���m��#���� �[p@  l G릹fד�����d0mԪ�;��tYy�ɶM�m�i靝��-)��N�l�6)UInW�P��;�90:sjeB�s�smf6Ɗ	�T�� l�  ��l	 m ���p   ��@m�     �`���HIz.�N&��M�/=$�Mm�Q��+���ܹ���u+����]r��Q膷v�[�X��	vsų�!	vn��-�tI�۴�6}v��ż���c�H�XD6M��B��Ĭ�2�H<���n�W��`M��B�q��s��� �a*�S�D�3k��Ʀ��U	�l��	�Kr�v��u�b��������Eð���c���V�д�k��/Z�t;��9�r�)XRT�IYQ�K��Ν��i�m��������v9��IS�xA��'���%kV�T�v��X@!Z�O�89�6�mr�aݐ�|�u���Y�ұ��i]�*�6���aSX�U�.6����8���=t)�&US=	t�m�����&l����Ş8�;tnv걷�X��ݓ�܍�Wm�+l����)`����)��]Z������l�C֮<��]�_
�͒�5���خ9�0�2:`�'�FE��V��t:���մ��kQ,�_thG���ВB6�d��;0�rv��m=����P6�i�ݐ�a��3��%�"�aؒ�^=�[W���9�unŐ�3�P��7��m�t�pr�M��EW����VAI�u6w���oE-@\��TKK�M{v��'��H0�t&���Xv3!=��kD.�V�#�/h.
m]��;lN1x<�m�2utb��m\`�8�8{f��ǐk���E�=�=s�ȱ�Gj:le�3un&�I�V\��[O,���ǶۘgC�KL-�H[Ca6��W\E:��.�m�T��x�LԘk=���@�@S�>���)�����6��ݾ��WK��5�:��S�^�<QGR.�tRYZ�&���	 e���Ӫ]Ht��ӫrf'&$wd�+�0���n<��g&�mE�l[�a�$3�꧳ʧ`���Q�k�[r�;+g{=`��'�pN�"��2�rL[�8�,rRM�6�ݓ�����)Ǎ������9:u͢�힊�Ž�S/F`�tc�p����{��o{���<��6�6@��x�g��S	�<�v|�p/	۞9SC��g�w�c��Q��5sV-c�Tr��d�P|H|R�$��]�v.����k�1nk�8�ǴQ�%C��$v.��W9XQ��5s��N~�O��"�Q��#�8���{�,.�Va����MQ��A��jG`��W9XM��M��5��{�^��I�M�v�n�'M�v��ӬS��,�}�g��;xN�"�kK���U����D�+ �ܬ ���x���6�q��Y��*�����jnV Nr�M����z�(��R*��Y��{�,�����K�w����<�Gp��4�(�D��'9x��`6J�57+ $�7GąR�nK�3]���Z�,�v�͖wbn�o�D�I��]n�pht�Uvj�����, �7���@��t]ct��(D�%D��$���ܭvf� ����3]���J�$�9QF(�j�u�jnV lr�M����X�"j���rF��9�����u`�%��&g؝X��Vo�4STH46�G$���W˯w���{^Vf� ������D�q�.�����X���57+ h���~��H%)��������M�H�����Wn����G7P�=s�[�(�]����X���57+ }O�`�᭺i&�Q��'�sse��ܬ�?E�jnV H2z����%)��8�5�ו��W�Iun��}�����QĨ�H��3������:��ñ�	��BK3]���J�$�9QF(���&�`�/ �ܬ�?E�4�E^�$ݴ�!���O�k�$8x��V�>%��"ж<�>���Y��ڠ��g��lr�M��S�X��`K�EB��A��*9%�ř��μ�Vf� ������D�q�#�S�X��`�/ �ܬ:N:��B28��QXY����,,�vu�j�5�ZcI6R��AW*�:���Ԓ�S{]�5�`vs|�~w����>�+$��fځ���Z���7L�^\���*�*�+n� �R�UR8u��q���z¹9��עn�\	��?�M�>p��ڢ�8��*���f�;m�9�ح��u��/d���Εʃm��"x�k\5��`������G��b.�<��A�h)1v�ud���`�I�]��l�ۻ����N���O��x�i�bWq�=��"us;��׽�Q�.��6+���L��G5�Ѫy�l����]�
�w\6�,i,�ǳ{`�j��R~��?E�j�+ 69x�q�(���@�;r������:�|���K�����v�l�HƢ��Q�]�v�͖s]���Z��F��TR8�Q�#�k��j�+ k��`���$�J����A���s]���Z�.� ����������	�#Q7HΝ�7�q�I�&���eڗ����Y���S�vm*�D�q�#�1w+]����`��`qw5��f���B8�U#���r��ٰ<��"�T���H��J+��g�����'V װm�bMH�7�sse����`b�V�����7L6���N�Jm�0\�`s��W9X���5Dޔ!�E8D�q�������u�����K����̠��[N9�qH(9��<m�������sN�4�L�Y���HV�\�u ��R�`�#N��8���c��j�+ k��`Ѕg�G�j��]U]� Nr�\�`s��W=v�Ƙ�B� �܂�K�3]��؝Y��	DEW��� �=�x3MT%$��`�G`j�V��3]�ose�ř���k5ԧLrD��R��X��`�/ �ܬ.~��~������`���<��q�� rOl�;�5ԽYzW[ۖ�z��t�qi^v^�(oYUu���Sr���W�{Pr��x���%�p>�ے����`j��X��`�/ ��xE+��/U�+��	���M��	�^����[�:�#���������`��`vsXTB!BUR�����3G6TD�9m��{�,,�v9�^��XȾ^��U��JҮ�����u��8c\�m�#X�=z��c�����4�DE)���XY��{������`��`�U	I"t�;����	���M��	�^��XcY��:c�&G7RXǚ�y��57+ '?K�	E���B��T�&�R�P�w�����`؟,=_}����x���%�p>�ے��ܬ ��/ �N, �����J�����uO\�h!u=����k�#i��z˭D���U�����qɹѦ��:�/N�ү9��<�emf���d��-[������h9�pݶ]��f��ī`i���pNS����ڹr�G�������*�;Kbְ�8�'t��Ի���ت4I��5��ώyl��;m�9W�Aj8�ў�vu����'o[['h��Sr�u�C�F�kV�p��E�&`!���.�֗�m�{u�����Ge��x=w�G���|�.g�
�j[�-�mۗ��8z��v�����׀k� Nr�M��7��z�"�*FE �u%��y���W�I�},��;z�X�4wLj�$RHF�� '9x�%`��,�8�	%���)���XY���CU��y��7���:��rF�q˫�s�,�8�s��jrV ����ԕD��iqk���/]]���a�<�P�r�t����z��:�<���t��	�^��X�dV��kLcN�FTI�`��}��%@�J�%EN;��89�<���t�i�K��|)M7%����`>vE�s� lr�Q:��Uz�*N�	H��CU��y��9������`s�+j C�NINA%"V2�X���57+ |�%�t���b�rm�Zsp�A�>�F$Nw88ġ�"�X����i0�7\���M�N�� :9x��`�İt��$wI��~R4�r�,,�v�m��Ic͎�I-���z���m�C��P��7I��I)�I/{}��Ic͎�ϕ�`đ6	J�[�B�� P�l�Hd6J`'	K'!B_X!��0�Hb�	�`HFAa!F$�M��h��4浡l3|WhM\`崬�h�`��H04���`����9�Yj�i�WP�%XT��rB-� &f�@�5�).d�,!�0�6!i�yf� ,��6B�ܭ,������jb%MB��c��p�+w��a�P��58�g5��F��3�$��&kLj� @��2�`�"�,U��Kqcf�	B���!B��a����M�( �jcX�{�2ahI���IR�Vp *US�4��U�P�(*� �)G}@D9T��������Iu��-$��Y��:c�7Q����Hǚ���[���I.��e�����9Ē[OMi�iҨ��ZUj�$�m��I.�1�Kd��$c�R�I--$N%JtF�<���박۶N����M�T�+ځ�N�g\�K�V
�J��u$�\�bI-�hn���5OW�m$�wӜI,mk�E&J*/��+�bI-�hn����x�I6��K�6�i$�ݺڈ�8��D&�7RHMʼI$�r�RK��F$��7��$�-4wM��!�����I�/u$�\�bI-�hn�����������k(ԄVCb�'乗�ZI.n�#��R�hQ��9Ē�s�$��}��BnU�I%��1$�7~+�����P���ݝvh��8��4=��v�;��֤��'f�(.�ţ��UݣIksCu$�ܫĒI�/����}�z�Y�]����žu)����	�a��BnU�I$ۗ��]&`bI-�x�I-����4�T`�A8夒M�{�%�f$��&��I	�W�$�t�i�K��T(�rs�%�۰��\�47RHMʼI$�r�RK���x�W��p-$�7w��$���ﾥ�}u�m����m�ﷹ7m���	B�` ��J� Ba d�n���{�W����k+��.tY���vҔ��U�
�cmm�ll��l�����=v��t���|�wϟ0�v�398x��n�r1=��>�X��pk�y�^�x{l�mA�E�����݀����=ӏ+�ONx�sL�5k;�΅k8,�t���vre��;QTv1X�^�vm�ڲ�t�i�q�E��-��)dx��;��[S��s?�{������??�~scnz���t���W^
{n_��������R��t%���rPN��6���Ҵ*��O��$�m��I.�,-$�7w��$�-4v�%)E����^$�M�{�%�f$��&��I3\��]��GA)H�I�I$�K��I%�MԒ8�I&ܽԒX��I
H*R�) ZI.n��I!7*�$�m��I.�01$�v��_<�鰍���?�߭� �w��~����I����Kd��$�:�zW��cJ���b�,*gZ�S!=��K�Oa�q�0�<ms�����x��:�7�I&ܽԒ�/<bI-�hn���ʼI$���MІ5*�)���K��辈���,H��ڔ*F	%(R�FRH�b%H�!aJBKhƺM�ۮ��I�[l��K36s��������⚧R��%J��K����I��ZI%��9Ē�l�-$�;�[Q'QE"�17u$��U�I$ۗ��\��I%�Mq$�i��1)J%J7$r�I,�/u$����Kd��$.r�I9���zb�As2/L'5[��:��bӣ{q�V���4�ѕ��^i ����ۉww{�%�^xĒ[$��I!s�x�Iff�q$��l5R��b�(��Qi$�I����}�z����W�$���9wE��܋5ԧLnF�8&�q$��~�n�m��~�9vǡT�SH�䷽�E�����s�$����ӥQ�ʃq�I{����n�s�%��tZI.f��Iz��i���I$�Ǐ1ЙMJ�_����RK���$�ɡ��B�*�$��f�q$�k]4o���"I�����6,�ۍ�t�;tq����ƫ�9	ݷ]A��&(c�EDDJ��K����H]ͫĒK����\��I%���ּ
�h��W`��7RH\�^$�\ܽԒ�%�i$���q$�i��1)J$���ڼI$��{�%�f$��&��Iy�ZI.�urF�%4�rI9Ē�3Ik�Cu$�ܫĔ�{�z�ɳ�I%�[5*))B�AI�Is7t7RHMʼI$��{�%�f$��{}��~�c�DJdn׵�miΓ�*)�k ��Qu�O/I���4���8h:a���I!7*�$���I��Inn�/�$��Z�IӨ�A8夒\ܽԒ�3Ik�Cu$�ܫ�����6�Y�ǘ�L��Q�rs�%���ZI.f��^���m�w�ZI%����Iu��Jj�J*"(�))�I.f��I!fk��Iw3g8���}�<~�)�I.�߂/��!�����$��5�I$��{�%�L�bI-rhn����{��#���|Yk�ɘv�
|��l[�WRJR��Oh��tmY�ޝm�R�p�ɪ�t�Ph7=,ۢN�.q>��[GRݵ���TP!c�3؅�Ch[�;B��i��]Z�)�z���Iv��ː݃s��;&����e����']%^ݭ��׷Y�#��Ϣh�m����k
��f�.�)��aK�k��a53RYL.kY���蛸n̺n�b��v�x#�;\���7���:69��#Wt�G̚��kq+M�.��)3Չ$�ɡ��BnU�I.�i���H�I�9$�K�v��I-rhn����x�I6����U%߯�TRR4�(���i$��{��$��5KK��W�~�"���s�%���i$�&�N�6R�
����I{睊���-$���Nq$��n����}M���C�I%�伛��t�:)�'��K36s�%��ܧĒ]����Hǚ���ܘ:lߜ��+�ع�Lu�spPH�t
�֩�B�����%�9�NK�NE������z�$��47RHt�I$�r�RK��=)�u(���BRS���ݰ�U_~ � ���04� 6��(@�1`5����I%�	oy`�y`vs_�L��OT$�29���`���8�Y�K��ߦ��߬,�2����I���rK}�˯w����9���͖w4���H�$�I��:q`���n^��X����N8��%H^F{L��5J\��yͱ�B�V� S�4��ۚ��k65���ܼSr�t���QUJl�$)� ����U�GV�=�9��5�F�I���tS$�s�g1Ձ�X��B�B��; ��� �k$�5*��i�`s^E�ks 5�x��`):��z�QQD�8�fm��ꯩf� ���9�uX�
ʚ5�) ��P�pn�n�;!]�n���^cy�J���%&7e� �u ܊0M���l�8�5�Ǻ�fm���<�i*��S����57+ �R,[� ۗ�t�.F�%)��i9��{���f�Xs6XY��������Ҍ,J�`���n^��X�a�{Հ���HX!�Vk�y��r��R�)IJA��;�����+ �R,[�����bT�V����[u���m2r�{��Ftp6�F�æ�=����#t���JQ'%�ř���R,[� ۗ�J+�R�W�+�Ԫ� �R,[� ۗ�j��`sǣ	E5�`s3l0���jnV��X��IUH7"��7�;������`s�9����{M��R�9N6�g1Ձ�����7����B�k�J;��8�#�NKH�	 4��e��@�uɁ�!8kZ4���1w���,l�y6I��I� D�����5(L��f��i���7�(�o��LB.�1$u��_4isY���GBF5��`��ZѶo	L�ڙp��Vqf4(�4˚2�G=��� �*!39�/���m< \]�7�7�bF��
e�i)�,g��#�="������V�%0���|�)����׌��YJ`G	L�x5�5�=`�$��)��p��d6	C��&<J[p��5E$FX0(@��Ѷ%�� E�]�����=vD3D��;�ww:���p 9�[@	 mm�	   m� -Zȳ�w
�U���U�QV�� �u��	Md��,��A�Y�n��v�� R��Hۗ���sB��Ƥ)	�L����t�ҬQU@P�(UFδ8-�    � �  $	�8�   �[p�l     6�-�m�j����v�'K`{�
��k����q��.����ŵ����׫��͸��E�WM�N�gD>���s��N
8:��1��]7(lq�x��g|5��:��v�[yRō��s��Ap�5�K���<��66(�kTax��m�\[�mem�ܻ
���l�^(V=)��9�����te.У��l�--���Ɠ��kn��sD���݂�E�ۓDen�L����|��W�)�n�dp�*�x�·;/m�JiYZˀh��%켘x�a���^Nkh�z����@]�iͼ� ;��]���N�jPm۵�<��i�عݦ/G"m$�n8��r�q�:̉�kv��S�v(N�;=�'��i��+j��i:2α��>��s/[[A�'.�I�m�]���|7-��!\��^����i�%��Ny}W&��S�������d.z��l�ч��ĳ���s��{[,R���:�8�b6j�(i66�nx5m�k�-�8w4�<]�H筺-�,�A�%u�3�6��lV٢v�9�،vu���rӍ��t�ã�����Î �*���� �̯��5���=�̞���EjW{�P��d2����7��q*���H�8#����{b8�Rls�0'h�n��i��n7Z�s�m/DԬ�����BMX��R��ѭ2c'����������S��U���v֙�>۸�k��c�]z��b�;Z����nZ��`՞>K���d�㍦�r�S<c�U8�!.���s�綠L�OC��Ͷq�����q=��4���6�6{t���������� t�� ۈ�lQ8�s�*�E{�K}ހT��Uu��6ڟ�.�|��l祺�<Y�rR�����U���������lC�w����Y��n혚ǭ6�sЮ��8ڸQ�E��q���7�җ�r��7J�n��i�]��b��1OϞur� �d��t�71�� p2c����lz�]����)q��\��xw]��X0vM&h�{v�l�nv�Q�]u֋5�c�[0�*��.�M�Eٻ;`�����^�뵲�[\�[m`2uA�z�m�۴%�3[.�{k���4�6?~��`���n^��Xa�pT%���A)���a`�����`s^�;��R�)IJA� r��"�6T� m��D�n�IC*$�9�4�9�uX����,�i���t9T�*+� �R,�d��4I���"�7�����5On��/kl<��.9��7���x�v56�p����I~�D�����@UZ�$��0�/ �R,eH�͚N�iț�#�[���6�8�Q�6�$�
�	RE�WK"n%��u�ݧ"X�%�����iȖ%�b}���ND������{�������(qvndj�r%�bX�����iȖ%�by�w�iȖbX�}�y&ӑ,KĿ}�u��Kı=�ݜֳ	4]Xj氲�ӑ,K�<�۴�Kı>���M�"X�%�~���iȖ%�'��{v��bX�'�I��v�]j��&����r%�bX�}�y&ӑ,KĿ}�u��Kı<�۴�Kı<�۴�Kı=>��u����Y���%�n�\k��z�x������I����;CfȦ��UUܷiԦ�RAR�m����ԢX�%�ﻭ�"X�%��u�ݧ"X�%��u�݇�Q�"X�'{�ܓiȖ%�b}�k�Y�0�3&�2j�ֶ��bX�'��{v���bX�w]��r%�bX����ͧ"X��$)m�.HRB����M�RH��CZ�]�"X�%��u�ݧ"X�%���,�r%�C�� C� �A�!RQ/���[ND�,K߿o��r%�bX�{��ve�e.�k$�Z�r%�g�2'�~��ND�,K��fӑ,K����iȖ%���'�}�&�{�������ZW����ݷ�����P�(K�|e�����$/7���Kı=���ND�,K������mrӛ��+&���Hb]&K��y�V������Ypu�ٝY�j�9ı,O=��6��bX�'�}�m9ı,O}�yf�yı,W����
HRB�oN�H8��#��Y����Kı<���iȃbX�'����iȖ%�by����r%�bX�{��m9lK������,�ե�&�ֵ��Kı=���ND�,Kϵ�nӑ, 	��=�_�]�"X�%��{��ND�,K�����Fd.��K�f]jݧ"X�~E�￮ӑ,K���~�v��bX�'�}�m9İ1!< Ў�lOu��ݧ"X�%��f��w0�3&�2[���r%�bX�{��m9ı,@<�_v�9ı,O}��nӑ,K���}۴�Kı/������0�ö��Eن�7+I��:�,���g�.�� e�o:h�q�=��ٻ�Ʈ�6��bX�'�k�ݧ"X�%���m�r%�bX�}��v"r%�bX�{���9ı,O}��vfa3R�S5�L�]�"X�%���m�r �%�by����r%�bX�{��m9ı,O>�ݻNEFı,N���Ie�j�f��\�ջND�,Kϵ�nӑ,K���w�iȖ%�by����r%�bX����ݧ"X�%����ܖ�3D3Y5�ֵv��bY�"�߷���r%�bX��]�v��bX�'��}�iȖ%�%�����iȖ%�b}�ݜֳ	4]XMf�nkY��Kı<�_v�9ı,>���ND�,Kϵ�nӑ,K��;��ӑ,C{��>��?_��+�m�ָI�QɵƸw�.�wX�u<9�T�v�F��yE�8z쎔w'+⸌:�M��'Q�2�`�[�~.�|��&���ɷjưx6��Kkf��mn̔�����ʶ���fi�clC˽��������Xvi�*����lv�c�C����y��k�c2�`�c�ѶƝ�Q�rq�r��q�Q8�[�K����/g�-�ҽ��҉̡{M]z�ؓ7u�n�p]��v�<�wZ�;�n�P]���b�����w�x�,K�����9ı,O>�ݻND�,K��{����L�bX��]�v��bX�'k�~�h̖kZ���˭[��Kı<�_v�9,K��;��ӑ,K���}۴�Kı>���ND�,K��w,�as.\5�d�Y���Kı<�����Kı<�_v�9�� ș�����9ı,O{���ND�,K����2�2�.�sY��K�lO>�ݻND�,K﻾۴�Kı<�_v�9ı��{�ND�,K�u;���pt�������#�Gԏ�w��9ı,O>�ݻND�,K��{�ND�,Kϵ�nӑ,K�����߼��ق䗧c��ׂ�O���y7���m�^�x=��~{����������+<��n�Ȗ%�b{�w��r%�bX�g{��r%�bX�}��v�Ȗ%�b}�w�v��bX�'{4t���h��f��Y���Kı<�����=P
	��c"X�'�k}�ND�,K��Y��Kı<�_v�9�H�DMD�K���Ӛ�a&��	��-�k6��bX�'ߵ���9ı,O��yfӑ,�P��5Q>����iȖ%�b}���ٴ�Kı;�5;I�e��)p�[�]�"X�%����,�r%�bX�}��v��bX�'���6��bX?���￮ӑ,K���~��e�֥.k2��r%�bX�}��v��bX�"���siȖ%�by����r%�bX�}��ͧ"X�%���=����lbiP��5�<q2���:k��뗵��v��Ӹ�k��G
ixQ�̷Y���Kı<�����Kı<�_v�9ı,O��yf�E"dK������Kı/{?O�L�pˠ��e�fӑ,K���}۴�?�`ED�K����Y��Kı;����ND�,K��{�ND�,���{!���`7�\>�}HK��Y��Kı=���m9�G���,��L��~���r%�bX���߮ӑ,K��~���ɭfd�f\՛ND�,��R*ő@�N����ӑ,K���_��iȖ%�by�۴�K��T�����6��bX�'h�~�\����jɭkWiȖ%�by�w�iȖ%�b��a"EC�}��m<�bX�%�~��r%�bX����v���{��7���_�ߢzb�As���Q��vPӭش����)!]*�*T��}5��ߗ�{�����)}�Ѵ��Q�����{��7������r%�bX��٭�"X�%��o�iȖ%�by�w�iȖ%�b}�jv��˩�S2k%ֳiȖ%�b}�{�6��� �Dș������r%�bX���߳iȖ%�by�������q�������G�y
�� ��r%�bX����v��bX�'���6��bX�'��{�ND�,K��Y��Kı=��r���r�!n�6��bX�by�w�iȖ%�by�����Kı>���ND�,W�RbH�R0!�D��&�6�K>�]�"X�%�{��w	�3-��C.k6��bX�'���6��bX�'�w��iȖ%�b}����r%�bX�w]��r%��{����~�~��0Wj�u�ƶ�<ͰtlE��G;M��GW��h��A������ߏ&\2��u3Y&f��O"X�%�����6��bX�'�}�ͧ"X�%��u�݂~��"X�'�����r%�bX��wg��ɭfd�f\՛ND�,K��fӐ�V9"X�����iȖ%�b{��~ͧ"X�%����,�r	�ș�����뫘])��Y5���r%�bX�����iȖ%�by��siȖ%�b}�{�6��bX�'�}���\>�}H���nio�O��)"�$�ӑ,K�PȞ���ٴ�Kı;�߹fӑ,K���ٴ�K��뽻ND�,K�S�N�.��Lɬ�ֳiȖ%�b}�{�6��bX�'�}�ͧ"X�%��u�ݧ"X�%��w�ͧ"X�%��"�*-��$UJ!$�R�R � "�` 	!��
ؖHA���Pb��������4�-U[\�����A�{jMvNh]�[�E��K����me��t���:q�v�B�pz.��6��WU է_Z:��O��͌���F!yy٭^[����V��G+�\=�뎺�S�kp(�T�맢�6��&1��/�'�7hHV��W�Ǫ�`��L��/��Y"[;���q���k��O�{vzL[�pԻۛ0�1 l�D�F�u�m�[d���,Ǝ"eb�9:�������'��Ǯ{%8��7�w��7��b~����ND�,K��{�ND�,K��{�ND�,K��Y��Kı;�_e��32��Z&B�jm9ı,O3��m9���MD�>�����r%�bX��rͧ"X�%���o�i��DȖ%�g��	�2e�k)�5�ND�,K���ٴ�Kı>���ND�,K߾�fӑ,K��;��ӑ,K���N�f\&jau3Y&f��ND�,�B��O߿���iȖ%�bw���M�"X�%��w�ͧ"X��*�_�����fӑ,K��������2kY�f�f\՛ND�,K߾�fӑ,K��;��ӑ,K��>�siȖ%�b}�{�6��bX�'ޓ��.[��Mf����Y��|��r�Qy������Nsd��:u������w�1�l�˩f])�f���jm<�bX�'�����r%�bX�g��m9ı,O��yfӑ,K���ٴ�K=������������5r���~oq�ı<ϻ��r�`���T�pHJap1�D�p�$��h��"�`R�����q��$HW	���X@dA,I�� ���+6�+��?D��K�~��m9ı,N����ND�,K��{�N@�AL��,O߉���?[u5K�.�kZͧ"X�%�����6��bX�'�}�ͧ"X� ��=��߮ӑ,K��;��m9ı,O���pђdֲS0�[��iȖ%��(1�� L��{��iȖ%�b{�_�]�"X�%��}��ӑ,K�@&D�~�ͧ"X�%���]��f�r�%�Z�ND�,K�뽻ND�,K_��� 
E�뿿f�Ȗ%�bw��rͧ"X�%��ޗ�)!I
HX�ʢ�b�L�󋜠��b�uʽ�/Z�E:�΂��=q�0���u��[�;"��tn
~{�7���{��g��m9ı,O���nӑ,K���ٱ� EX!"dK����~�ND�,K�j~��.50����3Zͧ"X�%����m�r+�� B*dL�b}����r%�bX�����iȖ%�by�w���Kı;߶t��2kY�kR��Z�iȖ%�b{����r%�bX�w]��r%��:B$ �H�	Z]�D���0�kf�b�H�<=>E�A=�����aǕ���֙� A�P����� ��9�L��_CI 5$��.��	W��	��
�>4?��C|�e�#~%S8�rI�yiY�l����#@�"�W��y�ɌV汁�O�V��zF")�
��������x�=Oa��F!�$�Zc$.&�����{i"a�xa��4�@�� !�)���0��3A��)��6ī,0�mI2!�G������E�?<v��Cj������P:�@4�	���Z
�(z����GX��n����X�d@�>��~ﹴ�Kı=����r%�bX��GN�K2��L�k&�kSiȖ%��02'�����r%�bX��{�6��bX�'�w}�iȖ%�E\��{��iȖ%�bw�7���35iusZњֵv��bX�'���ͧ"X�%����m�r%�bX�}��6��bX�'��{v��bX�'�v��yf���`�!y�=#�=47Fv�s��邋���ӝ&V>{��o{��ߛ��~h�ٝZͧ�,K��o��ND�,KϾ�fӑ,K���n��@ �D�Cؚ�bX�g��ٴ�Kı?j���Nd5���5��V�9ı,O>�}�ND�,K�뽻ND�,K����ӑ,K�����9Kı;�]�٘\ɗh�,���r%�bX�w]��r%�bX�g�w6��bX�'�w}�iȖ%�by���r%�bX���ܓ.d�h5a.�v��bX�by����r%�bX�}��ݧ"X�%����iȖ%��b�B(*�.H��w�iȖ%�b}�s�.50��k$˚ͧ"X�%����m�r%�bX������r%�bX�w]��r%�bX�g�w6��bX�'�[���\�9PRLj�*l8�����Y����Z�u�˺#Bn+���������y�̺ջO"X�%������Kı<�۴�Kı<�~�m9ı,O���nӑ,K���:N�ٗF�f�Y5sZ�ND�,K�뽻NABı,O3߻�ND�,K﻾۴�Kı<���m9ı,O��o;�h��.�5�k5�fӑ,K��=����Kı>���ND�P�,O=�}�ND�,K��{�ND�,K�&�hIB*Lc�����Gԏ�V��m9ı,O=�}�ND�,K�뽻ND�,U,O3߻�ND�,K����4\�ֵ-�u���r%�bX�{��6��bX�'���6��bX�'���ͧ"X�%����,�r%�bX�G�X �B�=�%�3��:Yk��gb�����f��g����%*�+n� �R�U]#�k5�lp\'[����׭.c3�Im����;�T&ݷ��h^F͞��	p�㞍lp㶸��a�7$�r���g���Ѿ|���ʢ!����孬���i찷�8�8!�#p�Lzx{9�c]��"��"Og�'�[�ƻ����L<�;�	�c��=�������WO/'��'-�sy��d*�%ڸ4�q�r��+s���r�8��sп}�����?:���^#��Yu���%�bX����iȖ%�by����r%�bX�}��ͧ"X�%��o�iȖ%�b_��gre�d�N����m9ı,O3߻�NE@�,K��Y��Kı<���m9ı,O3��m9�B(+Q5���O����&jaML�I35v��bX�'���ܳiȖ%�by����r%�bX�g{��r%�bX�{��v��bX�%�~ΐ��Y�34S2��r%�`��*H2 �D�����r%�bX���߳iȖ%�by���r%�bX�}��ͧ"X�%��tt�ճ.��kYusZ�ND�,K��{�ND�,K�$W߷��i�Kı;�߹fӑ,K��߷ٴ�Kı;�ҝ/
f��Me�[�.�z\v��l򽄹���k`�*sneln�-����U�8��������{��7�����ݧ"X�%����,�r%�bX�{��6(�����$T ���L�bX���߳iȖ%�b~������T�8�p���ԏ�R>����m9
!�X�AKH�P�"X�'�w�ӑ,K��=��6��bX�'���ND��O� �	  0 @P��" �&�X���f��MkRٗS.Mm9ı,O���iȖ%�by��۴�K�!�2'�w��"X�%��~��r%�bX��]�٘\ɭf�є��SiȖ%��P�(�$H�@�!��~���n	 �w��͉ �'����n	"D�߷ٴ�Kı/~��ɖ�&N�R\��r%�bX�{�xm9ı,?�"��A��T��@������ؖ%�b}����ND�,Kϵ�ݧ"X�%�}������qӶ��8:�)P�%0��g�*wv	��)2���`�9zSf�fv�Z8�D�,K���9��Kı<���m9ı,O>�{v+�! �AdBAșı=���m9ı,K��s�	L5��3E.\��r%�bX�{��6��bX�'�k��ND�,K�~��"X�%�����Ӑ@��E �G"dK��~'�[2��rf����jm9ı,O{�߮ӑ,K��߻�iȖ:Z�D
dL����,�r%�bX����7����{��7����|j�SP�m9ĳ�@V, �F!�EȞ���ND�,K����6��bX�'���ͧ"X�%����nӑ,iR>��C�$�7C��*��Rı=���ND�,K� ,�Y$�����yı,O{�߮ӑ,K���}۴�Kı>=���!�b�⼴��q�|=\�$n����=�a��8��TV���x�`��Y��Kı<���m9ı,O>�{v��bX�'���͂?���"1$��>DȖ%��~�ND�,K�f�K�ff�4f���Z�ND�,Kϵ�ݧ"X�%����iȖ%�b{�{�6��bX�'���ͧ ���#)�dL�b_ݟ��nRa4jIsWiȖ%�b{�w�m9ı,O~�yfӑ,K��߷ٴ�Kı<�]��r%�bX�{��;�d֌�jf�IsSiȖ%���"�`! dO����m9ı,O~��M�"X�%����nӑ,KX�a�$� 0Ả���iȖ%�b^����jf�f�\��6��bX�'���ͧ"X�%��Y('����i�Kı=�_�]�"X�%����,�r%�b����8�mr�7�b�v��c�靏�SYlB�vgI[�p�n���A�u�eֵ�\֦ӑ,K���w�iȖ%�by�۴�Kı=��� �	șı>���6��bX�'�������3H�|�~oq���Ǚ�{�ND�,K߻�Y��Kı=���m9ı,O>�{v��� EC��0R
�j%���MO�$���Ꙅ�d��m9ı,N����ND�,K�~�fӑ,K���w�iȖ%�by�}۴�Kı>���Fd����e�[��iȖ%���B`��;�y�m9ı,O{�߮ӑ,K����iȖ%�b{�{�6��bX�'{5����k,�ѪYu���Kı<�]��r%�bX�+ ��H���]��,K����rͧ"X�%���o�iȖ%�bqA����������2]��E�z��[/����1-++Uoa!�U���Y��scp�e���gj�"|�ce��ش��r�v"@C��{m���� �:��\JiKq7F����m3nt�(܅e���2j:E�&���9�-6,µs�����{N�K��;�%�������*�ql.�3��u�
Os��=������X�Y7���NON-��Y���B�l \��q:�gU�l�q����.�� �ޛj���t������1��w���{��~�]�"X�%����,�r%�bX����6��b�|��,K�����Kı;���?fY5�,�����j�9ı,O~�yfӑ,K���ٴ�Kı<�]��r%�bX�}��v��/�A�L�b_߻��Ja����)r��r%�bX����6��bX�'�k��ND�,Kϵ�nӑ,K�����m9ı,O{���&hѬ˭kZ��M�"X���(1 �'߹��v��bX�'ߵ���9ı,O~�yfӑ,K�FdO{�~�ND�,K�ݛ��֋.j��Z˚֮ӑ,K���}۴�Kı�"��s��O"X�%��{��iȖ%�by��۴�Kı:}��I/Ne4�G^�6;T��v�����&��ֹ޹��|���X�dݭ/O.�E=ߛŉbX����ݧ"X�%���o�iȖ%�by��۴S�D �&D�,O{�߮ӑ,K���^��Fd��j�2�-֭�r%�bX����6��:�u"��"
�$A4���";r&D�>�۴�Kı=�]��r%�bX����ݧ"X�%���}/fa�V�h�,���r%�bX�}���9ı,O>�{v��c�� ��j'o�ݧ"X�%��߷�6��bX�%�ӳ�2\��kQ�K��ND�,Kϵ�ݧ"X�%����m�r%�bX����6��bX�~��D�����9ı,N����0�іj����v��bX�'�w}�iȖ%�b{����r%�bX�}���9ı,O>�{v��bX�'���azf��u���rK���5[p%�<&���d� ��۴k�{��[R�h��{͐��S5s4R�֭�r%�bX����6��bX�'�k��ND�,Kϵ�ݧ"X�%����m�r<oq���?n���f롙������ı,O3��6���bX�'�k��ND�,K߻�۴�Kı=���|�~oq��������?�x8f���r%�bX�}���9ı,O}���iȖ:@�6RB�ԫU(Q�BRRUe�H���	D�H�0$*P��(4F �h��m�9��M�"X�%��}�siȖ%�bw�����a�3$�]\��r%�bX���y&ӑ,K���ٴ�Kı<�{��r%�bX�}���9ı���O�s�T'$�m������ŉ��o�iȖ%�b��"���6�D�,K�����Kı=���M�"X�%������]jYum�Y�n��5��^��5:c�\���̓n�$l�zyR���a5��3SiȖ%�by�����Kı<�]��r%�bX���y&���&D�,O����ND�,K��?O�2\�Y5�d����r%�bX�}���9ı,O}���iȖ%�b{����r%�bX�g�w6��)�X��L�bw�O�~Ʉ֌�T�d�5���Kı=����iȖ%�b{����r%�bX�g�w6��bX�'�k��ND�,K��ΐ��S&�4R���r%�g��1A�
1H�j'~��m9ı,O�����r%�bX�}���9İ1C��1Qt�jD�]�,�r%�bX�wGN�*�Q8ԍ���}H���#�����Kİ�
��Q �����ObX�%�����Y��Kı=���m9ı,O�5ۇn[��LS�.M�櫛T��r�wN�;[��U�:\j���ӣ���F�Jg��{��"X�}���9ı,O>�yfӑ,K���ٴ�Kı<Ͼ�m9�Gԏ�|�(��鸔$q_���Gŉby�{�6���T�Q���2%��{��iȖ%�b{����r%�bX�}���9ı,O���٣2�j��2�-�Y��Kı=���m9ı,O3ﻛND�Q��	��=�~�ND�,K����6��bX�'N���f����Mj����r%�g�$���ٴ�Kı=�~�ND�,Kϻ�Y��K�T�=���m9ı,Kߧgs)rSZ�JK�fӑ,K���w�iȖ%�a�c�~�ͧ�,K������Kı<Ͼ�m9ı,O���S�K�J'��
#�`HF&�J��ń)��2�0	"2h�
.)6t���e���2"H�!&�@tDa0є�'��f��0	68`!L\�[�<�A���5KRֱ�$ Q�������;�ϵS�����m $ u�6�m  �� qv4���o=��eU\ȫs۠�u 3D�=v��#�e��@n�)�ջ[�e^��9����'�a�˯BL�j�gm�vm�8 li6U����     � �� #i6�c��  ��i�     �`�m�O�{IGaYG�'�"n2i�a8�uƐݚ�:�&���!���BPnˁ���gbMٔ�����q��<�+�͵��	N,��>n���q����)ٶ��fn�>��:�+I��US���,�˂�x���`�,��p$�u���:1u5.[ni�j` ��՜�ĸ�L�i"9�wFwFy��gv���5�����v�u�^.cld��qy�ŵ���On�u��ϻq�w.U����wn5p�kl��Z#��C�lUR����y}kM�g`�x.NmT�PSm�� Ec5��ɜde��;
��N�ssA���f��nt�7�Stm[#V�/{n����e�z�0Yx68�b��,�5c��n�����o�3͝�c\֋�:�B	m�΍���u�k�ힵ��=O$���Rg�Q:l�Q��ՙ��쳗'p��ˌ�l��:�e��V�[ڣN�:�qL���I��';��l�;Z���jR�A�'�Y+zZ�'D�Ĩ�ke�-�h�;�vhڳm<��|s�M�k��� u�c�� 1u��mu�Ȫ ����dZ�� 5I����;[pثs�!�Y��9{u��4i��)��Vw6x��j�c�VA��ȵ4ں�I�Ι�t�����Bc:J�6�m��Ӝ�\�J��^,�= F6��P�Y���s����d���)�F��e��iy�.ΤOmbK5��Ɏp.���QA�֌)�k��Q`��C��N.k�#A���V��#<sp"c�9��n�9�z��(e�0\��N�i	���周�M�qt=�� z��/�v�C�b �E���[ff��tkx�F��/Dm'Y6��v�N�d1����V��W"Ӆ�y4^���	b2�.7n�=������N2O��[n9���<�bl���X�nm���1�.v��r��-��f���{�2��l��KΎ��9	豕�'8ɹ����&a�^8sm��s��%���%F�ˢ�u���9]g�g�y�։��7�[<��`خ�����Ӓ^S$ܚ�Rt�餪����ێs�d��X����3�S5�\֯SȖ%�b{���ND�,Kߵ�nӑ,K��>���G�,K���w�iȖ%�b^����f���)r��r%�bX����v��bX�'���ͧ"X�%����fӑ,K�����m9���w���߿���=���J&�����,K��fӑ,K��o�iȖ%�by�{�6��bX�'���ͧ#���ow�߽����F�fk��x�,�#������r%�bX����Y��Kı>�~�m9ı,K��w[ND�,KޓS���S3V�j�SiȖ%�by�{�6��bX�'���ͧ"X�%�|���iȖ%�by߷ٴ�Kı<��ߦv��[d�%*�n�X7n�6��\dutx������Ӳ������O���qT/$���{��,O��ݻND�,K����ӑ,K����iȖ%�by�{�6��bX�'N���eԹ4j�j��ӑ,Kľ}�u��: V�3�B�H*`,X( )Ij�!�1Hi*&�#�,!	�
�|U2&D�>�^��9ı,O>���iȖ%�b}����
HRB��4�(�Hs��Iu�m9ı,O;��v��bX�'�w��iȖ"�%�����iȖ%�b_>���r%�bX��O��n�e��k$��]�"X�%����,�r%�bX�{��v��bX�%�ﻭ�"X�%��u�nӑ,KĽ�s�%0֮���K�5fӑ,K���}۴�Kİ�}�u��Kı<���r%�bX�}��ͧ"X�%���oN\�V�)Ay|�عv�.���v��g:s�V��jhQ���CΠ��t2PT|�~d�,K����ӑ,K��o�i�
HRB���d�	.�<��`n3����)JG#�9,nM,f��ν�`��`shf��u7�R�����Ssg,K�JȄ���@,b�`f:�,$bh"X�G�(Q��b"#$��`no4�1Ҝu�LNHۦ�I�X~������w}�`v^:��!$��d�5m:�iT�8����r^�9X91�|�>�n\�|�6+�������!�V=��y��InL0Sll�2$necZ�4�t���pRHMs������`g��؄����K�k]y))�*q�r;���`g����|�=/_��(P�߼�QBa"�7&�E���+ �%����s��>��*#�_�֜jD����U}_R]�zX��vsv�i(JTD$�s�l�9O��y����]]�����s��>� kݖﾪ����z�ʂ��Q��n�O�pqQ�\��wb{z�fF֛s5�8�t�����ҋ-]�鸔q���֋:�U�s7e�չ���t�\��䉺o�3\���SsD}	%	Uo�r�s��Vsv�`mkǣcPL�)H�)�k��Q��9Ɉ�T� #!*d��Ѩ[e�krtQ����ߪ�{��%�����;���s�)9���������J�ν�`��[�y~��ܓK�}I"$�$�F0�(�j�"$l�{����^���άh��EH��j�+J��<-�[@:�t�RY-sjd����cJu�g��t�$�A�n����v�za�+��c�� &�*%��d����]\��#��l)��۶6(:۱عN���Y�4ڕZ�m9�;jݙ�c;��]�s=�9�ͭ�u�d�6$튣�1�3�r������gsvN�պ��2̦j[d˖�u��~�AP�AP �(UD`�b �X*�P��{��mߝ��d������^8���m1m�h=�T�u�YknN�;���p݉�v^�I7	�����`��`unk�UUW�qo���;�^�C�*'�(��|��!$��%�	U~ߪ�{��%��{�����)
DRq��K�r�rb0|�)�o9x�Bz[s.[�.]I�?����6ξ�l���ġNV��6���(�sZ��35��ܓ�3�䟁���� ���������T�iKB9RN[���s���WVzx{1���]'%�� /WE�,��H�J865�QH�)�s����V�&# }N, ����G�x�R�5��䜿{�o�T�"�UC�(Q�
����%�����,=�u���QS������μٳTB��=�y`zu�X�M�r�UUׅuV��8�y��5G+ ���,��c�P�J�ƤJH����aDB�k���ے��V9�1�S�x���m�xf�M"�n/ep�Y{v���5�����4lL[Lg���Q�f�Ww�j�V�&# }N/�ڀ�?^�����ԛq�v;�h�}�RP���/�s��_~M�?�?9`v^:�1�,��rD�7N"�μ�`��r��'���E��"���"�IOvo�U���K�YL�*x&H�M8�?�W�}Iw}�`u{|��w%�J^q���M���T�����k��;/XB_��	"~��xk��`��`�-I�HM�r�(�uuإq��]�nݝ�����إ�C��j�rSu�pEN0nG�3}�E��y��9������`���I�E�tO*�%���s�J(���Q��������;���;���9R�pr5$� �7���՛	BS8�nK�=�s*=�R��#�G$������ܓ�3߮���*� !��[͝�{C��ۍJ�
8��w%��B��g�{��;/X��{�#t�Q�yh.�=�<=\�&��ch��fγ8{!ɶ�R���<3<���ԕZ0���r^�9_��}���h�=^z�65�8��s7e�P�}�*�'�����=X��$!(�Q���$*��5G+ �s�μ�`��5v�֡��U8«��Q��=]V�{6�7��s]�n���E�t�J�3��$�С*����?o�`{�ի��M���S3]Vm̀��la�y����blk%*�+oa!��Z�I�+�e@1�e��f�k�vm)�;F��n ��]�<a��q��B� �n5̼m���l��&8���[=��`7R��q��]��ʜn�J��[Z��� ����Ǉ��r��V���<�(����y�W;d�Mv��^�6:G�=ff�o��1�=���ӎ9��m�ZsqZ���{q:��N4M�����li\9'8m� Nn��s�u�٤���ߟϲ�Q��;��{ }N,G�wh��H��%�Ź��UW�_������~�����X;�,�[L6�nE*+������q`���j�V�N�k�	ƔT�i2U�����nMٰ=�X���ce��YL�*`�!�4�f�8�5�����μ�`�?�-�l &�s[l-S�����cm�9�l�g��j�L�ں��w��c(a>�HNN���;��Ձ�y��9������Z�'TT�
�r�ce��
B��P�(@g��w6X[���U_$�� 7D��j�º���GS��r^�9X9�;���9R�u�I�������Uf��,���=����c��T{$E(JD�I�X[����u`g^j�f�;ZeJ��	!Q�s��N�=���u�CۭǩN�<�]���G���z��)L.�nE*((����u`gS� 5�x��`W��t�E�WTU���`�ŀ�Tr�rb/�_RG��_�Ơ�!�4��{��9~����|M�BZv��M�FV���\ �d�#��M�P�E��T�6$�����0�b+I"�"�G\��5��c��k �<P�%�g9���I��]���.C32r�ZaD�f8&�7���>�
ZJJJ²���g��VA<"���b��R^_1fb�DӰ|�I�s������t`C���䲲��.g��
��Iww�!���\V0�
JB� �� �c����A�)EւH��"G4`�ȸ�(`3Tf٭���B��5 �d� �"�
��0H �! $_�G�q@=�EN!��@��A���pQ
Y�b0�`d%*<P_�hBrX[�����μ�a睊.�,,�u�SN	20NG`w7m�q`�/ ��d�^�W��X#u�F�\����mV�T��o�G|���t�ݦ���!R8 �H�یN#�n=��q�X���P�d1�ܖ�⢵ �Ji�rE$V�ݗ��#���`f�֋:�U����J�"�G'9`v^:�=�ܖ|�S/)����,�[L6�nE*((�;���<�~��N{��܂"`
�9~���������mD�N"�μ�`yDO��:�^Ձ�n�2Hr��<�H�l����n���S�.�<닂x^�۲��v��e�[.K�r1�m�?�^�9X91�q`d%&P�}@�����}I�����{�`��`j�c�B�T�8��`{�,:�6}	)��w��ݛ �Ǡ	���j0Q8�}_}�~������l7�`g���=�ܖ�⢚���M:�H���9�����V���{�{�7$����"��RV�RE۽��ۻݹ��v>�pMuM��Ѕ>�t�{9"��[E\9�T�v�F��yL;�5�SJrr;�d�1���r��,q�qe��*�q���^�}E�k�_g�'7`۷l�Ün��q/ny- ;Wig��qm�k�E�s�]�'v�(l��X�+��sN��r��slf�pZyûm�:�V���6�s�Zw9wAӥc�7<��sp�q���9Kt*�{���w�]~~C�LR.N��5�,�9�._,N�{j��Wg!z��1��w��|��Q�BR$RH䓠{�|������`��`whb�a��r)QF����7rXu�l��,�77�%2=��z6�J2&8�qys7e��{���n�,�z�lI��UMrl��,�76����RJsx�X���12����3�uX��`)ŀ��B�TO�ČWj�:�����m�������Y�ny«���O7= t�-c���i���~��%���s`����B^���~� ��?�$:�TMD
*r���W�W��JD"�P�T��X�{V���XݔǨ�(N��)"���;/Y�P�q��V�{6�.S�8�P���9$�8�5���E��y��9�����Ŵ�Cm�q���K��%����o�r��oͷ���������Ԓ�V��v�d��u�!�{[����>�Gun��5�R����35�,�c� �7�����	DG�A��Z,W���A2B7
i�`��D)�ӯj�ǻrX��6 ��X���TrXY�����(��sՎl�,>YI�(�p��8������q��+ �n��w]�n��I'R(&���3+�q�X��X��K�	$�[~���sm1[a�;
�sN㋗R��C��ڗ�����w��������H����X[�����μ�`neG�JIE))$rI`qnk�=�ܖz�̀w��Dɚ�'U%SrFEvo�]Xך���,-�vk��ci26���&J��_T(�/8�l�w�e�D4��E@0���K�*8�&6��[�A2c E� ���
"�(��N�W�֕EO	��9U�T�&�;����%�׵�1�c>m���.O�l�@��u��^����:|�-�6�s�{2��eӜ;�k��	�r��u`{-X��?B�� w}�`yek�	P�"n�`܎��n��艑�=� ����x��2�E$4�L��:�g^j�f8~�ꤸ�5��z�`gvS�b�(R��)$�|�L������ڰ=����c�s*6����NH�����`w7KVz�̀w�q�
$D��=��~�2�-Uu�2�v˕)�����U�TYZ�8[M��;m%�WV��']+��n^��7k��q��6���L[6�r�-I�3���5`��5v-����=b{���H����ݠ��A��v��qx-�vڵǏ�L��Û]���5өT3�Yx�
r���ackm3�Ton�^sRA:��f:��s�(ջ��nv�����Tǎ��X-��T��3Ξ��⵺\s!�z6�s�6Jx�j<�������E�閛l�2((��3���S� 5�x��`W�R�i�EI8�:�U�s7e�Ź���n�,�x�lj	��SN+ �7���՟D$��O~��`k��lp�X�j�*�(�NK�UU.�o���t�`g��q�X|��&Q\DM����������V��. w}�`qnk�;��4jS���T�خg��c�ո���]Rc�iF��N2��<;��i�H��A8DF�Vu� �n��s]���.���c�LR�
TRE&�䓞���UO�� pt@�=\�;��Vu�s*6���D��$�X[����u`g^j�f�7�~z6�$dPQ�a���:�� k��Q��w�J_����Օi*/��q`�/ ����]XKk��� ��2ph�WVI�Żp'9��n��eb:���r�:S�2B7
i�`��`qnk�;������<��`�6�&�R9q���9X9� ��X���"��Z%C�#$���v3t��3�5nw�*C�)@*� �����B�!(*j*)�� A��"P $M4}UU������5g�; �h�#��բ�� ��X���9G+ �4��3��R(1J�)Q9�fl�>�>߫�f��j��Ss`}��[��n��Wvn�y6���ܢs$�m��;
2uh�f��;R�9��sr�]�~�� �!��T� 5�x�I����m�8&�9�����H�~���X[���F�Қ^���vU���`��� 5�x(�`�.�mlZ*��L�Q�X36X����e�D-C�ǹk4��M��I,��v3t��3�uX36X3ʖ�7EHM�o���@������z�շp��u�|Է,�ˮy�帹9u�qrSlnG�;��u`g^�n^�9X�-%j�jʫ-T_��"�n^�9X����u�JT�ʉ�G�s3e�չ���n�Vu�s*6�+X��ݫ���9G+ �!��T� 5�v����]F�6�q������Ss`�|�=/X
đ���[�I	P��J|A�`LS	q"(60%	�6�4Xф!H#	#�ʰ�YM&���f���
����qLᢋ0��Ѕ�AH$�2i�"D�����*bC^ILa�
�,+"¤(B��a
�SJrTF1o��l�hR ī#l�&��0ł@�#.���U$��H��B-1s[�m�!$V,R2D�@�+(ư"���`@H�B6�R0 �\E1���@���a����6�JA׋��s�[���ۀ�[@� -��   �` ;Z�ճVβ��� *��RUX�+[]�u ��(@�.�b�=9U��B�U��
����{5X��kIekڤ�8͓i�]�8 ڶ6Z,-[�:��[@  � � m�  $m&�    �K��m     m	 E�l%�:mZ����,�18��mr)����t��[��ӥ�u����76��R:��le�T����=����F5�Ŷܗ)�����=��Y�5��=b�j��٭�f����C��B�L�:LJ֩@U�5��V�n��[�Ì՝�;L��tP�]@F�̆�P vʻGn�gC�7,�x�ָ���۶r�Êt��Wn�"��������ڌ{Y�\i���Z�UWI�<;AƋz�e�C�6u�0�m�R=����`���7���n|��׍�j�盆Sr%����p'[g]xa��#]/L���gV�Y��dx�p��e��Ԛ,qDV����o9d%���6�M���7�Q��3H�g&��	P����˫��t�Ӷ�I$ҽ����َ'�-y@���-Dnkq�9��۬%�meB�b5����6��P�U�*��M[H����u&TC��0veٕ�7OX��׬��H�կP�%�eL6�ꎙ���vh��-�y6v�;i�'W�.49�̦�x�'Fu�aIQ;X�x��`M�1��+u�u����M6��<.�zy�j��VihBGt�jݼ�5�J�"�6�*P&���n,`�H�"c�H�l#�8��s�[��8�^�E>ΗS]� [V�l�nW��Rځn)ЁB�+�D:��C�e��\�fg�aCW=�g��ݳ�v8s۵M�N�0�S���7�v�/n�8]�5ٸ�=��9�yо'5�;.K�����/���ٹ���혲]z�kNĘ�N��@�2k;Y�d�����Y&�Q��"� ��J(z�_9�%��U��]\s֝v��Ȁݛ/��0���b�U��R\� �^������ܜ ��u�i��mv��g:�'W@(y�9t���	���s��f��ݳʃv�kN�2�Z��;)�XλjE��8G��;�csmkm\m�F;"��f^[==�0a�u�γ��v�v�sc���n%�Zh��x�'����/V�SV��ɩf��mOG7���b7LUW����!��&�i�����l�%g>M�I92%!\��M�]���R, ������k��`=-AT�d�����9������`s5ܖec����CY��J�H�q����߫ �!��� kr�]�u�T8�J��q�����̧��X�%`����E�*��]Q~����X�%`�.�}���
�_��@���R�$q���q:��qy�7i�"H,��l�x.����u��K)J�Q9	"�׾V���]{� �{�`{v�m����F��G.䜿}�nh���!�"ШQb� �I �!D�Ҍ0@

2s߾�7$���V1�q��߇Q�����H�r��q`�ŀj�V �R[)��(��I��ǚ�c�V�U.�r��z/
� � ��%V�t��5I+ �!��� w��N�T��A���$��.zY�g��C��A�X� ��VRj��t�玍�����5I+ �!�����X��:�*(R�q�����n�Xs�`���jlP�Z�Z���$�Q�`fV9�=��,��a
 @��	"��PʥX���;�������F�H�*(�r�&�T$��;�����X�2Ն��f�Xݨ�h��J#RJ�B��V������z�Tu[�)�-q&fܼ��������n=�OX,y�=�Z:9�i��g���ԕ?6ߟ��3�t��;�ŀj�V�_�)~�8EI8�1���W��Gu���������E�ͭ�ER�I�
8R����nl��VlB�8�nK��+ �4��&S�R�S�8�-�w$�߾ݛ�{�{�ܘ�6�
��,�vV:�*H:lNG`uɈ�S� ��Tr���W���m�u�F�\����q� ��p�/;����ݻ�է���q�ju���a���-�K�O� ��Tr�rb0��Q�ҕ*&�rE`qf�8�5��m���y���ʍ�H��H��� �$����q`�J�;�H��t�����I����Ձ��́��ua�Q��ڰ�*��*��Z���UU� �8�]%`���w���7$�1x��BV�����)H@�R�����ЅYd�T!F�!k���~���� f���dR;��JB7V�Jc�i�u����V��CJ��J-t�����S�9��R��ל���l4Z�Sa�e@Q&���NYH'^FWZ�u�����L�9�.�����u�'��vrv��W7����5����U�3p4��9�+/F^i���_��§�lNy6C�1�2V�w�K�A蓹6����XW	�j���CZ�R^,E�Վ��!�Ef�'(�`�;�sEї	x.1vM<-���\�s�^zc\%���Ղ�?�j��`���w9��s� HC[Hj�*���	�`qf�;����U������ꤍYZ����JAz�UWXs�ΜX���NJ�:�Dͥ�(*r$��U����S���00���t+��իU~��X���NJ�;���;j�;��:�ҊPG�(F5R9GY8�����/�
��8f�:�:��Ho�W*�iQ	$NH�,�v{�a`wj�8����3~(�*lq�G`w���7�v	'�	Չ�Q	eLp�>���A��IQmax�B���������Ala��Ɗ���4���If����ݫ��Ձ�8�e�"�5���U����g���y����OV��8�$Dq�H�]%`���w9��s� HCX�j�*���	�`qf�;����U����`w��6�@��$Wq�^{r��BJyf����R��r��5��:�GPJ�AG���v{�a`wj�8���,�vV虴�EQB:��8�]%`���w9��gsn�R��F5 �I"�8���_~�76mD+)@,A�H�+��(+
���h�1b�b��bD�@�P
������ͻz�U���n���Q	$NH�=��K2o������9׺�.��Čߝ
Sc�R+�Ͱ�7�E�j�+ ����2���[;RJ�Y;v����\v�{X��f<���QR�\�l܃���2Y[o�o�����7V�X�RJGd3�Xi���S�2DG�����RGVj�w��:��bņ1��:U)>]`)ŀw9��oT� ީ����2
8�)���sl,u����¡+���%	.�c���MjN��)a��U�ν�`qfk�;��;AYSi�J�fS�X���9���ek�y���2r��z����R��H�9�ν�`qfk�;����U���T�4��뻻X��`�``�ŀoS� �1#7�Ҏ���v{�a`sj�9׺�,�vnJi:�MB6��J�0t��5t��jnV���ͧ�GQ�L���"�8���M��;���5Ӌ oØ$�����.�8�X'm�խ.��mXӒ�����ۂt-�5UJ���v�W���s�t��N��S�s��;dW�ų��;E渳x��.�F�3�9�;wWd�'8.������xN�	σsq��cq�;����X����l��m�����������t�؎�m�of���n�ǝt�%J�x�eٷ5lvN{u����z{�����ݍ�Y���w����T>x� �U��7�r�jN"˞�;���f��w�ƹ�-��t�&�ҩH��}w���sl,c�Vw]�����)S*)�r<���]8�NJ�57+ � �Du�AB9`sj�8�u�Y������ͺ�F)D���ԫ��jrV��X91ǗK����@���JR:�H�,�vsf# �N,z�X��^�,���(T��3�{k�f�u�̇9�m�z�)����w0�����|:Q�T�Q�G`s�����U�μ�`qfk�;�)��](ۚ�%�Y�'=�~��@�z��~��lK{V|������Oj����'	d��6)��{�`qfk�9��E��y��ՋMcM�t�R*}���̕�oI��5Ӌ ާ �yנyQ�R?�cr;�ݴX��7ˀw�XY��mmM��6Sm6nk�&��k�cV��8��3���u�ۆp�":�蠡��1w5���V�{�p�33n�Q�)H�*G���q`���o;� �9Y��|��u)���P��X^�;�ɳsF \�Fa�J���0a
�!��̦ͤq�M,bGP0T�@!��@�1$"���)�� �6A�`@7Y0"HBNR��&e�����@|� "A&a���!���:7w�1��ٱ͎,`A�M��$X@/7�Np��H0���C��`�]��j�AI
.����$ѤH���(��	��@C�?!��� �*>�&���3�<x p �@�Ui*J�{�Ձ�M̀y�2���J�j"H�u�s]�μ�`qnk�;�)��](ۑ�$����:�;��6e���s`j�U�ӏ�ѝIV�w37=>5Z$@מ�o�0N�m/lr�[�l��E��a�i��?�s��`���oS� }N, ��cLc�R�S�V��y��μ�`s�5X�X�B�>�F�6���ާ ��X�8����5F)!B/��:�E`g^j�9ך�k�V������/mX�ۥQ��dd�E`s�uX���d�.����޼�`f�[J�	�I$���ʊK�^s1å�s8�mc%�^:DM&赥ʝ��v�PJQB�`o^j�;ך�]�v:�U�nRKi���J�jF�V�X��"ɹOf��V��Վl��i:Z(ۑ�$�����`s�uXך����OV�� �"#��wX������;�ŀE�V NţcT�l%"�G`o^j�;ך�>�Vg�Հ��
Q�2��S��j���3cY]ڣ8v��J:�p��E��UZ�R�	 d�[3���F[�8-�� /2����>v�u��Qۮ[���4n��kk���\��l\��+Eӳq�x�:�ӹr��ay�(_=�'���v^��ؐ�ղ��r�*�S��*ծ���R��wX�m���n6���ms�8m�㍢�ۚ=>m��q��0���r�S5�@��5��Na�\&��B�/+��㮙�\p�������<|�nf�#g$�ḹ9zۇz)s�h�m��V9X���	���9F��IR�/�X��v����5t��N�޼�`nf�(�JFFH�R;��+ �N,��X\�`�XQ�<�P�8���Vz�U���������Io�E)6����޷9X���	���x��e+ct�Q���;su�`;�=
���û<A���br`�:	ɑ(y��2���>m�ϱՁ��u`?V9�(P�!�Of�����d$Dq��vw]Ͼ����b��W�ܛ�=��Iϳ��j�k��-i1��T�H��8��qa��~N~���� ��":eE"tƛ�X{���ܛ�`yf�����'S� ��!%J���b����"�+ ��V:�X�8��t}5l�&l]S�n.m�"�9�9�X��	�g�ujx���j@�\ҍH�.�z�U�μ�靖<�|�n�+�	C�q8���W�Q
&Oe=�e����uz�D�n�����i����{�`j��e���^_=�7$���`wkm��q�#tI������`{)�����l$��8�l5[:R� �"#��#�9ך���V:�U��3]���꥙��^u$r�7�)�Qul��X���j�e�ٰ=^�5rM;.�ePlhi�ԤT��\���`s�5XslDD.�{)��9��ت#�\�H�Uv��q`7+ ާ:�X��!$ԥ�$L�E`j��`s���'T� ާ��h�
���!q���V���y����URՙ����&�5D�9P�7�"�7�ŀDܬz�X��	QV�w�\I�x��k�Ѭ"i��������,�`���t��>lM�Tl�|�~u8����oS� �R,�zUUz0Q�JF�+Vf��y��޽�`s�5X�z�ujDGG`oS� �R,z�XM��	�B��MSn�"�D�7�uX��V��v���ro���t�|��T�I9+ ާ9X�8�����`��L�uY�F)�oA����M�j��BR����RU*�JYn8�Ӏ�vD�\i���y���mq�֢�,ݱ�'�g���ŔB��La5kly1"/c7!X#�1�A�^��\vZ����qe���8:5�3��n..�s�ᮻFԂ�Ǫ�;2X�v�E����ٻb<���y�ۜt��!���6�=��#[���=����ҋ��`�U�rǙLq��J,��r����m�A�v$�֧ZܼX���A�G�m�>��U`���"�+ ާ��h�_�H�!�G`s�5X���u�Ws]�����J��9P�5u��7�ŀE�V�N, ��)���&�p���^j�5w5���V����[n���RR7D�X���7�ŀE�V�N,#����ā�Q�[��Ӻ�z�NL�8�f�e�1�+�%ݮ���x��L�i����}������BK�8��q��Sn�"�F�`j�k������@|�nky��rN_=�7!������t���訧)$����^j�"nV��]%`�R��T�N8*�E`j��`s�4�5wu���V�m҈�)ԌRȤv;�Jq`����+ o�z*J˶��:�M�1�ճ۞YW����ǆk��ՃM�
뷬g��P���m��6�ϫ� ާ �IOڃ�B�#�Jz�S��69�X]� ��c�9ݚXך��Ե�m8�%t�����u`w��Yq�
H�IBT�t�lc�V;O���&�Q8�r;�ɥ��X����lDD��ڰ6q֕CCT۩H�Q�Vu��y�����`s��Vu��~pH�$�:��/=Oh��]��g�
��v9q��P�z�y�X'�>l� $�Ȭu�w]�������`qn-�P�r��H"9��IX�`)ŀoS� q��H�"RI#�9ך��M,���]ǾV��������J���P
�M��e��V9�2|�XZQ	V)���۹$�ŷ��]a32eں� ާ �IX�8��ၿ����~�qs��f^VB�'n�}�lS�s=�Rg3�q�SR��"̪����y]���+ ާ��0�q`�<Z:R�ۑ5"��v:�U��ˆ�N,�����*�E*�z�j�`� ާ �IX�H����}H��bWWv`������啕��	%9���2tf�e5�|�ߑuv��J�7�E�tw�=��I��"��1#��*B��$2P��Õx@�H�YA+
��nS"�	��F0�d�
x�Gf�M$#7�& @�	 dA�¤ I�#$��cYB���� ��!	$�r�`H�d� i�����!EH�� ��� �X�D�1	Stv�DaJ��B�Bҥ��Z�4� е
ԭoY Fl,�HZ,�dX#2�D���S�!$�$)�HM400j�E�LM��{��vݽ�����]@J��U@��m��   �` 9$��jm�����倶���ӖF���k�j�5�5gJ�Y�@��طQ����vYTH��T܋hv�C$x$��*�>|����l��LK:����� [@  � � [@ #mm�    m�      �	 ����_�y��X���J��06|l�a��uƕ맗WbĜ%[�E����.�r�pln�� V���s�ɬ��7k�ۺ�1��m�ۀ95�%̴���ƭ*�[R��\�UZ<1Y��a�*� 4��f)P�̽p�	�5v\b��9���B�P�k�;���[���Wd�4�m��7u.�y3�͜t<WOgq�q���Uͭi�u��Rl&Lit�*1_�����)XyD���W#�a����]��,�v��n�r��qss�"�l�C�E��"D�F�|+=�\5<�`����Q��7���=��M�I�� 6�ͅ��]䃋���ۘ�l�*h�ێL�����uk͌�ƶwl$�z�n��Q鱚�ާv:m�W�76���۞D ��[�����ͻa�Ÿ�n��:��:�M]�5s���l��-З*����
b��
�X�%b�%�|	�f���Ɛ�����j��e^�:��*�����bSk�g��Wb���X��{m��\<��sA6��Ȃ�m����<����Kk�[kv¹4�q���a�p�Pܝ('6pՔ�,���� m�f�Jۦ��N.���c �mU*�&��p��e�{	���m=��)ҹJ2�ʫ��{(cRʮ�iwj�X��6q�7D�R��N�x�qX+���u���$����pe=X�w����=���F��t��\�H�"c5��b݌������m�zܗN�vNnX�ˎŷ[X���Ȏ���b��zO<�h�������X�^�� t��CH�����{�\��&����kXuZ�d�u�]�K���V���@j�i�`A��W)�u��ٍ��|��-��ݻ��t��u�z��*$�.�p'�דs��+�Rd��^��3kSӼq�.3�)����mf�F��l��r�i���@�p"6@
P�����s�|��7<��Q͎y�:�����v�m��ݣI���H십�q��7Q�i�[Cc�0#�br����������9����)�,qێ��c���uetB�q�QQ�)	�ӮeΫ�2P+ �)�XGp�;�ŀ5�VDԠƨ�7!@�Vw&�z�U������^��Im:5��M�ȣ� � �IX�H���k��t���)(��X���u���K�y���G�GJQr!��>r����腚�N��Of���ua���*|Xj����nyW�j�ntu�-�b�*�{5˞���ȓa��E�qryɰ<�=��6O�������+�5���G�Q%��;ך��7V}Ḿ�e�P�L�e��9G�H�9��=�`s�uXܚXܚX��J"Ta##��rG`g���<�<��.�v�͓�35D�ԅqXܚXܚX�����V7ʷ�u��(�T���8�m�r�m��Fۯg:!+���Y�6����Q5���8XܚX�����Vw&�1�m�֓�RQ(
B�k���H���tw�����=~)Dmʈr:NG`n?yXܛ74H���a,	�P��d(�D�L�� bQ
�j��&�w]��q֧Im2S*TR+��`� k���H����~h�"%Q���K�W�Z��|q���޽�`s3h)[��$&��"'=\��֌O�=;�#7G���=��狷웩Ar������ՙ��μ�`o^j�9�4�;ܕ�D��FGQH�����'T� ��M��'j&�b�)�⠒+z�U��ɥ�����μ�`nSK]h��T�c�O96^q��c�=X��У���P���4�P�~�\��I���f:Z�㔔J��5w5������V7&�V=�R�"#RH���@�mv�Te!���l��|%���K�Z��6T(�4��*!��9�����޼�`sri`j�k��U��m2S*Qx�q`� ����r����~h�"%I���ɥ�����}�W�j��=�|�#q��D���EJ��.r����"�+ ��vJ�"Ta#��r9#�1w5����nM,]�v�|�3tI���$��*�mYWS�t���AI��[�E��@j�U�����v�%�nm{�p����Y_c��+a�e啶���	�T8�O�!�ֶ�xö��<�n�|6κ:�b�(�dƻq
H�d�cA�{Y��ֻj�̷�7��`�n�)gkr���k�[����8N��hܝ�e�9�����!A���Zjhs�kG&�/;������۠f���7&�ZR�ݪ9�ڣ�d{��x8Lu:���g�^֡�:���''��*"��,�;��KWs_꯾���7�X�iy���Chp����2�B�6q�X)��}��e�h�m�)(�!`j�k�3�5X���nM,�ף��6�D9'#�3�5X���nM,=_W��7������b@�L�ʔG�����؈P����8���c� �eD�K�۫m��<�\u�K��9��^��C�o����|����ȼ^M�@$��m�����"�+ k��u8�Du��sDr�j�Y��'��~��D �O���xC\�`���6;����*0����G`b�k�7�5Y�朗�x�<�|��j�����*Q]�:�X�p�"�+ k��:ik�U1@C�R+��K����5f��ך��<��2H��)$L\]���q�r��U��;h�Q�n�g�݁�192��#M�RnGID�)Ws]����u8���k�E^��������Wu�5�V:�X�p�"���q֧Icj|�Dq�ך�}�qB$II	I!$��0�"�㺰�u`9�R����IA����ɥ��������`o^j�8�Xm��jR��c�bI�=���Of���2�ߪ����R�G��:����GlQm��Wm�����dR�r�vힽ]N�N	�:�v�N�B:��$|Vo���y������A��`{<���JnH�E#�7�ŀlw.r����#�%+�+�e+��lw.r����7�5X�kLu����Q(
B���V �IX�q`q��{�y(��7S��&9QGM��]�v����`s���|�+�j�B��Z��r�WOc2��"�:{;��x��㦮�Ѡ�\�u�9�%G`o^j�;�4�"�+ k��.u�>�}j�+T����tw.r��J�'T� �n=��u)|㨩GVf�w]��{�������r�6�TtI�%U]`t��N���0���N�&���JSrEJ'��{����� ��X]%`���r���UT]2�W�.�rp==�@Da�ᇴݵX��Ue}P� �^h%�:^�/u���gV�o]�H���u��ƛ�[��&F2s�Jw��ɻ�5�m��7��Y�l���S��.Mtg�4e����<����	Kl�v�ņ���:��4����(��9�^����ȖD�c-vޟ��d�;O$��T�.�d�m�֝=������wO�!N�w.$�<z���wF�)g�����u��[H��[xN���o�(��84���,X�`t��N���J�����±X+� ��X]%`�E�tw���_$n��'Q�)�rJnG`j�y��E�tw&�`G^�BAT2B�(r;z�U��ɥ��3]�������t���E(�qXܚ`7+ k��uH��*�W����]Ta�[�n7U��X$LH��ʺt���J�]!u���&�q�A6�m�T��Z�`����`���<��4������쯾����z�U��ɥ��3]���MQ����䊔N� �R,��`7+ }R,?Tˤ�TW �S\	�U��!DNk�,[�vu�Ww]�Ś��nI)U
�]�t��T� ������m��۾�{�=�H%(�Y��:�ޭl�)t��.��ݸ��ŀ�np�==�7Z*�uwX�`�E�wS� ��Wqֶ$���JjE`o^�;�ŀE�V�R,.��>+޵h6�;ך�]�vw�UUb��D�bB�3+����p#4�C3ݺf��Ɖk%��YP�!�� V�HD�����(��h�BB�����X$J֧����'�
1O �Ǟji6�E�@�,F�&kzM��²@�� \i�bs���$�� ��L�5��1�W��.h�kB)
�++)+��0`A���bH�F��E���R�R5e	H%KRL�4d,�y���>$'#l�*�!+,a)Lo��J�Å_)��X������
��� #�b1!&��sd7@�&�a��H����3��|B#%$%a@�`�)H0�h��Ȇ��� Dăh@���&�| �P��T�E~QG�OQU ��*�Q��y\���76�yM
u)|Ԃ#�X���u�Ws]�޼�`s�QDDu�8Fӎ��jE�E�V�N,.r��QW�(����-99�pvK�#�`z������1��6=c=Fb\㋖��1�m�s��wS� ���z�X�%*�:N���vz�U������^�5w5�Y�1�$䎓b��+.r��`s��wS� n����D���#D�;�{�����`w�߮���"�� �Ȅ���I��(B�~�nI��kbCM2B�)�������^j��X�76�BOy�*�b�L���z��F���:ȗC]Cۅ�6�ͱ�հ�p�i�*bQ�|�TQ#�|1����啕Ԕ.�l�ڰ2Mu�%���H"9������^�5w5���W���G�����Iԍ'��_�,.r��q`s��F�q]P�JRrEHn+Ws]�޼�`j�k�9׺�ѥ�D�t�'8��q`s��oT� ����{�����`�� �uW\���;f1 ��շCz��γ��e�����R��|R��nn�.'e.$�z7w0)r��2G���+�=�ònt݈�S+������n��(۲�v{q^i�e�.��oGF�mJ2�7��<�
q��5pu�X��/j[���w��lۧ%��B���q��{�v;o6�M��u��^�Om������(ꎹn1g�]��on,�N�;RB�2��n�O;F�t��C
r7s�e��+�1BF�$�'$t�r��ΩIXs���R*�׋J�֋��]]��R,.���3�M�`j�:�Ć�d�*SR+Ww]���{ ��X�H���'ʽ�V�@����3�M��7�E�E�;��{@�K�#�`j�k�5t��E�V��{ �����z���+��s\���.^���-�杝f����$X����4J%(�)�n;����s�u`{��}��{V�'6yT*��sZ�.\�nI���uSjŋ1 � �`��#b�
�����j��V9�;>n�2�]jT"F���9�޼�`j�k�8�����V#Z�BNH��Q)"�"nV���uH��q`ґ:����$u�����7�uX��V��vv�St��A(��I����xW�(5�f��h����s�J=7=�(�=6$��eJ��޽�`w�5X�5�]�v��F��TQP(�7��N,&�`�J�'T� �GR�#�_E ��V��vw]����c0#�`HF$�d �dFT	>�7U���U���Dm�u�p�����u`?Ss`{Վl5%;M�X�'�l���jH�N;z�U�޼�`DܬWIXƾ^��U��J�{ڧ��x�նqsf��m�n���q�O=�s���b�D��R4!ӃN+�y��ՙ�����7�uXX�k]	9#M6�RE`j��~���ꤎ�����~�;ך��$n��'Q��$u����V:�Xu8����Eν*�����C��׺���Vf����*Ŏ�H!�EHR�+�@ �@Q�y��䝾��w�ꢊ�)Bn+�y��ՙ�����7�uX�ڥn�n� ��*4�����)d�>���l�v�-���ă��.��v�����V��vw]������^j�9ܨ��RP�F�q��5t��E�V�N,&�`�\Q���A�#M8�]�vz�U��3]����`wF���#B8�a�DD�q���{6g�Ձ��u`qb5����4�n5$V5��������`w�5X�4I6�7*Hގ�Σ62v�`�"E;�U���*U�P�j��L���/]�Ѯ7�in�d�s�!)��c���]�	w]�5ƭ�r�š��
TR�dzL�Jd�v����K���A�yN#d�����%�k�GOs���9�Õ݄��/c乱�Q���]�Yc�&M�ok3�:�ϸ󂓄�q��۱k>;Z�o.��݃��������w��s��%�Z����lM�Tt��"j�='�G�`���O��eH�dT��:����$l�+�=�`b�k�;ך�k�V�͔��L�eJ*����;�ŀl�����Xoɇć�T���޼�`s^j�8���]�vQ���#�"��2>rl>J������ݫ'�������TF�)*�����Vw]��9X&�`)ŀt���b] ��t΂���9cm%�N0`�%�����e5
ujј�8�T��ͷ߯���97+ ��X�%`RR�'�Ƅ�䤤VVf�*�����u�S��	)ŀjh�����RUWWwu�IN,S��	)ŀrnV��[��7*2H�$V��睊u��y���`n��`j�=c# r;u�����|���������*ZH�T�D�F�>f��ınw^1�^�v$���|ݟ�6��v)� �ɇć�T����b��7^j�8���ך��q��"�)DI�%8�\�`G+ �ܬs��x��HHڎSn+�3]��s]����Ѐ��@0'�Z�7$����&�"j���IjG`j��`qfJ�$���X��B��"��»�Sr�	)ŀjnVr�������{N�;�*��k�a��w��Yy�N�1'��ֹ�d�9��ܘ��]�-�������t���XQ��57*��Z�uSnSqH�QE`qfk�"�V��X�j,#�����z����� �9X��`���Y��Z�ߓ��J���,�vr���;9��91�BD��HR��.h�:bHh!�i�JBD�!ѬȄ�Ma�ma! !.�J�P��_T޾�����(��K�Z,*�t��Sr�Q��5fk�7�*U����H��R��B=�Om���p��y�)����4���}��uѮ�HH�#N;�3]�չ�����`s�v�"j��T��&�ve��B��ӏj��ݫ��uz����#�ט��(�b��#�:�|�t��W9X(�`�)(	Uݶ������5��.��s]���u����{Σ��G�H�O�Ձ�Q�׵�2^� ����J
��?�
(*�PU�TPUh����J�
���(*��PU� E���B$�P�BP�U��P����P��P�T �EBAP��T B
�P�0T ,EB"T"�B0�AP���DT �B�B"�P���B
@T"�T EB*�T  @T �B
0 �P�1!B @T �P��P��P�T"0�EB AP�#B �(�$��P�"�*!P�+B ��T"�P�1T",B"P���P�B "@T P�B"$B!P����P����B �P�+P�P�+P��P� @T  �B�P��P��P��P��P��P�P�)P��EB � B B"�EB �B(0DX�
��B�P��DX�$B",B*$Q*��T"�E��EB�Ab�P�* �
(*��*(*�򨠪�QAU��
�EW�_�TPU�QAU��EW��_����������b��L��@8�j|� � ������!����s�,b��(���>ا@5#A�}π    b _f)Ul�@ @A)B@"�J7|i@[��������СFp�y4(P��n
xzy���^� ����F��z� {J ��󞷀�u��{j�m�ո+Ѡ�9�w���`��և��pk��::�y��zi��^�<��HR��ܪ���� w` �v� 9�w`>� ��� ��7�}R�w`��<{xu��)�F���
��(���% �/
��t9��^��t=;�q�MB���½i��l==zC����}%6�v�OM�纷���
8�k�O>��Mz���GB����á���MtP%@ @��@�4)*HQ�L d��a4�?Ǫ��ʥ4� CM  ت�MO�D h  0�  S�j�OE* d  ��   �����1�#��&�����L�(�� h   h �t�8:��̻{��h�TE�ݖ�;��H���'�� 'Q�TP%D\�������DQCb.?g��?�7����29r8���w�=?�����?N{,}�6t�ѯ9���?.OU�CHR*�� Q3å��\����'���("��S?��SbH4~��˯�+�vWJ �e��":���Υ��ç����,��������N�Mt����݌��C��q�p,�0�Ç�����cbÄ�ap�p��abp����2��Äal�!��XF�-aD�����6rrs���Uq@G�����"@ �QOAT�UK�����a��ʇ�������Ϛ}�������ρ����6y����Q�������5�,�#��g~�����uӋӁ��^o��-��0�pN��tr�/�q?A/3�;�ב���wĠy��f/����n��!Va�R�Wь����.�#�D#ɯQ���,!��P�����H��=��/�pT<WR�peP��aE�˝�x2�����$Pٖ���d&��U�@95G$��HY �ֆ-6�J� \�
�ڲ@h�tZ/�����O: ќ�I9!�]�>k���� 02��Ho��I�������Q66�� &��v�C��%ÁgHK@`(�#>��#�B��R��8q���j`�\T�#k�7e�D�.KRh>	I�R�9|�Z�� i���`v����o��1H��R`N)�`2R-�&��bHU%�@��D�h�*`�Z�,
.G��4^��_����;�5�fs(��|`»�3[�>�v�����l�t����d�Wf�&og9�6B��J.�X�0����Qd���i� �X��h�%�g
�� Pq!�g!�;������5�Z�A���sF�9g�'t���Qi�fa$��`�V�K08H� �i�XU��;fjW��~�䰽JU�Nv�=��HfN����iSs�"ŃH �'��@�;N���>s�o��<yi�_<L+�O��}~�&b���ˡ�D*�\�扜wW��J>4pH��h>�ԨA=�er�����N��tJ�崙��*�Nw���tQ�Y����c�"��
K$!0�r�/���KBV�j����臀�=�I�)�C)s��!�-�g+58RB��^�{>2��M�4�t(��B@)���P��4HB�1@S�Y�[����A}����y��X��*���ޥa���!�����f4���h%�I
�ؽz,�R�Ԙ�MoO;����bH!P6��B 勠S]����:!ܬ&�Ұ����Z>8/�녭0����8��C��
�!L�
�Vk9��K��ʲ\kp�QѠE�<j�q�f7��(���=���ϸQ��f��i�l��x%2��:4�Xc�C�XI�,3�ш6���Q��(�y��8���1I����4#b`ġX�04�o\��
�nV���C���P��%�2��a�`B>������\ѭ�sS2�����B���E�������a��F���n�n��#
.��ӶoY4�fa�����ed���*�C�_C������}^�E!��Hd*��I)�R������<�Wۧ#+�L,w�e
�;�Z� �F�^�� �
�ys�P_`>'�#1�t@�<�r�[�4�Ѕ�V����f�>|`dH @�-1��ą4�Ǧ�^������H[�l]w. 0Hm)v��aUT^Z#JI$�Ki�o�������Kc��a�|s�H1��#��>xu�
[6�|s�*�����TB��eᣧ�'�Ƃ�[�}�A�C
:���<o������z�x_���啉
�,�[fh�6r|�^� J�0�����o5���}���߷���6� :;�q��9��b��t(�����~><��ζb�������g9�o�s�/��&�j	(�Mn��+�r���3,�X��Y��ٷ$���9r�;��=q���!�o0GGI�����4���r�\x�:^�341߳�����N�L�3m �8       m�`H���p� I  [@   ��� h    m -�                                                          �x                                                                             <                                                            v�2m�m q��WV��a�;#,E�Ŵ�m���*V�ZR�і��Ec��Yxb���8:���6er�Q�Y�Wa�ƥ��a����ٖ� h��� 	  �ͳv�m�  -�l��[V��(<.� ��  �&����D�6�  �����-�                     Z�����Py��X)v�!���p Y(
+�Z��Nj�ٶ-�� �d;`�bE���m�O���κ��Ϲs�m�U ���d�2��Q�"U���U[)�*!#�Z��]1�� m�m�� �n���U�t��c��U��H 8b��m�UW<����mE	5�;m�Y��tK��f�&t��h�a�nS7[��|�\�U�*�<�PIL��i6m�`۬쬚������^���jU�r��3���kX$8��d��n�� �f��^�����]c�h��m)��  z�9%��rlMɮ��i�M� -��!�[S�C��Ht:�)P��jڝ'�V[�ӗ-E=v�U�áU	���$/|�x�!��z�I,z^���P����5��m 9!! m���Q��fs��UU)293���-��e�-��T�v�T��#�x:�;8ت��nM��ayg������[���v�B.���:j��!VN��kF��NJ�
�8� ��2q���snYj��ѧ��<vʣ�#b�imK֙�2��p�j�8꧘�vbÎzغ���v� s�
U���Y[��jFx �<K�h}F���G Ǣ�d�^�
�K�ԫ[U*�mP
�-�d��   �0m�m��װ  hh�[gGLȲ�� I# H� � m��.Z����h��K��x�V�9i�bImr��j�]�i�qDgR�+��݈[<0�o���@J��]e�ݔ��;	u��
�u�.�`-�:��tA�JBC,�VԒ�׷yy'���`���^�� ή�nj�`�^e=.�gBܭ�p�+�I���m����2lm�m� �$�m�������.
mTەv7��3��I�k�a�����l�5�B��%�,�m  q'ܗ-I���� S]cpUV6�4jj�͈��=KR�r�.:�cv��N��vֽh�N���n 8��6np p8p6� �MC��jܵ� VY��`�dq�����`m��[�.� ;I� 6�����9,�[kj�&^BM��$�����WL�ԩ�����,�X�ʭ&փ�p{q�lΠ�8{%�nλ��o�e�趀݆�$�J���:j���S���P�V�vH�� �/�������[n��ڐH �d�zrݖv뱶Ŵ �  �J��"��: u���I�n�s 6�SZީm�tQ����;�)T�g��)s�"
��l2�n5a��g�6�8����./^�  m�2�U]UZR������[B�k�bI�u��e5�I���l
�n������ z�z	m:`\�l]m��2�<�v�iթ��7���� ��;6ݽY���z�EU ywrh{uƠ��{�����O�sho�TNa��bz���?���x���s�yrx��ݻuݫm]��ff_���=�Ο/{��������ݻ���Iffffe����J�,�v ��iF��6�Qx*`�^:ڷ`:�"Z���u��;�gD8*X�	`Qx	���BILI16h)��Ȝ�� a� Y��`dPJgQ~� Բ��
w��ĊH6�!Y�d
(�:(�Q5b�Q��<�&�(Z�pD(��:�]�P>�ˠv6�R�� �/�;4/���}ث�M�t��+��� �q��
\V�߱A�	����xu:!�V)�P� =�I	!Gj�V!��h�Q����%��]qN��M`���ZS�@���Ч���-G�T^+1�D+�� � 1Z7�_E9�l�/{{@�DO��D�s��n��DE�&�j��� `=�#!ŖLX��E����#���J@9�W7��-��g�PM%uH��bs���ےI$�/Z�[m�$��           �               m�           k[v��`��"]3�mrG@M��u����m�[�m��70�     ���F�-���z4�΀��Ly�n�y��n�� )p%.��gomlo;@�q�셕�ݫ\[�)T�%ܻH`l�7d4�
�n5�pT �8�'&xE����S#�Lgk��(��fX����H��ƹٞ���V���n[��%�*�	��	�ݩ�q�y!SqdlHm�rB��vb�+�cWP�Ů���R�C�;��gC�8�)x����:���j�M�4��d�;�R�]��ymv����*JVף�L����q7. ��u��k�M7\�ś�l���j#�B�e�1�%*iRgc9�9M�sR�������nt�yȮјW�e ��[�� 缋�6{��p> (v�w@�/��ƍ�ߑn)�I$�m�  m� 
Z$�cQ�<f}i�WCɕ�hx�]�d��o]j���,�c;�d�v�\#d������e��u��E�|�
�P��Ͷ�)��-L&�-���I�&��4?��n�P��ʯ�8ۊW��1�u��F[���0�ޭ���bs�)8��w�u���иfu�\��޶0��3/|{��mkI�е�R�Q(K�%N4[�e� f!��^Σ�)�J��>ݪ�<�
��q�Gu׷]C��f1	ޱ�Ubչ�4��t�#<�h��|8k�1S�9�qJ��<@�C3_OVd�I!JAQ��Ɋ�⹚�c�a3��z�����f;#1�9��n�b�]fc@���h�
���^����*�@�b�'�p��У���h"7P�U��=���� w�]���\��1�$�	��
�c��kY9h��2ȳ�Ufc@�g,�#<ha��0���,�d��+3� �3K�Fy��\@�P�C�8+�e�{��1|��
N6!�w��1� ?_�I$�4�"(�F���\�?Y���L�l��痝����'��R�1�37k�_z�S���d�1v��O/#1���V}�Y1����[���u��fo��~ޞ�����u�{�       �\�Vܔ�$UAl�t)�5��-���T�'nqu��ۨ��91��e0Qk�<�K���Q��#��^�ܜ�޻��ڪ���،a��R�28�D9#p��q��3]���E���\F�
#�C1Vf19�)8��ǽT�9����pz�w�b�v����E�T��c��.�z�C��~`	YuH�9˯,����	���2�%pY�B�Uݺ����^�j�솆@�$��!J*�/烥,�S�v�;��e�Fx3{�xp���8G2F2�1��3�U=`�󉸸,�#@�cuV]k� s6�ե�fF��r�`a�"	�1qVf1f�3ÖXlĸ.�w�b�h����n+3����
9�`�X&�Dㄮ��=�j���^�c����U��Y�8���9�a	{9�.�l�N�n@�.�g��FТ3ʳON�2�u�ޠ3v����q� .�v���'3A'!�*��3��Wk:���a���>����.[/$�%h�Ύ���ˮޜ�iŵ#E�T��c��.�v��l�!+���X�A�v���3�;�YxŐ<�9i��ڡU����kª��U�zu�2�5��3�ۥ������8�      m�Y�7Vtmb��e�{v­����a�M�	�id.cPrl��6vs<8h��hm(�D�u��+��<b�d����`��Zs�J�T����o-�K��h�F�9�3U]��� �����*�R��c`��p]��|��h{x�4[�A�bլYu�]���)�J�:�ګ�c9��$�H#t����.L�ٮJ������C�U��Y�|�9i��L�p
 �tU!w�0��W�-��I��1�Vq!v����q�Y�C3fc��NF@�C�U��Y��9rI$���M���ln�l��D��\j��1d�=�O-¥fc f!v����z��)�J���]�������Ͽ����K~&����D �BLL�+P+V7L�jR��S.P�}(���9JФ��yxp�pU��L�%�6���Xml�,�ohB�XQl���q�l�a,�1c��L���m'��o[ֳ�6jxD�T��w�}��_��4)�J�]��T;�
}���W�+v����G�$o{�Os�Q��u�ߖb���i�3�[�*��y�s��f|���I$Q(�����+�q�cX[Q�{��^y�U�u�x�q��;�w{����RF~�N{��9���n%ᘻ�fn�}� @ s��
�����{��[�����=���uzI$�%R����e8B�D�h�aV��)�J����A������3���{ws|2�Sr��{��f�{�Ȥ>��ovz�^;�y}�+}�{���Ⱥ��,)��y��h�1�       [�4k�lU$���o�ݏ��:�� c�9��Ɲs;�î�#7[D]N9䎊^K�rP�	c�m-�e�1D.B̾���9��^��߭� [/Q�*J]��e)lG �)#?wy�,Ϻ7`��E���Ή��P��/z�� \��_�fN9���_�5-9������}��� n��}��'5�rI$�GQpѫ���ln��,�O;�<����t�E!��}� EP&�$��hR�I('�sQ^����P=��!8ێ�{�1ϰb
H��un�f9��.Ds9��������$�D�iHQEue�r�	Rb���W��I}���wFb�X#�\d�υV�c�Ӿ��ј�\���̿nڠ��C�[��C��n@��+����vX� n���nE!�>���P�Y� ���$�HR�En6,�ҁGQ($�8�n<�w2����a9���ww3�sq��G3������\֋�#����wx �S���{e9	Y���xs�h��l��I
�"�Y�x30���R��u�N���^��3/���܁�f}N��������nE!���oU��سA�q�w���T=��w���rr/��wv�P�%ߓQ�       	fk+c:��� ��x\F��<�����h��W��uk�-3)��;��F���vn2���[�˃M/wEA��t������'�Z���ٹN�r�쮺;w�x���D�Eȏ=��~��w'Wu��F����n���>�9	Y���f���y���3���̶g0� ~�C��fg�/�~�| �Uv�N&kiѰdq�q�H�;�}������I��^��Q��P�� � 9S�@�P��|�N{�B�s�:�r3��	�����:�A�GcE�|�F�#�Ǯ�n�������r��ݘxZȄ@�C����� J˩ms���I���<�N	��+u� �P�a���ј��~C����C���ǧ����Krj�C���(W�{�|k�?Y��E!����r�z�ƣ[�����cMIW�~���n������9$��B幜���g���L�����Z�s�^�~ �6gpz4\����;�<s�!�]֋�.�n��Ӥ��sxS���b�Ť%�\�h* �!.��^F�zodf87�Lnk�f6>ګ���$�Dds�XY��U���{z3Ѵ����y�[���/>;⤒�x�!��~B�y'1�y�Ǎ@s��\������	ŧw]f �����D�>��]���qi�$1U��>ƹ��>�r�Sn����V\�#����˺�a.�r��K�W.Q,���H�&ٗ��zBl)K2D��/2U����%�D�>�A#@"j�M�h�a�IAv�>�"J ]ZH����89�5�|&�\��F�� F!hB��Ca@F0(�aV%�����ߞ���$���7W�N�UUUT�\�[A ���۰                                       �l��;��n-��W4�c'm�`n�:\�	ѵV�r^a��    V�uT�b虸NLs!���M�۵�Q�[
��`���m6�\k2R��6��l#}����E�0��<[�8� �핎�{T+bA�.W!���)��lj��F#�sn�BY�cZ<na�s�2뇛��v�Y_0��@$��i3(	��y��3����vZ�����N�[lg�b����=��U�n4pP�����z��Y�n�rqp��+�0Y��.{��Nax�m�saYFb�G<)75�� a0g�c��n�U��:�T�SiK�E�6i݇���u�D
�(ˌ�ለ������{����W��n(���M 	��n�6DP4�Pڪ
���Q�g�       ��5�$���6R�![�s�=�Q�i��`�r�z���m����q[�$6,n�-��뗪Q�d�e�+�Yf����8�������ν�?��O׀��v�;W.��.ģ�$c�,9���u�Xt��uޢ��!JY��> f!���<=ϣ���*��'Gw]n�ڠxy�-��2��=�:�cV!��;j@�=w%m{�ZsU���'�I$�Q"-��%B\��Q��C�ƌu��z@�Xy�뻶V��g�H�E�*�X@J�J�-T>�� xY�'�G9�}���tU-��3�#h�Bw�X ~�1�	�t� \Cwe^!�i�СAn�w�E�NB���=�8G�Lκ�ՒI$���2�����̍خ�N�{�B�#���;�y�UVP�n�f�����y��V���Q"�}�2~�F�~?yH�<���bpNPC2�� ���+� �$P	�D+�~��o��yu2��
l �#O�*��!�����b�P�'�������_�r3��#�U � /A��uY��t-CQ�:䖺s�u^�0֮��Tw�o��s���p�P���Ź���|d_P5UA����`�����R�*�%VH{�n?�Z���=ݕ��o��$q8���C� E�
�{G������L?��Qq]�� �������ޗy��O~���0T���	���/�a�UZ��XF!��ې�����8�rû��q�#QR޲���rU�T�{��9������ R��?0����:�'ﾕ��'pz4\���P���r�P�T5�G>:=�nH_0�>n���Ƒ	9�}C篳�~�;X(       +r��N�\Zc<lZ���W�:�Tn��Ն����B��T����?j���;�vWX3qlƱ(��e
���Y��x� -�i��F��:��q����R8S��+������~�������q8t�B�#�CwC��y=-��ϻ�.��?����c���\ꉳ�B��ߥ{����@�L�gV�F;#��s��:�۲@[,�(�*Zm��4�Q�ުs�+�I������ڠ9�N��]K̨�o���R�(����[�CH�P��������-�W�ߝz�}UB* ?��,o4
r����Mf!��?U�����s���j����@{�n��{<�� Jͪ�Ѥ�!"�(ɅF�N(a�C��ϲ���ߒ��M����?�U� !�L�@�W��+�����MgEߺ#�  z��S��V$g��@�>`{�g�1�n��h��r"�@W}�H�Cf�� ����M��M��	R9[TG�p��]��ֆ��|��3|�Ҝ�)[�j���R5h"7P��t|(3����p>��}�!���P���5�Q�>���exhclA/W�lE�@��Cz�W��U�������:�d�uf�K|�UT�cZ�]�u��f�T~I����ygdI�wh7|��+J�3��|  ;�7u�b�P3�=.D@�A󽕘�H�c�[p�����r�P���n���^��)c�Q�}G�}oⱊ`T�bBh���U�Jǳ��E�?�s���H      T���1�RZ�·Z\s��l�ٌ.N.x��$彻V�ê3��G
'k]l�ͳ���\�.�Nεz�~���w�=�	Yfu�A���Sg��G���7G�{�o����=�Ÿ� n����~�_|���3~K�ȓG�wY���ڮٲ�fA�T>�@�Cª������<o��W⤌�`��]���1��_&��� 9�'�:خ�+�?���_��$��Z-��b�]}���D��:o���V�{�>��UՑB$��*�Iuv��I�@����'7g��o�A +^�/��2R�w6�
|��u�>ێ)\���P U
���C�c���:{�-�u��T �_+��1��\�I$�"��/:�&kiͺ�ڄ�y�>c����}@
CuU��l�������7P��\���RFx0��$6�
ewu�q$H$8�����O���z� �"ā�v�S�나�
Q�CE�Y��U�e]��5y+xE����(*�}A�8�|R+�!��P(����c,��Nf(Yd%�$� @��P�a7\������l��읎���{�~ڎ��6���W� 4��]3>
Y�L>Qu��N����� O��O�a_��o����yh��U w�7o3�5�xP��~:=�m¸>��G�Ɛ.�}�m�$����7X��0�Ǝ�>s�胧��
R�WH��P�|(t{�n��qHS��׏��g���P&�����S��>�w�~?|�~KOal�|*����}�.>�=�X+\*����\�e�+1���CwX
�����rI$�Gk��ƫj�R��qY�H��)#>��{����xYX��Ƌq*�1m�+��CH�㣿�+�=��k�/��=:��)J�C���ZMV��*�o~�)<;�31׭T4 ���޷������m����      ���M-� Ru)n݃v^��_��:��tl̳e#���x�bK��M�77=;zLvzr�R��D�C�[积]��w�[\4e�K��̐�+�o�E�U~�g:[���y�H��@W�X{g��pU|�����*�U����c2W�!�_�v럳�aRFx?W�~���?~��b��9�-Ă#u(|_�[�i��~�I$*8��m�ӮK��`��VVi�fau�Cڪ��_�C��܅)_�V��T��R������@�!��T*�1�~��E!|��������3�[�[�@e ��e�o�Y���[<��
��U^��u����������.��V������@T*6��Hc2W1�36������a�����|k���uv��?
���S��24[���s�c�UB��Y�� >��ۅpxU��}��C��,;h�
R��YB���fc�g>W$�I����k���/2VƮÆ����z�f=�Fb<�4、��{��7hY@ a��i�-��{��k���5U�һf@�T*�?�B��h�T�o�+e �ۻu��Ҿ���4v�(}�A��:�C���$�D��F�9I�ː��
���#��l�_Vu�{�{UT�����h�
��Ǥ^c@�_��~拐�+��%��;��:}�R��5�v��]f!��p .�����P�@>l�\,��n   �C�  M��#:�XFҰn�Uܬr��p�&z�G+ۉ�vZ��P���9��4l�p�b�6FL�5��r]����E�O< �Z)\T�]�R�ʠ�)���c�׸��~��n�:t��3%n��bv�UmR,��$��|t�z���1t���h���UxU?�^7���!��ߘ����n����+��> }�{Ͼ}�| [Z�Z�l���%�		�iHR��C�����g����!|��*�P�*pتT�������2f�uyx@]��u��P�_����> /�ǲ)?���k�-�g�?��d��C��.�z�翟 -�C�N�Mx�WM#)H�}UNqw�9#>9����03|���n$b�E�[�i食4]��l�����`0��#	I�R�Q7���
��e�۩y�R��:Fy�~[�����8�/��_ʨU�}��k1�$�mDTeH �,��r��s	<�λ��ݠ io��r)}���x��7V� �B������Dd��:@�B��_W;e�e��_����������Y�J�H�g�ZU�V =��Q�v��R�*�z����EUR��}�|@����I$�e�
\��]X��8�n����ha���\�)Wk��;#�>���7��dqH_�4��/��
���n�����?|���Y�o�U|����jG!�߾u�U{�D�!��w:T�I��;��"w�@?T�B2%���Y)�^�
ƪ�r�W�$q�����N��t��^�����s��v� �3��m ��                                       ��EkZ�K�܎���.���˦�m�K.)C�շ,3�V;p  
���8k�r9�1���)C���7$��#����$�Z4��LDQ�Q��x�VZ�����f�:wp:6�#r�c��Ty�n�a������3k�qt��,*�q&6�R�b#
V0���́*�m��6�B^�z%YnM5U�)*�/3�ԻZ�����`I�	��G=���'[F�3�-����6���`_+]�upX+�j�5��)��cy�i�/L�٠�3=���\�UAvx;y�
�y�Ġ]P��΅��9�ٛ�-���pғ��� =�4/3�n/Ji���nB��^NbN�U�j� ŀ��PL�Mi�X��� :ցB�?tO�j���K3.�333      
���i䥢	*�ᗝnm�E�ٲ\�f��YZ
�ҺWL��kXp���r�{<d�2෶{��ۭ�L˯f�^�{�|�z���H\M�db#8�sJ������ ;�+o�0��|@���Wk�߅?�k#E� ��;޺��,��X�0��p~  /�����}��~?�!����IK#�����s���$�晗0q�b���W�����8�/��z��|�Y�}^]����]��&
|��`H�`]�a����ʑP�x�y�}�;Ap��"��n��~�T� nۣ�J�09+u�.л�Wߗ��$g�w��>���}�{���� sm��M��M�p0�08�q��2��C�����@r	 ����I��s��w����H'�߳��
���\MD=e	 �'�Iq?N@�'����/2��BH$��R\A9E	#��@�^*h�a`4LE� �>P���R\A?w��H$��s��^Vd�&���,�$D��K�H'�߳��V�~�IpI�o����!�$D��.	 ��3�I���r���9r"�o�ڪ��f�ν��KNm�͖1<���$�{��A$N}IpI��@��=�K�H$�%}�/
�	 �'�IpI�$�H��%��
�w���1��'���z��˚M�$�$�H��%�$��قH$���\A;�W5u/&�lL��U���%�?U	�{0I�?z���kT���v�)}R	 �&}ü���V�pI�}�$�Hv3��@�OQBH$���\A9�A6}������.���9�no�u�7�w3$�В	"~�IpI�$�H��R\A;��	 �'�N�}���̗��A=E�`��5�>����	����$D��.) �Z�z�3hI�;�K�H'9��$r-D�i.	 ���(I�5^���yy�I�$��H E�>��`�	"}�K�H?@�e	 �'����	>��d���	 �'{IpI�$�H��%�$��`�	"E>G`j�I �'߀;�k�WYa@      Y��^S��Mz`2y�X�e8�ΰ�틭 2V,O���^&I��s��gt��h;7	��+�G:Ս��9�r��ri��I<�H#�1UH��Iϳ3330˪ɖ�ɩ*��nz���(�<�\�r	 ��A$M���/�����GT��$Oz���	�_j�^LВ	"{ԗG�()[�s>�A$Oz���	�$RD�k��YWy+I�$�{��A$N���H��{B=ώ�K�/ ? @>��R\A>�A$Oz����@ ��~�	 �'y>��/+2^�pI�T$�H`��ԙ�O߿f	"*'�IpI��oٙ�mzk1ae��n:�24Ue^fBH$���\A9�f	 �'{IpI�P��D�����̚M�$�{1t�|�D��7�D�A$Mv���	��A$Nv��"Tw��+�^VhI�=�K�H'(�$j'�ԗ�O{قH$��+��\�̚M�$�$�H��%�$��`�!�Q;�K�H&o��]K��4$�H��%�$ 9�f&�TD�i.	 ����I9>ӝu���UR�kWm�h�Վ�X���].�{��N@�ϗ��	"w�� �*	��A$Oz���	���s2K�	 �'�Ip� A��YBH$��R\A=�f	 �'w'=��3%�7�OQBHJM�0�@X�� ��($��"�fRX��fb"t���>T�&_��I�R\A2���^fR	 �D��K�H'�}�$�]R{~��$��>���I=�s꼼ɤ�A?{�`�	!��i2) ���$D��.	 �} !�������*J�
�ݻ���k��	��yy19 NQBH$��h>��N�s�I��_z��˚M�$����*��H�}IpI����H$��R\A=�VW$��hI�;�K�H'7ɘ$��'{IpI�$�H���~���Ui7�OwقH$���\A=E	"�4�����ʈ�PdP$P��4�d%�
���TE�Rv%A$J�%�$��c9rky<�y������K2�ŗL���3Պ)z�윁�P�	"s���Owف�D �=�K�H&�|�U�a	 �'�Ip���'�}�$�H��%�$�P�	"_�Oܫ�̚M�$��`�	"s�K�HH'��$D�i.	 �����L��ВH��'���O��$D��.	"���`�	"{���e�乤�A=E	"}��OR=�&��	���A$Oz�ӽt�����w�ߒ��|�       ��qwM[4vm�PN��y�Mus�͸v6�au8�`"B��Z�;t��5�qu`;SR)1���p�M�G^D�&�:���Ӳ}�����sˌ͚Z��Z��s[�dgS�A$N}IpI���$�H��!�I�$�H�ލ�ʻ�ZM�$��b�BPIޤ�$�~���Iޤ�$�}��z]��/4$�H��%�$�P�>�Q=�K�H'���$D���U�d�&�� ~�����}�%�$��`�!�TOz���	��*�y�CBH$��R\E9�f	 �'{Ip{��E	 ���<~�Ukk��ŌC%vYI	\ '��'��:EEݐQ �'>��$�z�A$N����	;��\ə��A$N���@w�(ꆀ��P�	"f�.	 ���$D�;_z��˚M�$�P�	 jn�.	 ����L�N����$��er]ea�$����%�$}��D�$��R\@�[BH$��~9�ʻ�ZM�$��قH$���ԙ�O�P�	#=�����9<��w�UV��T��;2���0N��/�uvo��I���2	 �QBH$��R\A=�f	 �'w'=�̺�&��5�$�H��%�$��`�	"{ԗ�L�n���d4$��j'{Ip������$�C�j�M�<Q��m�Ŧ�)TAq��fE�C�e	�e^����X����	̲Y	�"��!�\��2I,����L���/Zf�t�20!� ޵�5w�� ��d�JY��X�4�ܑ����lJ%he�0
�\.���>�g�����+���ک�"A@�:?���N�|"
��h�N"tM�'țSh0��~M�Z���\A=E	¨I9����&�pI�}�$�H�����	�)I�;�K�H��gg/+3+4$�H��%�$�P�	"w���N��9r'��{���ibƹ�lpʕ��4VxJy��=�cx��Ǩ�$D��.	 ��� $D�i.	 ��++����В	"w���������J�H��%�$]��P�	"~�~��^K�n	 ���I���%A=E	"����$�}���w3	y�$ߨ.'�ԗ�N�BH$���%�$	����KV�5��0Hk�9���d���=�7u�b��<rI$�(ˈ���c,�mr�'�_g���[�ae��q�x31ހ��@�U�t��$R��鯨�31�w��a���T>����[}��!��kŧu�F��{�;�=h��ɶ��ʜ*��P       lin��)ٷ[KB3�e�P�2���#��N8���M��3�:��]���dBc[�p����}nk�J�B�4F ��I>��%뾻U��;t���F[�������u��}�&�V9������=<�̀�WkO��fc�"�O�S����1�����<�Q���w�����ç�)��o d�0D�̒I$D�$�Yē�������H�]���P���u��ϘrFyg�g�P	��s�_�UQ�����S]-8�h)����0��G5��+���*Z��,>�̔[�v����n���?9$�B����� (ff:���̷��'}��o�B���!�R�`���=��f!�x��t��!���]�ў2��+'8p��$Phq3Nf:�j������K���1�P�>��$�Im�*�Ƭ�W1�3��M�v��ѫ���N���~c
X�:M¸31��@�Z�Xx[2��;�]�׸N��^^�� '�9�=�Y����&ʅ�����
N�~��=7�c��:G��4�uz��Գd�I�	��s�'R\O�kL�x31��ZG�TF�ӧ�)"�����b���|�ڃ/�
�wu��ަ�Zq������f!���c	�J���߾��>���hF0��Q4 @�T@��%��m'$�H      Q�q�s7jY�T�H��f�,s=�˸������.yo]��4vi�WRYq�����nmDl�>q,�J�S��g����o`�̼��p�=��Gu,f;gO�ӧ}��x���1��}+<M���0��s��u�b0�[��-w�}UZ�CH~?��<+ﾕ�CH��͞���U� 3��3	��I �6p�ZUL3F�Y�����S�N��3]���h�uA�< �F�M��@ɣ��n���������f@\b f!����{z�p. w�^uv�`�˒I$JTm��Q4���E�M�*֎G{���,��u��hio��n)�|�Ck����ו����F��b���B*@1Ep��~������q|\���<G����A�"
8�hhWn������Ύ�~�I$)C)�B\�J'T�y:���uv��ȻC��vXf@\�Z�@����f?���>ߓ�����uv�<�6�`�v�:z������_�l���8�<�:]�@�A����I$�(���ڷf���]��r���E*��.л�W�^X\��#h���u���0Dq�.Н����CM�	�W�}�ҳ�_�/���Y�;������SG��� �����s_��n�� ����)� ��@��@^)G��&1���8�$��1���,>$��)�M�Y(V��|B�*�i �U|��y��"لbp,�3P�!6"��)aC(�(xC+�k�������­UUR�*�m ��                                      �M�kB�F�^^�:�<U[*�ҩ�`f`Z�j���7`��   T�ηE���	h���1ݥ�^q�4pTi�g�-��N�q��)�#i1*���(��R��\"N�w6���-!uN.�Hb���Q�+O!��g���Y�ns����L�Nѝ��'��mrS�9IH�{n�<���Θ���Rĩ*N�WK���#�'p���J��m��"��7 A�]% #i·L3�49���:7h�W�x�y�ePwj�qԕ�k]����s�m.Z̕C�dV�l�k���<����4vHq�V۹b<�8Z��-`7"m� ���ѥn�/2�����޷�UWz)�)��� ߇�
D4?P�D��Er��]�Y�P       �5���M�����RCr��[��M��c��M��"v�7uy�&w\�l۹w,���l^���$"�+W'U�b�L�O{�|���޻�s���j�mwc���A#�"��S���|@�P�c���J܌��C����oP�?�$��8���~�a�|j�W������:@�C�m/����#<@��c��>���e�)͹�jk�Z��Q8�#��b�u���7�;�U�J��z�M��*�8W ���1��`vXr�]��@f!�̕8Os���@`c�<�Wh| w�c��b�]f!d��N�I$�D�1⠆J쫴b�@�����u���*���|�~?p(╖�Hh]�7$g����T��T�(� Q�Ou����1Ȫ� ��y�bC�֋p����W�ǵ���qj -�i-au5�֐�D&,9JV� ]�wn��{z�p.#�@�!���fq,r0@�C��@
9�a��58����]�@"����:S��˾ӮN��V^�>�p3�cg]e߭L�I$H�Q��B2d�)\�Q�iujeq�쓮���߷��9�#��;κ�B���0wZ-���m5�1凅��-��B.��(fd���&�'�H����Y�� hѢH*��>Re�$�  �   ��0tgMr�a���X�@�>�pA�ł�ך��ٳ[�ƙ4N��5q��a凒�.nKr���'�l�G}��YUT��,���9��G^mjT��u�>cf���n��� ���tۊ8�n��_�C3n�խ.I"��Vj���Y�9�j��!�n��}�'��d�I"J4�"&�ڠ��6f�s��֦ͽ�~�׭ ]�����%J�\�u+�j���
��Am��a ��Y��(, cC��u}'�����:����Y�31�  e�;�W�b�ޑ���3��C�\I,� �.���$�3KN�-C����R��3�]�\��8S�� N!����s�l��w�*�R6�T)��F���y,LEw�,����h���76U�@�C�|�!�42�����^:���I"�sL˘(����Q҄�8�\@�P���@Cu�k�@F�sF?Z��a��58���dz�8@�Uxp��R�ht�v��΄((Y��vѲ���aq�uv���UUt�5Yr\<��sߊ���a��q��>��b@ك��n%����ha����T��;h]�׺Oo���u�c㘄<��$���Bw����4�塋��čI$�      +r�1�S6�jvk�cS�x��(��5sZ�+��-sؼZ�e���]p���sW;VxA�=G���rV��,�1=���k�	�]�2�$\l,��kE�ntz�^}nw�a�Uٳ��J�C��.��C��MirFy��@�P�>u���,%�.��z��X�����\��ֆÙy�g��	YaZ:4I]�sB�m�!a�n����u����3
��o� ��U�����0��\�@@�C���,�ߴ�A�'f1Þ�f:�#<�r)Y�t�������ϟ$���4�d΅l�tN"i@�mS��� N!����O���R6�>\���Ōa('4wZ-ĸ7u׽n���+�gq����(9��!��^���^��đS`��U�F��A�����At����tU��� �ɬ�����k�UV	�`*{��1�	|�R�C���h%�����'D ��Wٰ�ݏP� s�d��Xn�fe��@dC�̕~'��䀮 s�fc���>��_��sX:�:�k6�j�)Q�  }��]n���L��bpn�ݱ��8s�8��Vw�3�fc�缎���=@����(�X�9�	B�H�6�{ηu� @��KQT�[˚j��vv[�hH�n%�����c�\���%J�Ǡ l������䀮 �9էw]n�{ծIu�vVf1��bq�����{3�M�5�A��O~�][��       %����%����7��dta�Qr�c�"v9�5����ՙ̶K��a1�laV��t�1Y��%�[�tj���s�I��I��Uk��wNrt�h�vG	IB$q7��1�g��n���F'�����3��nDb�]fc���֋q.�u�[@�B凅��*Vf1�:Fb1�v�\�IWR����)��Zt���䀮 >u����T+c
���yk��P{��D��Ti�N�_Wm�zX�4�gH���w]v��:@�U�F���PxP�_/��� }�}�gq�����:�f:��:9ܒI$�!$*N�^����GJU�t[�{�b�]fg�(A�	�֋q.�z ���4���U����*V�����L:6�꣺�nM󵙘K��@j�@���wX�ﵸ�� �]fcE��	�'��I$Q(�EFRNv�\ƨ��\�1�����{�cH��C�����W�|�.�|������n. s�Vd��19�$܊�̶=�:�aa�B��xP΀���h���y<�0���K�$�I"J!X
�fB"{46yp+3�21���I��r@W9�31�f1;����'z�3��xq�����]�ch�Twq��7�6\R�u����C3X��&�HےI$�H     hF�]����Pkg7c��GV�5����Q��t����J�:�B���quv��#��a�]��p���2m�����>UU�ŦumH�&�H���:�n. s�fc��bs�I��w�u��a�Ƌq.�u�[@�C%����*wXV��C��Vx�f�$pi�C3fc�q��I
�"�Y�`1�C1�;Z���Yd��D�]fcC!�<8�bpfc�W��U�EP������W��뉸�fc������y��Nۋ�H���3��
nH��C9�J��af�$�IHV�U���箛��h����^���aFK�T��c��L;�n��=��$pi�Y~�"����+V�]�&�ۼ�1	޺��>��y��NH���]�cwϗ������Ui�:,��R��q(dq!q�s����}��7u�����n.�|��ﾕ����~�h�9ޱ��cH8���\��u�[= T `5Cug�M,7	P|~�b��n�^x�I$*8��c�٘!� �:Psr���4��!���u�{�n)`f!���f1�fc������v�3����Ƞ���,��`�� ���W��̏�rF�> {�c3��1��m��G�̮ ��߽��g��u30AII$mE��`X%�!L*&j�i���Iibd���\�`�sR��FQ(�фHAY�f�2��)"	"�f�~��i|���#�	&��oz^m�^^km� �m�                                       ������C�w�zj�j�P��<ٮn�P ��Y�N΀   m��w׾!go�=�� �5�9KY�*��qmK�h]�B1���Ss���6P���)�����`:��8�\�V6Q;%س�`�i�]�k[�"��ct�y2Jcki^k��-�<!Դ��u� 7SaR���2���nP���&ڑv���h�f�60%�K(�\�����US2
�k4�6��:�IܛH�U%��^�Q��yT=7iٮ���*��-l��]�s-�b�z��������Wv�u�kfy�'���U�� ;�-Rm�wAc����^fZk���R�\�ϟ��?r��!�h��p	�����Q���C�so��I��B�@      M5�3t�f�`W=Y;l;�n�u==��,��N�9��=�gi��N��8���� 7kh���6�Z�Ĭ�˵t�6ּA|��rn���ߧ��X����kZnуP1nBx�pSq�7�s�u��a�Ƌq.�u�[@�C����J��<k㺆���〮����X�լp��Rg�÷|�����}���a3��tt솛C�7�������]�c�(��4�󉸥n��E�G��3���Cn����qpi�u�u�lNw�7�s���c`�4[�q��u�_��k�域 %e�hH��%v�X��6�h�R�1�3��^�=�N8
�8��B��3���WW��␠��3{�ZЍ�5$
d,�� MPg��k�����<�u۶0�����뉸�fc
��Cw]y�� t�#�F�V���P:J�r7;�31�f?�;��h�;޺��0�s1��K�3�w�iu�'��*U�1��C�4�\ҏ�4���>�}��/$�rv:;�֏��x��G�OWҪ�8�u�X͙��Y��3*�٫/:<�νzՙ���3����bpnۮݱ��W�g\M��fc'ƿC�u���jq��4�Ρ���1���0��@f!���fn�;����������       +r��Nf
"�xg=�b�9�"5ve�M���2��t�;4�
ƫ���ź��),M*�xi]&.��&X)\��	j*�M{4q�!��	2R4[�tg�׽laT+�n�y����%�^�zH�n묪���\@�Wf:�c���Rb���cj�V�6�q�87u��W� ��ň裸IQ��%�Cͮ�ƌrԋ�����ޞ����Cw^޽jq��4��eT� (tm�u~�'{����;�>��������\��޲���wP��z�n�nkU�7P��[њ�j�[`霳h���*�)�〮 s�^c��bg�����\<�u��2������]�v `@?%����5�˻ʕ��x���f:�/�n. h�;�V����P��$�B��# m��V�Ƭinp���'�vw�xp�n����n%�����c�X�ꑢ�J��<@�C3{��18�+�~=���ɔ� 'y���q8�N��f1�PsQ�$�H�P8J���5�ˇB�J�r��=�����la1U��qJ�������3A�n.��C3��1����&�@f!���f1��\Ƌq.�u�[@ϗ��w|�^���y�       {5���M��]&�wf��hK��I�r�mcM�-���<D��/�m�8t�٦�8n5����!�M�����ݻ�v�<� �����VY������Q�ɖ�^�}_G�@�C3{��19!+����3���ބ��u��� ;����N�u۶0�����c���fc f!������oπ��jn�sJ�h��.8�8�]8�f:��>�}��&�@n�!UXh )�y�w�0w�]��\��޶0������)7P}T ;�Ő����OV[�BW,��Bf1��ק޸�rI$�Gqp������Z��O~�{�tO<� ,��NH'f:��@���;�6╝�<k��~������?�J�M	I�ꨁM[.����FU���M�Z!Wu.�j�.� i���L�+R�L��2�(�!
ƨp$*&2&b&1b��CEDX#gdT���k�÷�Y�k��W�J�+`�sB���4�� |�bP�^m�b,2�{�>�-ֳ��N7��P����9��0��`f �����0�'0��I$������Q(��ۜΕu�f�|�1��� ���{8�4[��Y�ǈ�fc�t��'$%pa�C3fc�y�R8S��Q�r�{׹�P��Ěބ�P���;�����<��#�7T�$��{5���UZ+Z˸�3J@cDȣq㍸�}��x���T���h#q��\@�x�f0�s�]�Df6��]n�@���h��9��ܶ0֝�W�OZ-�T��c��3>o_���z������M�Ϙ       ˣh�vh��-Kd)7/ �S��&��43	��[���2��,�M+��`CE������/3����fk&������H���pKh�2Dᐗ�u^:��P󸤐 3�{ηu�j�N�8��x��la�����c���fc�3��S0��r. s�fc��c:�ל�J��F�N�,;-�}��9�pDq�?}�`����|@��wZ-�Z=�Z$H����� ��1�b�O-�T�1c#�7P��W�{���x4�<���n�x�$󸤐 =����1��.dm���+�z����hum����Nx/0���g?!��p��ȥ^� f!����#-��\@�T=�X@&���(Pg�1׻�'{�"R��ZwB��n�*��7�]֋q.�u�y|@�{|���	Z8��::W:WZŉQ��jF�p�+3�1�����}������h Q���w^Q>��$�;κ��0���q�831����9�X���aaVab+J�%��*8܊Uޱ�b��{��t ��Xqt�Ҥ�u�cJ$q7��Z����^�I���C����a�����-ĸ31׽la1_Ƌp����Yu�u��>��a$���[��NWwߕ]�       ��1�S�n�Ps5�&�Y�NGf�V���lX.��݊v��C8e��N�Z����ǆh�6�&sm����O�NH����Y��i�`���ͻ�� �8W8�� 3�w�u��a\9��pfc�ݱ�������{��J��x���fc�x�q7��|����'{���9�w��1� @��J�Z"�����ln���R���K�3{������O��*ھ_<���4���7]{<���!+����3C������� �!~�_}�ÝN8'f:�(P�a�H�����I��Z���I�Eu��e�#��T0��r)Yxǈ�fc^2�M���uÎ�1���0���w�k{���������1^g���>�.u��K�ێ��c�z��4[��Y�ǈ�fc��ՒI$�(������iV�UɭXk���ߣ�'|��^��뇻q��@n�;�Y��-��i�'f:��0�����c�7��l����r��!�BQ��P�BR6�����e_l��n. s�fc��c��I$�D��dE��)n����j�-��y����azt�F���-Ĺ[���@��c���U
n���E�
��5��fc�g���� s�fc-Z뇻q��@ݿ��k�n���7����g�v�%1ՄŊ�����Q�=b�����!��UR>���G,���˓C#=������dV�ջj辒�֤t$��Q`�Y#`��Oే9�Yh9-  4��BU�0�U�����bh�cXqEDFk�5ULEUJ�P��C�� �H�T"��(����(PPE*�,H� 4R�@-P�P�H4�c� �"9 k�"�T�Al|J�RYAHDE@(^j�LH���QAADDҹ
P{�#P�<��	 ��60�nd.-X�f,��R��;��|(UP��D����-�*�����/�"�B�EAj�H���Rlpq�'珲�˧�v�x�x�G�t��y���5�6`7m��n}�x\M���f�=\���0|��=N[�bH����]p���3��(���x���ߙ���������_���h����m��������������G��EAy�Qs%�$J�N�3p��;�|~)�w:'a�?�w��`��<�`������ѯ�s .Zx�'�9��v ���߬@Q�C���7㙑���i�G����oO22=�W��u�a�7#.�Zú��$N���j��)��u�v@�K���"ꯞ���i�����R:�?�4���7z��D���Tv��{~�>�u��^yl�y��fx̤��ֿ����-TM~��s�hn�p�e6S�!�
J�& ��*�Y�INd�B�F R$�)D"DJ�"Q�%FeV�ZU"D"iQ�T�@* �J bT&�R�(RHP�ZP)B�i�)�Q�) W/Le(R�R%*
P�!B-	J��+���0*�(��***��,#"� ��P*�
��D*+*��*T	
U	�BT%QU T$HDXRQ�P�%e%P�T! T!!dT)T"RB�B
HT)T(T$�E�B�BQBXDX	DY%d�E�@��&��%!WvFy1B��eo�%}�eh�Z���?��x��Gz��X����]�'9��QPk�r�" ��Z!hX��h2���s�y��GS���c������u�������]c�tf�"�wsQ3�'yG�}��ۧ�9�7��G�������y�	��u� �.�����l��+P5L�� �Ǩ~������͜2���ٟ玮i��oB~����>�C=��/�]���6���[{=6�����`�:B1��m�N�������������N�� �/?�q*.������Z�[�6������j�l�7`��I�iwKt8�Q`�E��#����g�'�ŀ:�1|�"����xÈ�� ?��>+�(������=�*&Qʬ��h;_��I�UDXkG����F��QU��8!�n�A���RH���t��Q� /��?�)�����k_�C����ina�?ՏŮ��c	�?��PQFxp��'_W�ϸ��Ɖ�<��S� Q�9���� |�:������hr�t-�c�+�����n�����<N ��a��yfE:��W�q��ޣ��1��z�oKA��yYS������uGq�W�7?s׸uLߜ�(����y�C�:���d!C�`0'y���0n@E��/ݠl _+L�����ǩ�����c���{���������<����Laؤ���py��-\�#.X�h��_3����8Mx������=��'co2�<lr��m��L�'��������wA�7���f�U%U������K��T2��vm?�?�����O�ƿ�?�l�>TF�;w0un˟Chf�>I���ޏ�{@G��s�}~��/��v��� 3�x�L(x -��ϱ��듹���T����l�lEG\�������������B7Ϝ�G�;��t�b5�����s��&����jr��.�p� 7�.