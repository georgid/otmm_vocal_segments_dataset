BZh91AY&SY�g�� �_�Py���������`�}`/�@ ������ @���hX��{���e�֔U	J ��J7��T�        �&��6�41M  �����&�L�4��     	OB�)�j�i�����& �(D��<�Dɔi�7�hf���CC5@�I&��i�jyO(h�M��@  2h4��!n�-$$�D�#Ң �@���~P�Q*	
@��/j��"4�OOF�*�"4�ъ���g+�/2�U]3s��1�  /iJRI$  %)J��@  l$��RH�   �+����$�   l����I    �I$�    IUV��H   ��m]X���VG[/�2�7�Ii.ˑu�Ւ�L�m�۸�xS��8Mڝ����w�ݷ^�Zy'�M�xt���/W�� ��E�Jy^�C���<����H��
�b��xˍ�`3��t�����ɉ�k��0�8Ҍ�"�6�-'0�JL"�f+ek��^\��D�ҕ-����s1��E��[Gg��dd�"Mmii�۔Si,�Iz���M6�i ��`1�$�1f�Ȳ���׿�����������g����=�⛓�}R��%�I��E��b�t�H�α�K�՛F�LY4LZaf����IK��L�[��V"2�f�]�1�3^���k+n�r�^��8��Ȳ�5d�WT�T[9�Ff�e]���BN������'���9qky$6�^�γ�IV�!$jg��?�� ��j(��(��(��(��(��(��(��$�HI$I!!!!'��>��/�dEYF��F$�#�"��N:���"
�Ȥ�,�`��hg�ю�IK�Z�
��� �*�
��� �*�
��� �*�
��� �*�
��� �*�
��� �*�
��� ��T!P����HB
��� �.YU��=^�rGL���tE���T����Gi�� �#1�$�f��Vٲ�۰ 6*�����Xʪ���[ޗ������Q"[�/�V�Mt�Y���=������ѭ�+�M��Ml�k6���R4�L:�<�/wqO�Z�@�x��HK��o�~���9w������ �h������r�:���
)��n���4@�rF�Xz+��p#�rnj ��>V#���	���p*p E���G>��7ݙ������m���v�{�y�NW���J�JWFh�7Ms�ҳ��6���_�}�}��w��=V�C ��I�ʙ��D]�F�@��a݀;s F�B��!�E�>�� n��H�%)�癈�tDQ�s��_���| `�7y���&|�Cx �� C�� Y�X����陙��m��m��f[m�0 I��WړL�l�)FYZ�`�DR���Ī���;-�́r��m�,�+�׀�XQղe5=��M��o*� �}� U�o�E.���{��E���m�D�\`j��4��nƚ���DDo����@&N6�����@zV�B�8N�_<� #;�'����<G��JG��1DT�@7�ۈ��%�i���&fffu��m�ۙ�m��V!F�@6"�oS�}�R !� � ��;�tut� 	�Ax�H"|��O-LB�#�?+�� B~�v��d�E�< ��a]� D���x�٬b C��J��y��1<��x��TcYQ�Ç��f�@� @����s:��ι������m��s33m�����������Y1H����r���$�w2K��]vVI�Y����~rF/2H��Y"�A���׀=�{~Zi�G��y��|rϱi��5�#�l,<��s��g����:��àG{9ݟ@���� ��ÿ><`<NK�bl (�j�fz�`B���#Nb|�<�y�9KLc�sV�=~��P#�o��J��q ���v/r5���Ebr�v��g/�@����I.L���km��m�x{/��'����4�ܞKՑ��s�e(��O6|!棣';>d̰d��<σ3,#�#'La<�BHR@�@�B��w����FFtH�@��2E#�8=�{���;�>̣F�����'V1����2IL
��ѧ�K��D�\�+x����q��z�e�R.�LT�J����5N��f���� 5�:e��5�H�U�G%TZh	��
��^+�XIU�n� 7UU[m���9����y�xAyT^��Q�A��Q�$�*2+)��XA��H�U��ʷ���;e�˥�ٮ�i%�K=�t�&��RX��w�Y��� ����w-��WH�Ӱ��k�ގs6 	�䏡!"BA���ݮ�c{��\{A�����g���`L�=܏�((������Ol�
�潶��"�{n�I�`3[q�":�PBS��X&����u�8Ѣ-�͚[^z �UUUU��,+
Ό�6��Yy��K�P��y�@l8�H��	��C�����=���/��w3���a�)���9�]�q��EҨ�y�2���\��Q�0�=���]cisL�Ū�L���M-����^;�uUUUU��A9{��y�EPy9yO_a����X�A)l�|{<��k�6��oN�h���u���'����ڠ��Sr|G����o�]W^T؊��y�7��*EƵ��HX�49� &1���Eɐ����0p�Ĭ���/m��Qq��3v�!�Mi*$��l��$��2D�۞�=�{yD�v8��E�����#B�j��]� UUUUY�"#LI %3C� Rzc,�-�h q��iN��Y Fs�B1"fH����@��	�h��/���N�<�����}��*{ƫ|��8D�	�+�4�P`�����=����� mz�u��Ǹ���|��#�#���'�����FBs�$�@� ��;��=$1���g�;�/���3̵ײ$|U!fubR����RIb�LQE #"�b�Z�
B��"�a"�HH��F*��A�`J!��N;�P�A���@^�(�!�hDZ@o�D:�s�/;� �"��xl���$��e�\����D�����b�e���]=3����EC�PN�D�*	ܨ'��_XC\P}��(~���YP��p"~����%\�}p�*�|�y��i�:r����I$UUUUUUUUUUU9EUUUUUUUUUUUUd�I$�H2�I$�*	��Ϡ��<�7���o�6d���B7}{��9�M��6gǓ��a�D��r�^�ҏ��dB0y6XB;�H�4��un��~��6�{d85Ϋ�D�[ߙ���P�j���𜈈�*�ʿ�u�Gg�F�.]�R�5���{����*:T�k�x��+�ir��i�ݠ�{�9˩@�I?mŎ��sBׁF�6�
�h�#��HE���H2ER)D�IA�-)��Ѝ�2��U�n}�9��)C� r��J-�*��+����0�����1���hx8�F�᰺�m�R�1<˫�즶A�Jӹ���#�Ө�9::��ͫ,���n٬�ۂ�9K4��M�`��n�8����y�e��F\XQz�Bʤ�m6���+��.V}��r�g
�iJ���q��yM��Y<0�s���2"����Q�� ��ꮙ!���I�����R*"m�![��5R��L�X��UBR 1�c��2*�Zꔶ:rh���-G��h!uKrrvw�%uftGqe;z(����o�۸��OƦ���f�Z����e�h�uM%�#�h�����G�xB.�}'��G�/���9�����!P!�����,�,^��h��<���6N���n�=���L��S��K��:n,�Z-g��jRZ����a��ӹ�B!f���K�s9�Zy���S��x0D�΢�K�5]6�r)�	^{�3���k�qʼ�h��x$N�$0}�I��j&�@5��9�w$S�	f{|�