BZh91AY&SYݪ	� �߀Px��g��?���P9'g���a$�6I��O4)�=G��M��P4 ��=@�Ē���  i�� �4�)�&�&�F���B2�&MLL`��D���S&�h�CS�4� ��2TG#���\P�V����G���H(TR������BA��c�N��}�(�H{�P<ۏ�ƛ�p���L~�ƪg	ILm�`��BZ�&Ve��̑��),"��g3�+Bl�ni6�������x
��+�Uf����=��C���� KӃ��D��������A�Y�6)a���)j�p�XLN�&(��&h*�6ݘ�@;�4�������Ut�o ��M���#k�H0�lY �6�hY�a2i@��B�K���0��D��2u
����-��IH�P�[���K��u;�MfV10D C��Y$�˩�NȆJ2`]�ԥ <�m��(��6ɒF����ծ�u��F��Ж�����`��y���z��H�J="�������܏�i�-V�-(�c8(�J�����ND�Я$�!	�dP���N�]F�h��*YI�|��H�yz�_j�������8M�I��j���2Wc%/2@���|�]⴦_��`/��6�2��.n\E�$H:XHo�`�U�lU�?nJ�S吧㻃�!���{E0��d�|�7��(�����8��^�Hx`�W�z����By:/|]8
r�izP�	=o���|睒؊P�@��	��,��3���`%�9��L��)�_���É2~�5���3�k��_��z�ѭ�0�Q�U�t��=mٓƘ��©�Б��!
���5�а�t^$>5)�Hp8v�W�{">��8��A�`����b�a��t��>�"\�w���G(�k+�HC�5X[L30�,v�YT,\���J�S�@���{e���)�KQ���7�B�}�h��"�~5����q� ��{�OA���k7�m�`[�#f���GJKș���3	 $@�Z�_U%�u)��.���o��,U2r��=<<���sC{�H��(C��d̡�N'Hc�ގ����)�θШ\i���x&���>��S��%N&�s�D6�^�\�5�7T��@�mR'�βE�[\�ls���
ڬD���H�
�A7�