BZh91AY&SY4Q�Y �߀py��g������`>z�7<
>S��S�m�Ela]u�ƚ ��)]�޷�����/] : �S	%=��Ҟ��OP� �   ���4� � &��	L(BJ�   h  �T�ԪL`P�	��  �DѢa0���e=FM22mP�4dl�4!iT��I��=@���A�2 �Ƌ�J�:�T*���?��D��?6̅�A@>P  ������$�U �@w��d��0n�A ��E�=�C��οS����w������K�J���bbl�Ĩ�-2��+�QC-˙���%.;���-2�bcM"�X��*)��C2�̳��335��2�-B�L��he��LC6��%`9@ͳ4b0�)�^�/M�&�T+��Ѥ��Ƌ�Q�VbȚ$Će&w�ugIS��Væ�%�����<�v.�ofC�*4���.BW!RW�)E�����&�Jy����ņb]�yq�YLV��2�U�X���&�baK�5{)�f4SH�� !�)K��L#A\�9r�c 8�Q!)#yK�B�"� �"��"�d��C(Ɉ����J\� R�*�-�m1!�b�R�Mmc�br9��F�� 91oeM>L����3,�%5N�l�nﻪ��������K���]�+�qړ�u�Xܑ�[�E)S�4�X�M2\r
�s���a�����=_ �pAꀹr��r�m�d���!p�=~�[A�3���q��H$��;�b���2ژ�Ƌ^R"�H�xؓEc	i�S�L��!����9g�ƶ<hB�]�L��dk��	 6Ұ�n�n�D�.3�Ds�D�Q?��-��󦾾���vffe��f^�fff���ݳ5������UVd�������f]���f��l�ّ3 ڨ�뷷T���I��,��LF=#���76�Ax��l�M��fgm:�Z0�	nŻ���9�C�HH�	�c�p�SۈA�Pɦ"��!�P.V������f���ky�B�4���Z�iA����M+T!b�Y��=�9�wŞt9Ǣwء��.��Cc)T>��!�B/sͱ9I�A��$����@+
㖀���K6�xM흋b:�����)���DB(Î�7d��@�Y�S��=Y����nL4*v�!B����ѹuٴ)d��o�-�I,4yt���J�I�Z+2��	��]U]�Y4ѣ���I�GY�/Mq����Q���^s3�d�֡��:B�
*	���/̈́�q֪\I�N�ޛ��%����sa�����}Ӷ�4�yyH,M�N��:a�q��Ç��ޡ<tp��P��c]���l@<��B��yD5����u��a+(V�=�o[cR��������L8x�ttXp��Sk�аߦŸ����g��*��d��*DPQQ��V���Kv�H��s�*¡�@�ED4W:]�Ѕ���&R����(Q�L�(�T�b����-�qbK�卼h��\�]�t��o��d̑��IQGd�iv���c��"�Z�
�c ��Mq�IӦ"�y!�!!
Q&��Mf�5{8B�v�y<�б�=�׶�sEG��$�K��#�#UǺ'cE)�E:ћ��ٌ;6���D4#��R��s�l�8v<���WLF��2���:9�60a�8RgY�y�Xnw3k��ę�	����I�=C�T�(�
�n�1$dU!DQK0���s0Ѡ��"3��dKtsx��V�.�}��>����0��̐������m�7-�{Զ�!0�n��8oT"҇����0N�{.Kg)��'
�����5ˊ�9̆��2��%����K��<�Fy�k�)uj�_Զ|Y��{0T섥Fd�l�P;v��%�pT�W�6��2�'w˘��Q)I�W3��j=d��Ȯ٦R�t8�(��������,��+�����Q[c��$����mԊb�1�c�@YH �^heCKQL�!^ލD����{3o|�O\{9��}WDvH�au���r�1C
�?U�T�
:�Bl]�
�]9�3H$VK�F)`���Ia�1\£I�TEA�T��mi��
�mEC'�Q>x��|���VFSǍv���6dJ��%#ᛦm�8"O6hѽ:��8!DӐ�<�f�����Hϫ�,ܖ��}=W�a}��D�J�Y>?.�j����jr�>P�S�0�*�����I/��f��Ȳ�²#v*�+��@�;_��T��JNc�P�*��S/u��i���QŅX�f!��0����5%�˄x�uK��U�ι,:QW��X��8�u
0�ĳJ��v&MQЕ�a��l#�*�9D��p�����5b�y�T��)�� ̠�xr�R�B6�9Q\�^{k�=q�� \%�刦"�����Eٌ-~`+Q�
�HdV��;	[��89JE!y��T�C:4JvI���9�C��m�^E�51B�iK���i�V� P��g��, w$Z]�cV�--Hmq��!'�����:Y-\��u��[�=�O\����K�STյ�R�4_[A�����+9̩�J�q
�/Va9;)�rf�*��M=(�h�Ġ�O�ue�)�^�<�X�M�X����fR�:�6�b9V����։p�;=)4D�Տ��K�kJ�/'����,{�PO�x_���v�o�(0�&w�h������D,�Ie����-w$0�*��[�ү �?e6�wpj{�u�w���7WT^�c�X�c�x�to�a`��a���#��GК{���20���7�z�rJ��S���U�V�U�Ωx��řw$�؉�٤�2�C��8C5/I����Ѯ�Y�F,�/��P+S:'5���Ts>S�4��]���m���ˮJ�3��O�-#^�(��U:]=�)�B*�9.����갤V�Jt�zZ��۰d#��H���۝'@�Z��H;Ȩ�
�����S�Uz�p��H�U��ܳ姬D����y쵡�g�m
�Z�r�����ș�{���v!�1����I$�I$R"��t��st�-���<�BI��׫؋�A��9��ɻ�6�$1p�X�ED6,��
Qb��iY�Ո��*�Zj�[�X�bت��Gi)ER,���(�IK(��PF�AE����M�,�`��m�U!XEo�/�X����%@Y$�BE*�_u�J	�#F��,8�m4\�S0a�H�a!��$=���^K���-�F���aa�����4ik���p���w�߆�.H�P;�|=?�658њ&uϞ��\l`�2U�� �|^����IK��<��`��׵+A��� �>���[����b;>�X>pA΀�~�Q, Л�Н������7!�!����RYR����@r��~d7�aҀd_r�~K:�@v�������,C��#qKR�QR�|���v�D�1$�%q,ا.e���N�%��L��`\"/l�W��]b����e�z>BU���9���x}�����I
X#����$AYdT�[��I$@E�H�E�P� BH(eH�w�F�)�4J�(B`��Ay�(���Y�t�Y���	��0�@���	Qj)�"��H��H�#-�epݱ��LiZ�a�c�$MN&p�����9L���{��Pa�xC ���� '�-��k��<��;�ۉ�8`��M�
;��=[C�ȆǢ����H{�MA̽�k��3p��jpP�<tP
��h�Ao9�˔�ꏏ��MC�}  �:@o��;��C�"�LS�3���R&&@���:ho
8�3E,nC���� td	pu�ʹnD�L�I;d�%RQ��7
b�g$1�h����%��bdKA4�0���@(/!�eui���8^���x�{��֊5 =�������^������<w�����۷��'��H��y��C�5&��1�@�>u���� ���@o=���ß:bzs�1 �tiL�bH���>�T����d�$��lGHs��`��_����DEPlQJҡBpQJY�) ,����[�n��6�.�n�HŠi%��%��^&��1�3��PX�xs���e��r�æ��GY&Ȭ��X�r�R mE�zlq0vM��g��@��� i�,pg��n����f66'DC R{��]��B@�F%d