BZh91AY&SY�4���_�pp���g� ����ap@>�   
       �  �  �    ��   � 
D         P��� ���! ���$�$�E( ��R�D )         �a  �  @� 4��K&�g�*����*\3�X��{:��6�Y�Җ�@�L[�9��  />� � �  k  � 	 ���0 	� �   p@ ""�
 +�5 ;7�����|�#]m\�zz��Ӗ��/��x���o>����P�-�-�j��k� y�[ռ'�o����
��}�-��۞Mu�/.�����|Pz��>�zy5���/o]�צ�>�@ $$@  6�
^yU��/)������|�'T�����9��Ox�x�姯O/{j_zT���;����o���y��y�+�z*�=���7����S�J�ܚ�׽�(��j�׾��Z���z综�U� �|     �6��=�U����k��&��o�T�z���W�m���o'^��oW�*_t�;���}���ﾷ{|t�ҹ����E@W=)�����wW��,�{o>���z*����Φ�]�o��}�/_6�����<� "*�  m=��>�r�eg/<m]�}=|���R�z�[��[��+8�{����sy[�E@�ֹ���}��^  =�����^��<��}��[׸�wz�����������Ё�{��rx�������;�y4�         D�Bjm�J�@     ���6U*T 4    Ǫ�JFS� �M4` ��UI"�6��00�O�(������F &# bh�D�FIT�1Lԙ='�2��jx�Q>?��+�����Q��po����D �s��T � @�(* ����  ��������W�B" �T�O��" {�D@���A@ 5�����ߥP^�������^��l�e%�]�l{�������x���9�NMe]�w_e�q�x꼚.�:f�=�x{c�O&v�[�)
�JB�>�����Z֫�I��F��Ȟ�ܪoi]=���,5�D6_����V�4����t�Q4˲Vhӆ���m֦���|n\�]^��Ufѳq�=9u�5�Y�Ѷ�xa�°�=�~��}�yD��	\2{	W�a,��7!r�7s���Z�+7�q�kp�Vk5T�.�=�לKً��}q���5����!��A�4F����"U�h�f�����Q B��u�o�v��F�ˍ���K�⬊ݫ��蛝̟-�g\{+s<��a�$��,� �jPF�����R�X\�����PIt�D����[z6�A$jY���ͦK4@��HbY�����Qt�h$�M&K%*R˹P
�"�j�@<*���[�*R�P�)$*�<ۨQ�9
l3&���Y�������o�������'cG豅kk
�F��Z˼t7)��'ُ��p�Î�Cw��*�Y�40%�$A2����l.�aw�R���P�*�³~�5=2�kǛ8Uˆ���/<Ѣ��w9,�͐��|�HI)�.@�wK�S~xV��W��ɚ�O*sw��-���^V�{%��y��E��T�_*�JM� ��RU5Xi�5�����aYf��|)��Gp�5福P1�HK3[�xzh��Pr9).E�	f-¯��m��i
�r
 \C��nzB�\�Lj�ѡ��$��J������RY�z=�KѳTl�uA�q�-�)-."J�D!R�J.�.b_�ӆM���J����hU�B��HTeF����%A%HT�F� ��RU�Fɞ�7���F�󜛖k�q���zj4�C5�o�|�	���y��W�x����rCU^dM��o2�k&;���ގ����^W��_Eҙ�#c�&R�8��ȔY�M�$e��F��ѩn:rR
����ٙ�y��6Lַxh!�|Z��1Ѳ���*%�f��-D*�Az7�a��fAJ ���Ɇ����y�,�j��I����w��&܂H��fj�n����n��vW���5�T97(���$��HUA�J�fX@�R�B��l�&�V�P�H�e�K�H4� X�%�Y�+s��_��z��u�$�zT/+f�Y��d�CF��4z��Yp�n�Ơ�KXU�B�Q�����R��|8e���Pٸ�%��E����I,������ATPo�"�B��i���-�1�E�7�GbI=�!�6y�k��(�p�l�k�{�m�I����5LK��)��p�O�C���k~>ĸ�HTp�K�38�P]� [ F0)�$�4�H5I/��{����2�&��!��p(j%%JI�xT!����/F�ߵ)<�|<h�'�C�5+^^�W��z�j��kwG��T0.��Eii�sZa����{�c
���z�k~�=ג�B�s[�>k�^&aE�d�l�{=�sTzU�a�x_����7���Vd�*���j�-%����F��*���L�\�X$��/��;�[�yp׻��r�
��[��^^������P�Y\0�����=��2�Sp������6a�V`nVjo{��&�\�U	f��E�r�^^�zza��hh��E�%�a�.7�"Qm��C��n	'�U�6h(j-�n�l|�
.Ri�h͞�"�sZ����
��6CN���51ёӳ�#�J�dnG��L�G�DX��$�)l�T��.p�$��av�j�Idl#PI�Iڪ��s&�rL��F��ƃ T|,�-A�TJ$*	 ��p��u�Qī�ߐ�Nn8�(��(I�.	 Y�\!T$�*���(���B�HV�$�SKP85�
�
#��PѧG��IUI%
�����\i,�
�**4�$�G
�Q*E���Z��YQU	5"A X�ŅP��H$�H�JnbXl��O<��<2Qa�M�kW�I���5�Sf��I+2Q~�$՘B�\�����j�����U��rШb[t4Q*Z��THƪ��E�*�L	P
j	 �	 �j�JB����F�Q��(��w`J�B��$���H��PI)
��0�(%˔�e�.�/
2%�$�H$�IEQ5�����n�7�R�Y�[o&�a.-56�CA�%���"Yfd�[|�xx��NM̂H[�2���,�!�@�	"TE�5y�DZ�+)G|M�L{�t#&悥]�����
-�a/ �I�0�3<(��2XƠ�5s[+R��%E�T�4�0��P,0��f9e�p��eF�kU�*�.7uxz��Z|���;K.w���[��Q�����Cf��!E�p�w��p�1׺�/��^s~o���F>���Jl���<�s�aWZ�r<6^h̔Mюn�����(�5�l�SA=.�n�Ʃ��efku�_V�W��iͱ�a$�������{��{DٹE���
����C{ᛚ�n�m��v��72	!hߞh��k!
�!�����W5�f���K�<��@/E�+݆y��B�Q$�5)��T�����I[Zj2H� D�	AH���.H��&d���@��$$�(n�*\�ۄ2�ۭ����%X�-����SZ��ײ��8�T�2xe��_a��*����=�{c8��ao�~M�|�dA��ND������Z�A�|�a&],.n���uI���ZQ��A2&��
���7W�ܫ��<_fߐ�R�	ljHQp*�]�]�#��ND�٬�TL,�*W�wc�#3�GG���f�T\hޠQfnj-�xK��e70n��E�6ʂB�67TѢd�s[��E��W�@��wI{*�\�r�����B�֡ j*ȁ"���������/1(Ʌ�]�5�Ѭ4FB��U�+=9�
���0��5u�uFh�
����r�$'��jں4�tX���O(�A7 �VzSx5T���&�pn>�q6J�P*	 ��PM����&��	pK�H'�p���ʐ�\��*�5����j	�M�����|�p�4��7Ve���=�y3��\����J�H$��
�H�5Ȥ�n	�A$�I�I�Iʎ���F5*I!21�HD�E���PO�˳}6H�׵�mH^�P��.n����h���ÒI��(��#!$�$Y�5�5B�*TC*�䢂��@����\b+��s[���.�]ɫ橕��2&Z�����$!O�ެ�3*�(�kA�t���57�a�`��#^c�0�Hr�ܩd����{�z�W�.�.�Č���Tn��¡E��!I�Za�Z��.U�J.Se]�l��I0�CE�c*�4�J��V�j�ٞ:��Tij�\��g���L��c�Y9�x�F�yy�'�ߛ7��8yK3[7��m*�ޢ����q����Iw�|��h�B���T H$�aPI�
���	$�%���Q�eB�K�ݠ��	0��P�	$�H�G�f�ȕx�q���TJaQi�( TA��$ �	 ��˗.FK�!
�H$�H$�$F���I(�#P
�)��QQj��PI�HE�U4H�Q(�A$A$A$ �:�7��j��K��
�r�RT0�!q�$j5 J�f��<�XI*�va�%y��D5{�jp���*T-ݙ�@�L۶/�^GL
�M�vՁED���A��E���Vk[5�roe���B��QDZ�%���*-B��S T�ܗ)#���0�̳xԙ�F�Ե��nB�Sm�ɬf�+e9TYU��Q�āP,j-���%B�ZT
*%B�[�/F^{���'�f��r��L�+aAe��Ori􌺣�3^{�e�<9
�2RD�K$*a!UDo�VJB�n%�^5W��	���}͖n�~zQ=�>�.�'��Y���I2��6�
fk!A��Mj�a�w��*�y4h���zk�$�2�&1�Ͽw�񏋭bM,Lb:)��Ncx��N_N�KRqɫn�3�J����?��~����0����B�_��"7?�s�����݇             ��                 �   ��               8 ��   6�     �  8  �>               -�                              �>                                                                䄎-���      m  -��      m�m�m� 6u��V��@kmM �UA�llv���M�   ��m��5�mm�6�;m& �$t�826ȳf���&I�Pl�l m�.��AÎ,q�$ � Hl�� �v��`t�km� ٶ-I�B;^�@	;%�Qm-�   I m���nֶ�m�6� p  �Am �6[P.�f��  $�]���h�cm��h�  ֵ�mt�P�᪕j��݃���   I� :񤩧Fm����uPW>M�.�����Wh╼9�e�Mһ5v��V*�U�
�U�V��w[e���[@     )[l�hH	6۶�#m��-��    Am�m:	V�ٶZ�K�          ���J  d �� 2 R���� )@A����� ��   � 2 R���� )@A����� �p ���  �J �         pd �� 2 R���� )@A����� �p �@
P`8 p (0 8��             �  ��       -� �p �@
P`8 p (0 8��  �[]�t�         
P`8 p (0 8��  �  � 2    �m  l)@H           	�          �       ��              	                              �     |                                                            m�     @ �[d�� ���pK+[t��sJ�ղ���R�U�	���-�   ���e�    �j���    �t��[Ų^� R��$�  mt.�  �  n� �J��    6����s��8  � ��	 [R���m:�
�j� i��5�:uą�/��i�d����n���-��m�^�Ѷ�ɀӶC���+i�/���cC U]U �e��k�V�T��'ijx�n�ad��ؚTKMk �WM���X�I��%�4�!+�M] �5Z}G����h  6���[@8 p (0 8��(0 8��6��  �J  d �� 2 R���� )@A������0 8��  �J-���Z�
�q3���F5F�ujK�I�n϶w�}�6�6Лc��	u]�Ng*	��cjX���(��n��*Ze�L���gR���Gn��z՛XK��莭P��rZ�%�ֱ����-�t��Ǯ�I�m�i��l$�l��,]�����Ցd �v�hh���  ���͍��`*�h�.�aem� �iaU�  [
T`�k���U�kH'M�� h�@l��� �@mٖ�f����`�b�H     m��y�r� k��� ���v�& ĐgXa"�A�Ö�V�U�W��`U���5R�UU+��m�M���M�cm�� ֤��NH�z]� �݀�E98d���p$u�6�v�[n�6� ж�   ����[V�H��a5PN5+֬�VU�wX��e͵�A k m� 6��m:�ݰ[G6�o��ݶ�۶�����9����UTq����S�*{����`���y�b8V��oQ���5Qրn�k6]n�M����&���I�E������6Ӧl�5n�[לp�� $ p�i��V�U*�Q�y�@��չ�ye��T�۝] Ѥ�'GM=rb+���U��EX90ӫi���)��;6�I�ڻuN��ki��YƐ*�^�$+d66���+�����h
�<�l�@�H��-��Uۭ�D�I@7i6 I����ȸU�T���^��V�-Aƫ)WVS��j���K@�h&�e�˶����  6݇Ci��K���i;v�JͰ�M[0㤒B�t�o
­DC� �RX4�]]����{m��Ám6@�<l<�J����j�h
�ʪ�d��U]�U.-�t臵�[z��,�WYTl��5��u�m�%���#P��-C�9o-/��%�j�k` �.�R�� [E��Ӻ�0�\p[Q�B�U�Pq �K�psm�m��U):b��E�mYY�o]�&�'kh�-/Z m�n���L,K��+F��t� 4[h��$丁�<�Z�j��͚A�� �;E��cm�d��8 �� � �C�ݶ�7e�nnP��8)v�j���n�*��scl���v�mV��[N�8�-�I ���U�|�+��7;*��Vʜml���s.��V;��^ڪ�]�5!1�ʻsj]��B�3��5[R���tu�Ժm{mmדv�|>|�Jg8S�5uU! l�5�!<����UeZ�ſo���,��v�  ��:v�4�ce�HbuȥJ����k�"h25@m�U�^�!F6�lj���93iocXiv�av#���j$պ�s�Nv�e�;V	��^���&� �)Ζr�C��gs�YZ3��.vP5����%@j�C�m#���U��@T��*Լ��+۵A¬�۰�m��d�z��rӓ�ۭ�J �O@�ޮkZ�ml�t�2���*V�F�m�r��%�-�   Em�̒�m	6�d���p���i
4+U�UYF�2�΂W0An�T�������Zf�hz�u����)m�6��t�lJڭ@[D�hj�cz���j���b����ΦĀ:H�z�p�5� �[m�v���pp��mn�$��|�OO��o�����E K($ �ۭ�k���&�����6[&$^��m�v	l      ��7m���>�m����6�6�6 � ��p��[D�v�Y��܉�d� t�K�m�Ӯ�M���pr�1�Gq:�Tsq�������};}�ٮ�����v�\��e%yQx�t���v��P z5!�6�vw�aވf�J��=:�Y�2N�uUҲ%*�G��b�km&	-t�d l��`��մI�j�m�kۚ�\�A�//J��R�mf��讕kj��Ņ�"��
�AJ��Umq:�W�����6�p:[�ƒ!z˱��6��֖��j��E�V���9T7/x����+b��5��WB5��98^��'��pB�@mFRz����YEv�%��W`�@��V�l�����J4�����	#b�V������@p�x����W]��KUP��r��޸ŷn�&��ٷ�[��B����b9~U�Dɭ�[� �I���/���W�
�Ua�v��W�*�U��Im��T:JZ]��U�m��Hq�Xu(p��[vԶ��   m���9jjr��m� ٖ�n�7$��Hu�A� m[6���85�� HkgFp�K.�3��-��i#�}~��ְ���h�f�[Nh kn���`5�� j�@u�6� $
X3g]�Y�Tu��&�9��)'��;�3:eZ	�V�[V�K�l��l [5�\ m�l5�SR圥�$t��`�iVU��V���Ԫ���j�pW RQljo�����w�AS�O���� ��9�����Dv�JG��D�䂈�?���-���-��D?��A5� lD؃�E
� ��*�����pS�=@�"@B�g��X������ D���BT�R�JO5������=G�M"���D"�:�Jv��|a��4� �T�"�D��lG��Tv�2{�����S ��<�5F&1�@�PZ�8�x�&�;�W@��#�pP�m@/��i�[8Pf�Nze�6� 5�⏦lU(���b����=	Q�UQ�� D����P�D�ABE�0#b�$#�A�E�`B�� ��dF!"�#�*����aB$I�$bB$."�i"A���Q�b���`�����de(J	 0H` a�b���`őX� E�B! �a$� @�[Мѐl�O�M(r0X1#`H!  ! H$RB@A�� W�\@t�H��_ "��P��E<0ߨiL���k�g��d�0�q�L�M*hU_}PN�Pؒ�� /Ңz�sx"�P<,���Ĉ��PpCJ�J�t��@�]P/�(H�*P����U,6���AS�Q�Av` z�;<?������ �O���K��F����I��"���$�H$�H$�H 
��$�H�I*�
� ��,�H$�H$�H$�H�0�� �ȨH$�H$�H$�� $�� H$��$�H$�H$ � �
��	"$�H$�H$�B	 ��"͐I�J�A$A$A$A$A*�I�I�H#pK�@I�HE�I�I�Y�I �aAD�A$A$A$�hA$A$A$A$A$I�* ȀȈȩ  Ȅ�� �	 �	"`�	 �	 �"H$�@2	 �	 ��H$�H$�H$�� �	 �A!�I�I�I�I�HA$A$A$A$A$I�`�$A$A!�I�I�I�I�HA$A$A$A$A$I�I�I�I�I�A$A$B,A$A$A$A$	�I�I�HH�D �	 �	 �	 �	 �	$�H$�H$�H$�H$�B	 �	 �	 �	 �	 ��H$�H$�H$�H$�H$ �	 �	 �	 �	 �	$�H$�H$�H$�H$�B	 �	 �	 �	 �	 ��H$�H$�H$�DdDi�I�I��i�`n2v���u>  � �P �m�   m��m�` m�H     ��           
 6���:޽�@kf��R���g�6-.�J��@��u�;%�U"��:,��q�3v	��5 :Q��^�m�6[z�nك�2H �0 8��[L� d � 6� "�
P`8 p +� �m� � �p �H�  2 R�����M�� �    �  m�    m���       �  $#mmKz�L<m�ml\k����v�`� �k�U��9�k5��[ ���mm��Z�p�Vu�b�M����l1���� m���];�}�г�E���:bŚ�ܶ���rv��8�q�6ۥ�Xt6��q�+����e��U�H�mPPc�TU���V�T��4-V9��7*�C�ȫs�'ew�\9j���;a��K̾��M[ ��4�Q|�o�|��<B�:x��h��u�%㥊�1���V�t�L���]�EV��F�;
M����:tlFw]��.w::e����u���-�.y�ǔ�Z�Ô�њ��1iD�beU�ccC`@6v��O.�$������#g
q�!�ΛNN��V�o��k��lܝ)����{]�i۴��;�a:�v� ��벳�:�d�T��v� �9�ݖE뛜��p�Ue]K8�;�H�D�J�}k���<�T��a�ں~�*����Y7�n�o�c�ѝ9r���8��b�R�ŷ] ޵�����{s]�����[`�m��q��7k��ܝ�_��}}}��y��;�u���曘��Ԏ��s-e���Z�yb��.#�ꛒɿ?�����O�8�M��U[JP){,�I��@S"�ꪭ��(˼��
�]��;=~:�Q(Bj�j�C W����Ъ�ex���Y�{�e�kv�	`6� m�����]lV�Ե�Ju�  �@6�d ݻe+�n��[[knHZ��e�RJ�u�ٔ�jˇ�\F�] v�M�WHV4�v�N`L�c��9���rXp6Y�=�����z.���V�uv�ͥy%�M�7��՞���m���%��y"�P��q]����mP\0�=�j4�5�%Js0�P(B�t^V��ەvXێ�l=��v{r�� q��;��/��l�UY7vE���8O�l��xz�.�g���,D���>nE�5{u�.W�.V�*�8qJSd�6���swX �W�.V�*Jp*Ur��7ǲ}�`���)' �lӀ%IN ��� I(�(�A�%ԗ_MLV`	RS�)� J�������V��dC�B'�Qb%m�seg$W$#f�V��n�b�;T����v�Tr(�"LrE�*�_ 7wg �lӀn�����x�h6�Md��8� �W�>���>�� i�0�9����H���cs&6��' �c0�)��U�	%x�)ʩ��*����˚� J��O%X �W3�v�ۢ��K!#rO��p<�`I^ �E� J��|T���4�>u�����EZ���X�N�ڡF]�S�u��;q����ʗ�$u�M�`I^ �Z=�	U���U�/ǲ}�bBǓII8�f�u��{�����#w7(s&)>qA7f �78*Jp�>����#�Il�ݚp��c���r)!���pT��I^�Z0�)����Y2|�n. n���٧ �{���� gO�y��<Ğ<q��<�Y'e^��h�^�pٹ� Yu<H���5�lSvϾma)�$��LMc�N���pT���)������T�PPM�we��`	RS�r�� J�Idp��|ib&I�|܋�{^��I^"fo# n����D'鸹&��n�p�ȕ��9%��%IN�}�k{��o��>�1"4��b�)' �F �%8*JpJ�*�Rtvz��Cg�$�J۪���p�+Y������ ��xY\�<�mq���;� �%8*Jp$��Ѳ	���yq���r(�"L�G�=�upwvp���os�Un� g�j4r&�E�SuW8 �W�rK# R���%9�=�x�I�̟6��' ���?u�j�T��I^�Jr�l�
��j�����0)*�9RS�	%xn�3�?���~��$I$���H	)$  �ʹ��έ�ۡ��խ�m�U�%X���}��-(m�����$H�z��[vͱ   �lݷ8�u�6u��q&�%r��G I\�/$��݈�&x����{�� ttE�Uɕ	,�bۃqm�δ�|&E���2D�����@��ݐ[VS����<�Ǒ't$;NY��޷73���gk����l��;���w}���WzD\�=:vȪz�Mx~��|�x��qO�� �h:f�3B��,DɎ8����׵s 7wT���g ��u�xkVjb�)��K������_L������ �IN{>0�.���S�b�)' ��F �%X$�# J���A�%ԗwW0Mـ)IV�,� I)�=�4���Ǜ���Q�D�$��rK# J�Jр)IV�GQ����a��.K��d��n��Gme�h���;.��m�n���[+Buג.� J�Jр)IS���"6A6�8ׅx�0��1�rI�=�4�0a!�A�#�0
"�E5���2 J��S�Se@UA7�ݗ5f
RU�rK# J�Ji�?{��񥈐q?���/ًm�� [l��4�U]���UeL_%21INg 7wg �٧ ջ��n��8�tm��a	"`8�ǎކǇd�6SYP�Bt;]\N���[����&<g�E��RN��N�w_ ���pwvp{=��G�a'� Re%XId`I^ ��c�菾��:K���j9�D�$��[o3���R�<R��H2s����r��^���Q�ۑ5�&bn'3�>�H-�pm� R���Y*�TJ����������9RS�)IV�,� I+�魽�LN8���<�P�S�v�g�zR�{]V�Gi��㛙B�˨���,]��U� �%Y rK# J��}�6�W �����H8�����,� I+�9RS�)IV ��S
h_%21I�� n���{��j���=�����d�TČQ��)'��C �" �V��[u�rK#�ӿ\g3��;8��f�1�I�#��)IVQ�-� K���)�3�\o�����O�a��.Km�@e�i2�vb���fulN7n�\��������!�IWweh�d`\� �IN �$�����mȚɓ��8��8*Jp)*�9%��r�D�������jj��0T��
RU�rK# [8��\mA�7�O�q7 ջ��rK# J�}D�m���r�bK�����j�Ie� �W�/RS�n���'������}�c1��i'$�؛\   6�m%<��C�,�6����ƀ+��[@��`�T�ݰ��   ��Y�$��A�5�/$�ֺۤ �s��ݢ^oN4�8,�tm�#v�U��j�d�
�X��)\Onz�f�_p#ӹ-Nۮ�g�����#�Xv�m�Ty~c�۝�wc��OG��Z�(_FsS��<�}w��;�����䝹ʠa���jZ��+9���^����5v�Է.��٪�:x.�U����}�[��%8T�L`������M�F(�D���{^���}��E���6��������hs)��8�98%IN�,� I+�9RS�zE�y�ڎL�9�H�>�Ŷ�� +n�T��	RS��� ����������0��`�)�;�����ͷ���ߥ~Ip��Z<���sc�Z�]Zïj�)6M���Ν��&�^�����W��M]�ʒ���N�,�}�����WPx��M��=���k���HE[�|֍�s���9�����HFHE���{}��t������3�^�����S�L�RA�9�7u���dwO)��rȕ��Sq2D�a7UUu�.K#�}��rY$��� �W7q�<��fs�hv��W٤4&�m��헙��)��t�;H����3���S�.K#D�}˒���
*��˲��j��~��dh���rY��\}}t<�r&�d�Ɯ�~-��o�x�����?/گq������U����"�2�rY����Qfh��j�(ŊE
����"���2%]Ӗ`%Ţ�QcJm`��B�K�j[E\�ie:�f6Ai�1�)H.�W��^ѡi`4�)�*	���kp	�%F�Vyd�DnQYA��q �$R)�^�-��"6���7X�B�%@*�
$X"ז�(�}Z�UMO(������h��2^�XF��	  �J�dKuz�B&���B�w��&1�pb�T��	)���m=��&SD�HH��{`��AGl
H�H*���{�X�b"\P�Ke0���!���02 L*o҇ �w�P=E<E^E���󨏥�9Z@��R�f;A6 x�z��T�S+J؆àTS���ZRE$M��wC���s�N�].L��jʼ�Ғ"s����qI�/��)"�';��C����W{�Ғ) ����wY5�Lµp̽���X�)"���dRE��@;�~�C�RE=������H��rןt�����!Rcr4ci�J(�pښ%sMԫa��V��=SBire�݊����5��컪��U]�Dp9�Bi��)�w��)"�';\�m?# ��"�W�~�)"�'�O�~���a�+3%�f�qI��ށ�� TRD��߾��RE;]�ץ$RD�y��w�E>��ՅT+.VIYww��I�;�w�w�NW9�Ғ?�茂���_���dS����Ғ)"w��d�S,�%�/*Mk5c��������JH��߻���$S��{zRA ��'�m�O��n
 A��.�����Z���)ʟ~/�wYy30ʫ���JH������)=�)���"���1G�������?��oҿ�:3�Z<�v��OL�E8r�P��e�Ƹg��Y��;�w��]|����e]cyuy���Okﾽ)"�';\�lw�Ns�և�QI�w��>E$R��}e|\���T�^zRE$Nv����'�Z�w��ZRE$N�߾��)"�W{�п�2'���}wY5�Lµp̼�fj�qI�����)"�'~��hw?$j)>��f��I�W~��qI��vwRꪳ&e�f7��RA~ ��w�;�H���}�RE$Nv����) t#�Z�~ޔ�I㝟Q�\��a�+3%�f�qI����)"��"'������`2)��kJH������)"�E�~������l����UUUUUUJ���8���r�<q�[sv�4�5��JlHv���k����|  6[%rpm����.c���cb4� �5�&���]6%���ԆAt���e�^��
���\�l��ۖg��w]8�r�t#�9�j�Ӱ�{��u[�e�j�ϱv�w;gQg�1�dǍ=v��
bl��d������͂G�>�:��y�p�V���@g�Zlnp�$�qy��ŭ��~?��;wѻ��]�d�.�3JH�������;�H�k���I�9�w��y�I�>�4��H�t���2��f7�&����RE;\�o@�䄊\D��߿hw�I���f��I�k���@
�{S�>.�/&fUxff^��I�w�;�H���iI�	-D��߾��RE>���Ғ)"zw��;%��Uц7�W��$Q����)"�';\�sqI�s��) ��y�~�C���w�'�W�ɘ]�K�Y��$RD�k�����@�A��߯JH��߻���$Rw��4��m��{����߭�}��"rK7<��*��A�����r��v�V��.����l3w��{���ኁW�V��&����{�k/+y���)"�W�v���H��;��);�{�QC���QI�W~��qI���}�uUY��/+��Ғ)"s��t;������H ���A�EPj)>���)"�'��w��$S��v���(�b���?�~��\��a�+3%�f�qI����iI�9��;c��} R��W{��I�;�>�C��w��*�*����2e�f���(Dj�߫�}c���}]��ZR��';��C�������4�H��òt��V1��5�Վ�)��;zRE$>�������I�w�恑I��w�;�M�w���~����:����#�\�ɓl�B:��*L�p��U�ݪh��|�?7˟������*���Ғ)"s��t;�Ȥ��iI�9��{j�)"��s��$RD�};_T�K�̫��˫�c�RA=����h�E$N�]���$S��~�)"�;��C�,�r����\���T�u��RE$Nv����)"��s��$|5�<�nB� D`"B"�=[J$b�H� ���z�E��wZ��;�H���iI�;�{]���¦aZ�f^V�5c��� ���}������}��ߴ;�H���}�RA>D?��O�W߿X�)"���~���U�.���/JH������) ���}�RE$�W~��qI�s��)"�'�@�rN���xe�>u���ӧl����l�gmR�$�.��6�랩���ʆ�?,F�����T��2VfK���I����iI�9��{c���v��ޑ~B�"E$N�߾��)"�rt���U�.�*��4��R�s����p���B��~���zRE$O�}���qI����)�R?�#7�?|t�'�YXL��ֳV;�H���ץ$RD�y��w�+�и��}�iIؕ�V}���)�N���Wy�30ʫ�32���|�0*'~��hw�I�>�4��H��s���R@�ݠb�#�]��JH����vNɗu�yY&7�W��$Rw��4��B�X���߾��)"�W{��I�9�w�]�$Ry=�.���VYyw��e��I�W���3�z6nlc�]OK��<��]���=���	7���[.L¯.\��ͩ"�'~�����)��;zRE$Nw���`}`2)>���)"�'���}wFMc�V���yZ�j�w�N�9��'���'~��hw�I�>�4�H��s���H�_�� �S���j�UfK���j�/JH��߻���$Rw��4��*@�"}�����qI�_}����H�=�����+�Y�.�4;�H|F���٥$RD��߾��RE;\�oJH'迈�b�Iq>�����$S�g�?�
*aVd��Wy�RE$Nv����)"��~���Ғ)"w����qI����)"�'��d���ʪ����*�̒�`  �͹z�u�7=�.�b-v�cn���a���p �a&+v�:��6Ā 
��Vx#x�V����7Gn�Ι�e�
P�Y#�m��x2���� �1��n���n�ĝ��t*�i��כv�q�!�&n�aH��\�s�Z�q���<!\�vVL�ӑ��t'$�]���x:[v,\�$����-���w㻺��~I���m�l��+n��+-��+H7���;�Pam�+.�2�Q���(EXR9f�eL����/*Mk5c�E?W�~�)"�';��C���N����	"1 ���b!��D�H���;�w�w�OO�3�mH�D��$|��σ�۶�>�?AXEF""j)>��f��I�W~��qI�s���U`A"`"�J�Ȝ�w�>�.�2�Lo.�4;�H���}�RE$��w�;�����B�?W{��I�;�~�C���r���w&aW�7uu��RAW��TN�]���$S��~�)"�';��C�����Eb$T���٥$RD�߾���ɬs
��L��k5c���v��ޔ�I _�)߻ߦ�Ȥ�O��٥$RO�j�^}��>�୻�D�D��ӧl��Zؚ����ݔ���P;j�ԜSu�� |�z2�+w*�2]e�cW�zRE$N�߾��)"�����$RD�k���"�)�w�^��I㝟Q�]T�XfJ��u���RE'}�s@x�p�`�� �
TRD�կ��甤�}]ϯJH������'��~  �	qOݟ��(��Y��%]�iI�>�_~�c���v��ޔ��H�1B
TN�߾��)"��}�iI�;�Ӳt��VYE�I�f�w� � �� �`��}��JH��߻���$Rw��4����1����w���X�)"��|g���fT��eUᙙzRE$Nw��qI��"}Ͼ�)"�'~�����)��;zRGݷ��������u=���3q��v��!�e�L��ڴ'0q;IȽ-Ľv�/:��������Kɛ�re�f^V3/4>E$R}Ͼ�)"�'��w�;�H�k���U>BTRD��}��qI����0������JH���+���� �� \S�}��Ғ)"s�߿hw�I�{��)�����{�}wFMc�V�je�kXj�qI��߯JH���;��w�lBÂ���, �����3JH���+��X�)"�zr�+W%Vd̻�Ư2����)�{߾�C���O��٥$RD�����qI>"_{��I�>9��U�*V��0����RE'}�sJH���(~�����ؤ�~���zRE$O9��C���v���U���U٣��v��U͕�)1j6�n�;=F{��%�uI��������=�\q����2U�fԑI������)��;/JH���;��w�n%w��iI�9�H��QS���ֳV;�H�k������H������$R~��٥$RA�����pG����>.��2��L��33/JH���~���);�{�RA�D�k�}c���{���Ғ)"{����2�/+	�����$�?��~�)"�'~��~��E<��$}S1�FD�T	 ���"{���$S�8s�]ܙ�^���fiI�=�s���RE�-{�~�"�'���;�H���iI�OA=�N��r�
����Cg��[l��Z�χ<ԗK���H�<8^]�fT/H����u��2kµsS/+Z�X��I���4��H�s��qI����
!��*)"w�߾��RE=���V�J��f]��YY��$RA��t;� |����N�f��I������)<�;�EO�""�"TRA��Ϩ��QR�̕�����);���RE$Nr����"���dRD��t;�H�=�1�aEL��eL�w��$� (A(�D�k�}c���O~�١�%E$O{�wC�����@�U+��٥$RD�ܑ��(����/(��j�qI�w��)"�� ���������I�w�٠dRD�+���)�S
<��K8�Gi����]1�eUQ.�/z��٘ %�F!��ׁz��hՙ��h�!AUd��E����X���(��Qe���VJ�0e^���]���bs��4�h���,)(M��I����ԪX�T"[)�^&�0��m>đ-��w(����U�[vh��t������M�� |�[tm3�/6)�hCh���4�.�9��� 3�3�c37�P��I$�  � m�     ���  m�-�                ~�| 0��m� I���'[�ڊl6��#�NY૦�R(�*����Y�mJ�l�2�a�x.�	魺�����4v1c���=��\��f����s� � d ��-��@A����� �  �J�    �� )Ii� `8 p��m�M��  �  @  �               � p [@��m���JIq��������n�J�UT ��n�3�[�K�`�jlc;<�΃-�d���J���\�P9mR���`�lA�� p (0l�3�.�ѱ�Ӵjب�Ҏ� =����Ƙ�h�vfp�ʇ%-mR◭2c-.Y�T�[@4�D�nm�*��
;U�����Dv^6��TԲ�pF����1cl��v�H�"ԕW#�7�QDҜ;tU�a���|�5�hݞ����`P�er�W�%��nt�(2UI��aS	˷n(��=M�w��te� ��T��U�/<Ê��*Nabg;k�Y,#��[�h�u\����N���K9_[;n�=�E��ЮϘ͓y�3�^���vJ6^�6���v��#/��ب�(�{9���0g������A�mUeZq�"�5�C�E��
b��qS���;Z����w����@ઋ��,��GS�����U�d���϶�y-������Nֺ�=�������f�ᱶ�\9Km���%.�@���n����۔؝���M�l��ǧ��w&�q\^i��uXw�8l�r�7.�f�Uҹ�iڔÂ�y�+a��r���LQV�RJ��2�Vͬ]������4����)�������������!=�h@��⧂�Q� 0��D؞ 4����� A�ӛ�eUUVfd�MfU���  6�m?4��o�}�Z6²�mr]��� �ILmmlj��n�:�ݵ�$  PJmr�`)�����ۤ�m� 2��׵�x�0T��M��sӳ�gRefv7V�b�s�����q��q��x�[gr>//�y��<r��������n�sY�	N�66a;!��m��s#�v5y�\
���w{��w�㵹O�wb���v.m�@e�i2�mT�����gӴ�6]��8���+��F�٭�Uu�P�ɕW�u��RE$N~����$Rs�w4��H<�w��C臑I��߳JH���g~��2�/+�Y�y��RE'=�s@ H��qI����;�Ȥ��f��I����� >�Ý����*��3JH���W{�����w��Ғ� *'>��hw�I�>�4��H���ѓX����z+Uy��$@'��s@Ȥ��{��w�I�y�Ғ '9\�j�qI�ӕ�Z�J�əw��eff��I�����)"��+��٥$RD�k��c���O;�攑���/�?�cѣ����,N62�6V�Q��^[X^�����fZw@��W}w�r���*V��2�Vf�Ȥ�N�f��@�n��Q�9�r���C�A!�����'��b�F�Ȉ&����}_}��G�W��0R�!rI�`2(k2�*�A�4�-%��Lh��� r�/H����
�Ϸ���z� 7گ���5x8�.bK�����6�+@9�x6�� �;��Z��%ƛR!I�6���0�i��� J��Й���|ӼQ�#jG�,y���l� ������y+��|���";��U_Ip��Z<���uqԭu�.��	d��-��%&�5��i�;��}��|�\窦����ku��W�>KV>DD�DG���@^N]Tř|���.���k ;������i�sw�%\�h�����D���18����ށ���槄[�V������c!$ �"�HȌd�d$HF2!1��B2"H"
HB�"*�B����^��>�5	8{읝��T�.ff37�?
�)�X��s��^�������rI��jM��� ��}�RNrt��ªwTeL����I=���jI�`�Ds�[��@��f��U�7C�SJ�i��fs�hv��W	٤4	�Pb�m�6�]����x��ȶ�oGs<�o���m�y+�%�0O���!���A�BS���n-�MT��7vTU��]��՘DG!�A��n�U�� {�_`> � �R{�Ϥ�L����ɕ,˼�g[����U��G"��n�ͧހfe3sl��I��$mH����Dp�M�� ���%�0)r �c��[UT�>�� ��߻8����YϤ��p������l�$��O�������{$�w���$�����Ԙݍ�oQ�ŉ�F�]%v�n��%tZ㍻MZ��n]�h{v��N�f��n�&��� ~��O����n׵W?s�"9 n�}G�扉&��f�໼�=>J����$��� 7[���V���������S2&���7 n�:��� m=�:y����ߢ�F�x���}�Ϗ�l��oz�m|���7_����-�q�ԈRb���' �{�3>���n�m} �v� �~�Ͼ�f�VH�I9 F�x�m�  �m�IҨ���1�Ȕ��W�����(�������sE�6텴-�  �>��tvj�I\��Esu�i��� A���9*NG6���J�,�MI��9)l����.bK��ٳ5CGe�� c���6x�`����Z坴�99�znEz�8ݳ�r�p��v���o]�]r�&
uf�y������'o����=A����HGh[u\��tS���Hⷑ6��k����y�5��ڑ��y��[��U�րy�y}���h0�;��bs'Ͷ�|u�k��f������N����LY���L�t^^v���%�0�ȎA��u:�	V���?{EG�$j5$����}��S���u���u�}�ǚw�(�*b�FH��	'z�m|}���������;n����N��I���39��j���CgւX799��w]C@�`ؤ��gɓ9�Č�ّ�&����k@<Ӽ5��>�4<�`	�|��EL�˲ey�^��󹯺*D�܈���1� �5]v����Ȉ���[��������*���|�y�l�]`G�@�ru��	i�����M�\�rEE�^a��U��@J�:����3�?6�`0�;������QU3wXU�ց��>iށ�������~>����*��NIf㇖�N��vc*�>������nf㞳@�:��n줥���w3�E�yy��i�����N�>�?�f|#^���=�_��0JF�RLR�3RM������O� ˟W~�z$�}I�� �j��ʡG�扉.������7�'�߻z�Nr��or��Y6�JCeR��Ҡ~F�{��Nv����r}TČ�k#"Mǩ?AW�(�w�w�׹$��f�����$�����(�����������}�:�t*�����{��w~�����9����#�V�6l���X�ͳ\���� 1ۂ��(1�^�w�w�;�i�"JLpq�$��������*�������w�<�`���l�"����6}���~�&B#\�u�iޤ������*r��>����+.B��n� _�?ՠi� ���O'X�Z�j��q�bd��@�0�v���w�'+�v�$)��B��׼��~����)�I1E$�����N�u�րy�x{��S��K�:���N�N���u����W8�/j3�n�[��2��w^�I���zƅ�)��N�u���d%�y��=�&PS��ddI�������g�}��N�֞`>�]q�r	Zo�b��a�8���� �]�����W�_@��[��M�Rc���/��|�f[^�X�jU����N��o�mH�F4I;�5{k�]���4�o�Y�TEs���Gy����wo���@�c��W��W�  mok��t��9�k�ӗ��&��ڐ��i2 dp�q m�8��ͱ � ����צV��Ը�uۖt�[l��H��:��\(q�m�M�C<�g^өRcH%�4����9��$����k����0ʽ��� �mA�,��38��Ո낍��cƝͶ�<nܓ��bpr��ݎ�њx�M\����]���:�'ʞ�y�Y����;*��SFr�3j���]v��]v�3.q�2g&6�LQ�(ڑ�?������f�
y:�;�˪�o�{�.���k >Z���Ȃ"AkO0:�t*�U�q�O9'���%�M���M���@���t<�`뛭�J������"RH);��_e{]tu�� |�_A����<��.)��1���7 3=W�}�l�뷽W���36�i��E���bK<�'�V�W6VXհ������<���\�*<K;���Ϣ�r<"Òq���:�j�gګ������ �(��j�2���ywY���N{��o|@q��X(� �*/HjL�wW�	��m} �v�|t�
�#�����U�<�j�:�"��N�@|�y�yf���	1L(ڑ>te�:��ի0J�N���uS`e���.�ʼ�4� I���N� �v��୻�&���<���N��Rׇ�[�~8x�e�o��WF���3�b`"G$���t����5{k����~@+�p��R�,Dd�I ��O'Y s��h�w�$��qre0X�LPM�Ė�����sSG;��l��vz���$��c"CY�jR�Q%�i��� �l����!!HF20����IH�#L��aL)��Rʂ��BPD� w��������H���o����I(G	"�K� ȒDa"�T H�B$��DB�� �&��F,*�C�)�UA�n�y��MS)h��T"�`F\��6��YZS�TT� �v��z���B+\ ����8����[��iUC� `"����U �= =x��J3��"��I��g����+���F�q.\���]�0e_k�#���N�M��#gګ�yR�� �6+PMTȈ�q�$�������z�����9�~��jȳ���1b��l
�����y�e��#��g�OV�M��ڑ��h�w�g�^���7��u�-V�2AkO0�P��U�M\_�USwX:��@<ӼsOt=���fb"w�˪����=�}����� ;��x������&�@�"h��D�6I1E$�뷽W�����v�'��O~dk���R��P
X]�+A 0D50��(��i��R�M���Miv@&��`��k����'}���\��d�I ��@��8��^t��8��ށ�b�m��$�$��X���lɶm�	jf'D�i���]�Ii;:�ǌ��)��1������z�����8�Վ>�S��`.uhq�\���\�\���k <����kO'$�u�ʵ*�?f��	�"���Fԓ��g���z@9O�`롺�4� �sU7P�ƈ�zj���=_�} �v��|o���,��a&&�O�mH��s�n��;�4�@S���[��$B
h�V���<���=�������@U�x���  �ʹ�K9�Z��JM̫�J���V@�I��p	�vu-�fؐ   ����'����7\�å��r��B-��;�>.���h��g�d�=hv;ttGUW��g�x^��V0�,���X�}�V���1�k��6ER�Y�cc�`�̅����9^XHS�w#:�t��cRG]T���;��{���~Ip̽�Z<���dU=\D��χ����Z�#��%�
7?~��K�\m@9>�\��q���9ԍ���gګ�r9��[���K+(H�d�RNw��w��f�m|�����l��>��/��nz*b�FH��
N�[��W�_@?]��o����re0X�5�q�3�9�7Z@i� ���)�� ���E�&����������]����_ 3=W�}�6��RE𡏘f�p[l
/)٤4��ZDy���������]i�D�Ɏ@M�$�'RN��{��u�s�n��4� �sU7w��*S/7�I����im�)R
S��@B� �F�H�HH0bH�0!$A,�R���4
;���w{�O=�sRM�՘�"�Sn�*�&���wU7u�5�����;�}���Ot<�`���VI7�d���5��ܞ
�Ŀ���H���϶W;!�^J����� ����$�p�뷽5{k��־�~�g �_i1�1��i&�9�s,Qsek%�8���v��G�zK�tl�v��"bFFH��
N�^������a��}v��o��()��0ɉ�����U��TӾ����@l�Uto��~��q@�����l����r�mc(̯y]��s����$<9�h&Ԉ�aRN�v��j�םUy*�s>i�@����M�\�q$T�����U��9���4�jݽ����f��_i[�SR4���%6S���k�I=��V��b�T.ԜK�<�6�LX������d��w�kI�}�)�����M����9�]��yZ��	��@�O'\k���ٟ�f�.0#��LQI}V���ju���[� �j����*bFFH"I��3��^��$�o���$�w��I��0!甔+!5o�F��	�&&�.*�j�z�[s�D@�w�&���Npæ�{O>u���Z�(͔q@dPa�v݆�˶9I�+���m��q���� �w�&���Ns��nt
�M��6��06���^��6�Z�n��;��P��Y c������ O���Ӽ4�����uTq57˲��z�D����i�@պ� J�O@ߒ�U6_.��"����Ӽ M'�7i΁�e��>ߕ��6�NH���n�  ��i�޷�"��]�l�55t۬� 
����86�8��6�Զ�   �6��0r�6�:�t���N�k��@
S���6��4��p14Z��� �2�E����t��jJ崽V:�$[����y$����NmV�/(ۻimc�Z�pl6S[;q���õ�|�`�����Z��Ѭ����ެh���^i�-D���B�Ó	jn�\q�EN��3s�.���5,I�0#��LQI<����@��\k����s�
T�K&7$�Iށkڸ�>*���@�����{�|\�AL(œ�ȸ_�U�
V�� ��Y����Kv���9���H�q���*�_ ��ozU�z"%גw�8QI��MܗW�sSwX�Otn��ϒw�9i� �
۱��x�28<yQam�s��N=�gq1�\u�,]�+;�U���^ѥ$qd��D�z�j�?n��*�d��_۷�V\�6�LML�H6��Nל�s|@Ұc�C$�k��I;�s��%Z��"#�'ɺuWA�]��"��u�� �]jB�G���9�����/�U$Q�I�� ����'8�mށ�`9���1�I!$�@��\�[g@��|��ހfg�$VݎLjc��q�<�ӶQ��54h%�s�:�ҧ]CҘ��fw�bd�gL(œ#r.W���Uv�wm�@��\���ߢD�ɷy��9i� �ot�9��nw*B�ǴjDG2,q5#�v��I��;Z��Pr� H�I�j�]��:�����¢6�qd��Bs�*�=O�W�)Z������(�Ѷb�����Wm����v��
�����ZejIcMcQf㇖�N��vc(�v�\���H���U�2W]����aو�\�I8�9:^��Z�`
}��H9i���,��]��wSw]��� �S���jW�*�ָ���Ҧ���$���$�� r�w�9�� m7� .\ ��bn���������cM� �S��;�w�ܞ�T��(���z�y�C�r�K*�l.L��o S�U�6���?����*��t�֝�dX8Ad ���#�V�6l���]hl�15�ː�!6㉗�(��a��M���R>wm�@��_ �����
���?Sw
�ڒ�b��RM^`
}���29���u:�v��,��a&!̟F%#�y�zt��&�@rӬ�n�U�vb$1r$�|�����]�{�*�_ ����.�T\`"F�RL����K0�C��`u�xU�z�SŲl�R��}�� ���n�h�b9�(H
�"B
�,)�0��JQ����u�%
Y!)  L�$"@�UHƐ�2P��7�2�����*ev�K�wI�|    � m�p    p [@  �                   0`l ���v[`���Z�Bnd�޺��ڥYIiT^�-F�^����d-V_h�á�ntV�J��3�I[��e���ڌٗ���#h���  R����-�E� 2 R��� ��� �p �8    �p (1-0   d�pm�Y��� �  �  h     6�         [@�m���fn�E�-�Ƶ��i5u]mv� � 6�&��m,��rVQ/kj[&)�ͻU�����;u�C��F�u�@�m� 8�� b��K�2��e��kλ�r3�v�5!��toK�4p�m��FN&����s�65�s&ۗL�mFq��z�T�������ض�UfZH��m[���@��L�������z�Օ���ݕ�����X�g��I����i
z]�fIcO;�d�ue:�s�ћ]Lp�ez6��w5�kv�m�v��x�	�B2E�����[ ���J�G8|�le\v��zWY��<k�n!�W�n�qX�s�z�M�<fNr�����7N�]��r�n��f�Xsv:�Fu�lE�8�盃Yd�rp�.��52u�/g\������j����7Xf ��\�I���ԑ�]��9t�v^�8��L����wW-ΝU\�-f��9x����n�ѷc=� ub:7g��Z�V��Ql��Ů���)y).��ِz;�Wq�Ԣ����Wv3��r�g���7[X��)�P�=q�I7=ku�]*6�]K�;d-���D�,q7*�Ai��z��U�Rܪ��2����s+30���@�v� ؼqP�y���!� �n�Ne�j	�b@������e\���M�bM�   (v1�;i��ӆ8��3k$���(���@�`�9ā�l-���  #e�W��孰XY�wKcZ�� �*����f�d�l�6�4On�%f1V{WB��]==v3�X��fy��x9���WIpqۣ`{���Mړ,�L�F���QԎ�mg<;����I�W�֙Y7:�5;����!_�t�>u���N��*��h'X�Eb��;(�$g]d���tg[�".�e�2Đr^�V�|��΁kڸ�oz��>�`�JɊG|��΁Uj���%�����&O�7�&,����2ｼ�Nz�	f o����n[:��jDG �ģ������KM��kw��J�*�=�n��R8����z��p�ϳ1/�o�]'=y%�
]2�U.��"f���n8yn�Nʽh��9v�\�:��2ݕՅW����:�\jפ�_[o������:Npɽ��� D{�Ӫ�¦d�35���f����ՠа��F@:�"���ŉVʻ�G�D(�ǽ�w@97x�Mށ�h��5�dM��/���}l�{m���\�É�M,�$�]��|���&�@�I� �7���>�`�Q�&(��' ��l��j����}l�v��k&,y ���<�ԭ���V[��J�����S�(r����W%#���>��7��s��z���_[{����U�l�ˎ�M�*�ss5W=y%�� ���Rn��ڸ���DmH�ɓ��z�{�ԓ��w��^ؼBB,`/��n:~������Pnd�/�R]]�D�I��5�s��Y��g ��]n0��H.}$��''@�{W@^If o����u+�"#��h:��%�#��zt�T�]�Y���O���m��fN�7;,��f���b�&�������@7��V�z���~�hiSHDC��d�N�}l���$9����9�u(��(�)�'�tL\M�M��>I^�Z���&ZM� -n�{�ĹdŕW6&_{��<�{Z�w��w�$��jO3�E)�0�z��F�[t/�{����=:_;%]�e̋I��ݷ� �[8^�΁�������ٴ)��Ia<q8�,.K�l�Re�ۚ����s�������v��L"#jGL�4��� ]����[g@�{W ����~3ٹcM��!>�K���
|��ʵOG��G"e��`����?~��q�f"As�$�99:��=n��9�kw�̐s���5Cu'B%$ț��]�{����U�l��j�=��M!a�#�+���� �w�s�� i7���{A: �����]�eT���%^��l   6ٷ:�I:ٹ�K�����mn� 6���M� g
ݫ���ͱ   �lݶYV�Զ�[��9�ݧJ��(	uA��m��5��J�����I��sr�cj3��oVp���x�N�.��7%�ݛ�:{\68m��q�f����<��3�l�n�ѷ1��3t8n9x�M�in{0��ۆ���{�����7��U���U`��j�l��y�AӢm��I���4�P����}c��!*� ��w�yV��u,�`�����B\�b�n�K��/���<�T����o:w��q�U�l���jDG2/��j�p�{���7�\�u�t�u�y������������W�)�J�O�WA�9��`0�C�����B}#��U�l�^��ݷ� ��g �ȭ�����px�1@U=DK=e�0ظ�m��F�*�Z��ny�Y���ݕ�]V]�^���� �ot���z�:�-h���"I�� ������	�,Eʓ��椝�{�����������M!"9"��'��נ9\��<�`&�@\8����LQ�I8^�΁��]�{�޶p�����nF��9ɀz}����7�5'}O�+�#���m��;�*=��0��%���2�Bn�B��F���e�l�[8���s[
Q���������� >�W��R���T����ڎD�DBD��@?z���n��N�����66��(�QO�Drp
��΁����|fG|(d�DF���-�JBЉB��o��0�0`�1�9໭^w��O��L�n���:����ݕ�]���������=M� }䯠��ڝ����0HD��� ���� ��g ���΁��_ƕ&7cF1��!lpڗ2�6V�;WZ���6��g/be�N�y�Ԙb@ȚB&!�G$Rw��l�
~���=>�O�&D�j`�78��b��I�*��y{k������l�H�o�Y�hQRs��
Ru�o�=�sw�9�'zC�tjDF�,qE#������l��=�sr ��4�7U�;z�o���HڎD�DBD��@?z�p����?V���/�m�@�Ҷ������6y�	M�T��R�֍[��D�[3ۃk�x�9��l�y2F�Q(��F���~���=>�]}�X�Ȉ����kw�7|��]�Dݕ�]��e��<�F ���~���U��g@��xc	��$Wu��՘����eϵ;�6u:�=�M!"9"�� ��g ���^����8�E?j~�6/�nbI�&.&ꉻ����j��9��� ��� ~���w|-�$�RH	|�Ĕ�I   m��u���ѧ_G\Jr��͞ڪ�ȡ@m�����5�7�gR۶m�   -�Jmr�`�WUŒ��m�:�#���/�ٴ�a[����o��ʕ�������\ݻ]h�6ݹ�˰��=��3'��bRn9����J��l�e�[���ۄmf��n�Z��;��M����j�뎗�=���{���`���<��fs�hv��6Q����ְ2��au�.�÷����|�6no���Т:���^������[8_��tfe�h&Ԉ��X��>��o�sw�9��<�`��ڎD�DBD��@?z�p>��@��� ~��@�
��M�����R]]�}�ށ��� ���{����-�0}>R�I'''@�����՘������j��$X�h�v���!4㇖�Wek��p�[U��m����s���5;v������tMu�`��������y7zO'X��M!
8�Rw��l����1O���"8��͝ŗ�}>�]������'��,B�Y1dxԏ�U��Ο�ؖ�N��O0��W@�x#aL]M]�rl�e�<�`�=�=<�`}�΁��ڑ�����_{oz���Ϲ��:y:��������Z<�v��5�E8҆�jn�c�xk�<,nyT�[iI��5�+��m�9���������'�L(P�b�G�8�_�l�^����g�D}!���{�)��V���˻��{��t�u�>��ODG��&*��������]�V���ȾA�łE�X�5�eʠ�^B�1&.� B�4aaֱ ��d���e��]��qH�D�=�g�D&�P�PA�eQYmGN�'�c=.�V��e� � H� �yB@$A$A$f�$@�Ф��IG���Gzܕ)�=K�� ��yj��P�*��*ąS7�I��3�@����ix7ŀ�Q������%"�Ԉo��q|@�;u�n�!���΍/m+g �̊9$R>}����� s�n��;�{��ZB"�qIށ�z��*��g@=�����{�Em��jc��q�>gi��Gh�u����K�w%��m:�KҘ��fw`O���17�H�_�l���p�m�@��k���7)��!1Dd�{x�ګ���L�uC�ӭ�@S���s&��6U7ss7aw77u��y�zy��������������)��);�޶p
�z��{]8Nz������Wk;�7$�:w.��*������� s�n��;�r{��l���V���4�5�b����z� �r��\��ہ-iu��+���n�)����+>�������� }��2{��W�l��V�09�G&8��?L���@��u�9�7W���~���&�M$�!�Q���[���_�l���p�m�@���Qb�&&�������ܞ��n�������Ӑ��:�9:�m��3�{����n�����Ȉ9ȅ�o����ۄ���&�  Jʫ���f݊PV,�2m6�M NPmm�m��� m�h[N   ��tr�ً��a�.�s����vWc���J��h�m:�=��9=��p�9)l��u�t�"ėe��B�*��h�Y�:{n�G�5���$��� z�l\6�絴��������[x����d5V����q�������w����;Y��t6y�����M�+.(�76n��v�s��6�,��A�=�m�(�+k���������� s�n�G�z}2n���=���F�r,S"1H�����u�9�6^���� ����
;i�$'��>W�[:���}�Y�}>J���{e:�
��ݕ�]���2�)���'����Ϲ��;i[8�`�#�L�H����@��k��[g@����?f{�5�c����Cg��;dU;����#�g��qW�Lh�ֹꍪcrsl�@:3q0�����������zO'X4���.�󛘙XC
�.�/RNW��s
�4e��G&D����w��^`O������������LqS����8����~^��
�z��=��h&Ԋ% ]�M���=�=<�`}�ހw'x�zЍ��JdFI������Y�7zܝ��=��R��&je��V�@C�)����u � ���X�Pݴ���=H���v�?6����_�^�$�^ �����`�	��V���˻��{��{U��G8H=�� ��u���"&MLuGh

����������S���U��o""��ʛ�vt��8��
T�K"��I�""}Z�t>�� ��Ut��f�/���)�LM�R>������_ �}����Z��֝�d@�A�3<�d;R�깲��V�0-����E܌�2�IHбx�(,�'2c����^�X�'����O6�@�Sa5S"�H(�|�m�@��k�����<���Sv�mG"S"2E���n�<۽����ot�P��M��!2���m� �����������������RO~��j�+H�����3//@;���ot�־����?#�[u(��6y�ӶES��Lzw��#ሶ��z��[;��ٜ�8:!ȣ�RN��������+��m� �m��4���D9�9$����� Sͻ��� ���D$n_��	��[g@=�p�3��&|�,��u�3�L)�b�f츫�o3/@;���otO7X]+nt}q�	�"�Hi��=v����� ��w�t�����F|g��%UQL"����H�0�۱�{~~��9���
�V��  m��M�oo^x�k�9x�,��IR0h����� G݈[[-8m����[l\q�P+=:�Kӻk���� $ky��f]z��V�u�p"S�	�=����#��.��톸8��.g�e3�O�8�7���vc��m���EpK���m���nqf��c9���]:�*^��%�Y�9ߏww��>Qݧ�a��.Km�@B�#T�]�sX^{\u�m��-ɧ���f�ⶔ���(�ށ��_ ��t/m|��{�<�srƛQ"Bd��6y7zO'X�otO7Y����G�E�N������k��gS���Գ ��k���΁�l���rd�w]������=:�t�jW�z}�����M$�6�I��}�����)�������R�d�M_rv�D0qYԵW6VU�Ә�E�N�v�M�$��|��>��n�^J~m�Sɻ��� �M���� ���Ü�e�^^T��{�O}�sZ���"90YKR�guW@�V�X���s�&��8a5Sw73V]�M��CM���W�7�m} ������#j91)1w77y�}>J��-��|Χ]���yf��6�D��<#��o��Xz}���R���U���:�wE�Rmhl�Ӌm�T�q�Yn�<��8]v1��Z��nT�t�~7���7ץ�}?;^J�]�f��*y �Sw�j�?�8�`�E�"���m��<���
u7x�ګ�#���$sS39S	$�N�-�Ӏj��:LO�}�I E��҈�\��oRM���z��O���17�H��[g@��� ������É�6L]L��Uɷ������u�kM���� S�l������I?�N9�Ʀ����vi]���g�p�-�G��({z��ajEp�E#�����?/Z��[g@����=M���H%�(��@�|�ůu�xΧ]�R��
4ډ ��>����{]84���n���	��3ꪼ̼��[0i��=<�`K�"#�P����k�k}��<�gn欅�x\�]ŕvt-K0�V�X�m��l� �SRcv4cx�M�bp�s,Qsek#�t����lHcQ�e��.�y��v��Ф�F��I"������j��t�ت��oz�O���17�H��mށ�V��otO'X�&�1u3WaW&�f^��V��ot/m|W���{뎅��bNbr��otO'X�m�l��[0f�ڎD��Rw�~^���[o ��h�Z�c���F6�!D�O�	�2Q(��:B�@��!@D!v�h��
��Ցd$
,�U��� "9�bȁ�]��D���e�bF���#
HЄ(46e5J�B�	�e%0"��Q�$1#	�T�$IS{4�4%k4�Db�AJ;����� Dc	$(#@@!W��HĪ��(e��#!V�����0B��#�mQ	l�Q"E3#�g<�%mܪ�d}H6��⒩3�q�	�[���PJeA��B�S\=���]������  /Z  �    h   [@                  8  l �lN���]�\�Z��]9K���W=m�mP D��%��j7]5mA�cb��m-v�4��N5�Zn��'f��T�n̶D�'m. �p �@
P`�C (0 86� $� �p �@
P    a@A���%h� d ������    � H   ��    m�        � 	 ��f���I+� �b,��I��gYm��f�( �
���4k�\�"��v�'CAd�i� �{�aز*�$u�@�A�m�J  d �4uU�j�)է2��5��I��"�v8,�u�����J�b1�S��r�R��Mm-�<��Ȓ�UF�Tzq��+�.�sS^�kiQ��f��� W�l��q��Հ�l����ܙ��^��3ۛ��l,��T �,qf5��$g��v���� ��jh �]�b9��#�Ҽ�/g��j�=<�{m���5�U����7�n�w�1�g=��u]x����f'S]nvP3͈櫕 ����ݥ槐ֱ��]�1����M�n�qn(��s�۞����#��=��\�FNCo&,���͎G`�V�J��K�g\���c���p�Z���@��k��K�ʊ�-׭.Ո88��l�,�-U�3m����gw9��s�D�F�a��)�jx�pN�k���u�l��h�;&��=��%����)��*��z�7'�!ۂ�bxy����m�e"#��;���t�ů0���T��S��ke]YA4n5B���%���:�����s����,nF�UU�u���o�{��|8���>��OS�`b(z��<@�ҫ��{��3*��[�Im   fW��/bۮ��檆a����+5d���0�a&Cu�ԛ]�m�   -�f�Vl�H
A���- �b��6�L%��G���9d��s/d�Bn�K��r[qڞ�*݇�j���g\
���8v���8�����ˎ�S����u��g�6��uРַ9yQ�#�%'�1��GKl<06�;k�^���v������+Ip�I����HJm��D��u�p^���\�N���Y��q.��<�6�����q�?-���~��pT���N���n���>��>������=�ـsM���� N�u�rel��9�G'��p�oz��~ϳ䶽�}��S�m�A�i%��0�������� �&�@�+f}�J�o����}TX�0ɉ�jG�6�����c4���=<�`����#�ߴq�<��fs�hv��6!� ��7Z�m�<���4�lsF�CM��:A�������9;�`	��@��u�#��>�� �>�N��`)�
�������&�&���;������� !�"D7'J� ^��ֆO�c0bL.�n��nɘ�����=<�`	�n�r�`
��\�Z�j�	�xG ����=�ـ&���>��#��O�`Dy(�����>��>������=�ـ&�ށ�{k�^����X�����4��p��J�v�Þ�l�C��e���.i��a�>�#��r}� ۶��~^��׶����)�6��4��ڸ.��n�@��ut��ܭ�{oz�~�U!L2bo���m}�y���jg��Rڊ�;�~�{�r�ϯRM�t���Q�U��/޳W�>Q��u�@M7���U�5V�X�R5"Q�	I ۶��~^��׶��K����=��p��ȇ�%����g�r���mZ�.dŵ�U����c���U\����H%�"�N���_ ����?y�\n�ށ�.n:�p_HL�Auu�5V�X�����&��������A:}7f}UWY���{�T�Z�`�gө�@N�u�{P���\\�]���z""SM��zu:���ɾ�"� �C\���P�a���IdmL$�);�?/m|�2""��|�����R��*M��ur\��fs�NӶR��i�6p�ւ]�-ט�u���-v���ϯDq��\/%?6߯�Mց�� M7����z/��S7w%\^v�XޭS�"i��<��>��z�A�"Q�	Is�5jY�}>�]L�I��=�����ڎD�H�����1y��|:M���T���� 9�CAN�j���xG ����?y�\n�ށ�{r�s�j�I)$�RA��  m��-�zg�ˊ�ٖm���e� 8RS�[@@� �#�v�Զ�   *�D.�yn�R�[-�NIڬu�� 29m�k�[���֕����fW�^�\m孱�Xy"�c<��lM�6�B�G��Ԏ��J��Ct,�="k'f�MA���k!b)׎^�s�AtS!�6t�zI�Iz��aXw��Q"�j�Y]ffX]�r��-d��z��Q���s�ۧ�]7*���l�s�FF���͹�����{]�\ Գ �}��s� �&� �ԝ�dM���.�m�@�������xޭS�Ȏrd{*&I.�n�����:S�Xt��Ӿ���� \��@�/���)�LM�R>����>�j���If�r}Z�t�8\spL]L�ܕq{���{�9�6�@��u�z����Zv5�`� ���'�V�6l���O7Vn�4�Aw��ae��&8ܸ�������.�.�z���Z�� ��u�=^���=��m7hF�r% "eL���W���O���!K*���u1D#l=T������B�� �)�$�0WA�-39�N���'��{Z}m���H�?���m8/��X��>��u�}��="93���3 ��u�;��Y.�)|ۏ��}���p�K0�ګ��]�� �ԝ�*
�������pͽ�=<�`�7Z��\���ݎdjc��������iT�Kr�l[\H�0W3 m��U������g�"6�HI;�?/m|��~�ڸ��ށ|_��E�S��Ƥ|��U�&Om'=ko0�ګ�2f�S�"H�2w���{^��7����X(=�!�z hu���������'\[5w3uUe܅��C#�������yV�XޭS�7�M�H���N���_ ����?y�\��ހ~4�j�bO8��qr�l� �&Wm�Փ����X�wig@���$sɏm8/��<#��]{k�z�O@^Ic�#��S����n���ưɦ��5���I��ּ>@S�Nȋ����>���n�����'h
��.j��ww=ZK0�ګ��DL������?�nm$"2`܄�tO'XT��ܭ���&>�"�����o?t��>�,Bs,M�R> �&�@�Rs�>m���� �1���ѳٸ�3<�d;R�깲��V�R��Wg5c93�V�Y\�&8���k�75����{�9�6�@��u�5I��=qܠ�R%p��p�oz��]{k����i�B6��)�黢��@�� ��h�9�7{���[N�!<jE�.���Ԝ��{�y�s�j�n���>��>������Rs�>m��I� ��_@y�f�nM�F�I� 7�ro   ������Si�.�a��Pڪ(��(���@�`�9��v���i�  V�۵̒�� �5Wh����kl�p�g	Λ�	�~Q�? ��d;]`��+,S7w(�h�[����]�5����Ƿh�m=-��\{��������<W�Κ9wlv�:y��;'mw��Pu�
cM����׽��96U��ľ����N�OW,�wEA�;�k���=)!�1��9�Zoh��L��>�E�?��?���{W ����7�j����B#jawv]��t��Rn�Ԝ��{����'�?VQR��vU�V��v���h�9�L�m��I��/��\]ܕvgo���V�s����!�W�p�������ܠ�R%p��pͽ�<�9���h�9�<����twi�f㋒�`P���&Wn�P/=�hh�pj�u7Etft��;jŮz����Γ��Mր����ot.z�m8/��G�p\��_f��B(��(eH�Ȁ5
����B!���Q	AU^�B!髹��v�$����ڸw�k#��!ϛjs���.�� |��Γ��N���n���S#nO��p�oz���u�o���-�M�ĄF��I	'p�j��㜈�Zۿ�[I�@[�f~����۾����;r�8��C`vM�e���!΋��z������<��1�|�"K���������n��j���R��{W �������L�!��Nrt�Np���<�9��N��DD�ߢ�0��������B�΀ַ�ʵOK|77�ߜ!5��SeY�����H�z	yXF]����������IE�6yv�J0�-Ov�xJBY�="�!40$��m+���
@ڧ���=��� �mKڀp,�ڨ�z(�JP�-C��*k�<��A\�-��N����s}B�j9�>R2]��I� �w�.�� k�� �⢶��B<xԋ�U�l��W ����~�j����cSR4��=8��N�:����yV���z�\�E�I���8��t�Hs���|���`&�@�� sͻ�=��I�CR�>�E�.���ڸ^�΁�{W ��M�ĄF�b�BIށ��s�9����9�M��\P�DǓx���U�l��p�n�!߾������W�H�uL�(��"FlT/�}��������1%���Wy۾���s�4��Γ��6�DL�����*=�Ϙfs���@��;4�p�ب��[�����6y��.({\�[#@Kf6+t�y�yV��
|��|�F��������M�w��j���"ds����sЙ[�}�d!��uSVO&캊����u�x�mn��ʵO ��-d`�|�9�mr>rt��p�{�y�s�9����l��*�n����8ݷ��{W ����7���I4xE��6	rI �E���.��J[%$�` UU*��[n9[��x�Yn�5��8���M� g
ݫ���ͱ   �l�E�A�	[���Sv.[,�R��8�;:��'�J�(m�-ջA5Ɉ�y��U.v��[�,��<�s�rv"v����/>
�]���Ԃ�����]]�q˺���m�[�6.�ȼ�e�,Re��)���ow�����w{��]���/ԛ�� -�6����6��CE�\�:v�Dg���]c�;5^݁��B#ja$��7�Z���z�}����@�/�[X��&&�U\�y�z�l�M��I���7��H�'y''@�l� ����_=��U�l�����(��]��&�@}I� �w�>�� ��B�j9�>R2Iށ|��W�����\?%�-�@�h�����6�6y��`wI)]@���7��vM�u��'[�M(��ZyqGͷ���L�ժz�%��9Ȉ�A�'=���e�[�^n�f������B�r"9

'uf`ժz�$�#��C�	�����&��ws�M��S�}��}2�<w�.�� }*	�.�n�����#��;Nz�m���K���wm��/���V�2cɉ�M���N��ـ5���I��=���{O>u���sӶR�!� �rv�@U�m�3�	�$�捬�6z�]�3u9�����o����,�>U�_9��:�����s�jD(���� ��{�>U�z�-W�o�������&)��Jd�)��RG���\�[gN���� /���ԓ|�{��!�gjv���ݗQQSw=�r]kn����M��I����.�t�j�>��ˬ��+f �ot:Np<ӽ�������&�p��J�v�%�]{l#Ѯ�,��=N���9���j�W����ot:Np<ӿސi�� ~�	�ėU7��wy�|�T��r9ș�N�����,��ˊTɑ���&��z�}����@�^��;�s~�`�d�rw���|���5���I�|�>�" � �BT�H�P���[:�=�	�"j`�!�/���<�9��N��ـ{�
����skhl�g��W0,Z"�����3Zz㶄��Ĭ�����R;jŮu��?�t��y�z�l���@!�0���5"�z�}����@�^��/�:��t�9����N���G@[�>t��:Ӽ�R��`�A5'��p����{W@S��Ds��u�^�"eA1%�M�wv]�`*�=�֝��l�}oz��s0�ǜk��D�JI/��m    m�^�un/>�� f��Hxj��1iCm5�6"G�gR۶m�   -��m�-��,�4�˺��m:�#���/ V�.u	��Ӑ�c�����<Ղ���$C��N����d1�����zL�7lu������q=��.��O'nsvNEg��"���pռk��нr��ntK|9�����I��6�1��:��y�;`U��u��ݺq��*�S�+����ȗi�ݍ^��q�v�^?[o�_����-]f �o0��=~o�L!�F);��N�}����@�^��*��t��ڑ
5;� i7��'8�mހ�[0�QȔɈ�N���\�[o �m�����5����y5qu5s�9���	+f �ot:np�������}��*s̳q��Y'e^��c(�n�t=��ۃ1J�>�=���#��v>���Ȣ�*�/@I[0�{�y�q?�����u�x�s3]�"���"j�*�΀�R�Q��~��"9�;'{M�@�u�}we9�$n���b#ja$���Λ����+��""e%l�&� �;�E�P	��NE�*��tݔ�v�ށ��W ��f�T�bjBAI�w��$��I��<���n�7���G�N��P[hl�d�	[s&M�h:7g:+B�l�2u�^]Rc�˵�4bj��p�oz��\��׹��=@�2�Q���������M�w�ҔߦMU|�@��� ^I�C��8���<x���v�����p���B!�4XT���H�G<�O}���������'M\v(����X��:��� �v��:I��mI><0x�!�Ȥ� �۷��=�m��`�h�}���]\]M�+Z<���"��4H��v�J�v�r�m�!ۄ�q�c�8<"6�HI;�?Wj�5�N��� ^I����nbI���&�� �I:�V�y'���\7�R�u�n�o۫0q3�M�@��N�(�9 �!�7���@�]��v�s��5�	���� ,�	�lH��6�|{��f椝>��>.�/2�"�7t]�`*Jz��V΁�n���kVH�I���b�1�0 !ӆ)2�m����n%oN'Is�Ƒ�t�:u�ck�F7"F<I��;^�}we8�ݸ��7=�7%�N%\v,����X��:�d^I��M�@�[��{jI����ndRC�o��ށ��� �I:�V�(8l�&$��������ϝ�=�I:�7v��7��ށ|;�A|����NL\����V�y'��78�r�C�"�9�9Yuʚ��H�pm�Ā�
Sx������#�	��J���L$IO?��� B@2�0���)�R o`R�LF�0,]��b%%�<�e(�^h�!I���r2*zɐ��0�M꣠1���HD�B����"�y��ֈ!�/~B�SuU�-x    ��  �    H l  m�H                   0 ���ΖYd��"F�n��[��N�N4�/l�R�۵u<�F������1��f�`bSB��	:��?>n������d`��3U`d�I. �������� )Cm�G  d ��8  8    �JYy� A�����M�� �   �  �     �         h  -�q�,h�^�U���my�$6���K\ �l�ZS��
���PK�x��f�ں,�W�Z����5G]�t�M�$ �c�� )@A���u�27i꤮l�[��dl
ii���ogn�t�qO����n�ZD	��ֱ���	Kv�eIf��e����������6� �'N&�k�L�gR���a�2�5�2zS���w��riN�7QYҩ���kc�=Q�[$Q�T�W�δ�c3��<��g��z����s��^zȼ�=�jw<�s�v3�lh�Mmjn��ζu�$����<���yny�vvn�0Yz�D�nP��W���؞Q3t�c�Ʌ�����4�Y��[i{N5粧���bA�G��uJ�v!�O�n8��=;��'<��Dᮺc�B��gJ$XƷl��!:M�bx�1h��\�$A#:�b�.˩�m���[���ゑ�fj��w]�Y�vCѻ:ې���b7&���Ѝ��\�\rӸ�tC��#��ZM��n�||W��ǒ�Tn:|C^��$��)ܖ�87.�ӝNӻms���]b3a�%ڪ�,�b2Sgp���v��v
B�.�ok�Y/e�A�<UU�S`#*����:V��Ӏ�~m���)j�"��E�Q=6��l�űu�	�k2���2L�n�&�   ��t�����՜:%X��0�p�j�P4����86�8h�ݰ��   ��G3��gH-�5Ƶ�[իI4� �GU���q�%���`��CaqB�R��=��#�Us���΋����N�km�S�-�ݍvU�5��-���skZ;�(�����w.�v�o�9�\m,��>.p8������y��>�z D55�Woԝ:��fy��v�m�f���Qdvꌐݹʜ1��KêLx�>��	Z��������/$�@�� �I:�9�Рӑ� rn���ڸkݯ�n� ��t.6��)��%w�ʒ����U`�h�9��<�����Ӊr$LI��;^�}%l��{�y�s�.��PN�%\v,����X��:���ș��|�'X���S����n��e�YQQn��*�k�K>��X���k���zq�1��9�(� ��.Ȫ���������b�m��l�8�i��<HDs褃���<�������P��{��_^��m�~�Y����iO�9�y6ApUD����$� ��o۫0��������ՅT��ə++<�j���Uk����y�}���G#�?;I��)G�&Ԉ��X9��oz嶾��k�ݔ�>�A�Ya<q9����^f�/>�J����AJ땈�5Z��Na�a1��L�)$�@����;i'Z%l����z9��������.	��]$�@�V�{����v���U<��N�SE�Z�K�FK+Z�^����ԓ~���s�4�B-Ah`����]����~�����;�@��'ǆ$1�]��or{�zRu��>�o�h��0�<Z<HDmL�LNN��v��RN�%l�7�=�H�3ES��!QVC�-U͕�κ��$M�����]��]�|�		�dP_(a0oq��{���m=�X��G���t;/��㙉r�)��z�Ngؑ�v�w�y[��=��뛔9���8��� ���@��� �RN�%l�~�QȔ��#���ݯ���^O���$��Ϧ�Ë� �B ���!C�X�y�}�����ͧ$0R>��v���}��x���� �wUt�U;���)6�6y��"���R��Xn�y(��`]m���:����c��c���:����� �V΁����>��S�쏜��i:�7o�I����nHp�ٷ�����餝hJـ%�$�PU���M]��I����hJـov����T�92I ��_@�V�{��ғ���_9��$��蛛�̭�[0�OtJN���k��)��H��X�% 6�   �kzY{KgN{&nͬ��mZ�T�(!��R��G݈[[-8m�����u��F�Vn��˺�d�� eYǕ5�#��WK�"��J��Y�6nm�ejv�x/<槇��K�����Ɠ(:N����ղ)�.sv��hMF�m���v���K�|)��ٓ.�Q�8)��ЯZw��n���|z��b���g<���
^3�HG<��,س�u��Z�#�Zu�Ի	�LMI梙�Ń������@��Ut��U��C�[:�4*���f�������ғ�}I:�<�� �{o{Ͼ��3|TVӉ��) �W'Z��`ܞ���`j	r8��"J�Ȳ�s/+@�V�{����U�|�9?z�u�{S���AEQvEU�VY�or{;!�I��";���x[?��M*LnƌcoI�,Njh��.eX��k�l\ݼiz�8�g&]a�U��͞�G&''z�_ �����?n�g �oz�w����#��}�n���Oc�Q����tI<�?-���{7�$!�F)_8���G@�y,��DL�uޤ�`Q���ڑ<��!�;�[ށ�m��~��k�ݔ�?]���J}>Rdr� �u*�9ǻ��_�[:{�f}�m�5�	D���iE���6IJ���e��n[���:;s̳c���/&�`�]�%�5u�y��:%l�s{�zSu�5r8��"J�Ȳ��3'@䭘�otJn�>��{�y9��x`�C��}�{�?-�����!ɨ�u�3�rN���jI�H���bK��.��j�0?O�7]�m��9+f ���qNsd�6ApU�]��@�zҜƥ�`u��>�J��B�ӑ|G��A���y	6Ҏ"��N;=Ղ�n�az�&-�S�����^���蛹�����+f ���қ���}Ȍ���n~��5������ʹ���������`}m΁�[0�~-aq��L�I�Iށ�m��~������N��[ހf�VӉ�����8��r"��q��&~J���ܞ���X DX�B�?AI%w���I?|O�T�\��T�4d�����9+f ��� �n�>��@�;�ߟַ�~���&�p��J��ҍ�mW+� q���3�U��7���n�4]�Ue�ـ-�� >ԯ�|�iN�9�N��t�1�����.��j�4ɲ�>��@�V�w7��T�L��N��Z��e8�������/�ٿU1#�lR'���rV�w7����Hy��:�r�15"'q`�8����fd�7x��s�{v��?r=̍�q�Ֆ�hIo�%�  J����vvz�v���u�cn���f@�I��pd7]�I��fؐ  ۶n�:�zآ^�o\4�݋���A�嬲Ge���E�VX�lp2����vƋv!F�<&���uKͶ�]w��x��'-z`�6۞z���;�����Jv9ƭ.53�r7�.h!��Y�Y:�{\�$�5���w�������g�{ߏ���#�N���Z<��pJۧ�E�j���$Y���.	��cs�Q�.�)9s����-�?��?_KW@�� �z��7�Em8�� �	��?>��@䭘�otɻ�27ȗ3WT��eV��[0�{�n���s��Ϟ�s�G�9��AtE՗wf ��� �l�ϭ��<���_aKG��GQɉ�ހ~ݳ�y��:��`���2?$d������>u����v��V�4�9�T)�{n��h0�u�tfi�ç*_T���$�/�?��`� 7�^ �t/�MĢ�2]�̫�j�7U�9����w�� �H���nT����ܒw������w���ďg����&�C��,� i~����}m΁䭘�k���I�2LrN������t۲�}�{���
�q!�A&���֔��K���y�n���?����O���y�Y����;*���˭�m.�����l�5�ak��f��\\�����Td]L�fd�Jـ.�t�Y�?_KE�?{jK�x`�Fdp�C ^��@<��ϭ��<�� }-�J(����@?n��?_KWg����s�tkF��h�<4&��搅X�$���j(r���;]M�^� ����FW�!$� �$�IIL*$�鏀�$6%F�hw6±�!$f]�
�[��b��@�D����$�Q!��Le��Qa*�I��!�5e�@��v�"x�z�<� x���Lh@cD�v��������*P%ޞ$
	xXxVg�cJ����IdQ���f��<�Q�iZ)%JƼ![ނ$H4�h���缧� �c),��&��� $��4:Z���_�a�8�f�<��E�j�P�H����YAĉphެD�01@�>�Q}U�;��xp����R�D��@⧏�������vj�m��)A
l�M�\we��@ϕ� �u� ��{�i� �t/��L�5vUsu�h�� ��{�i���S�n�i�k"��@"px���J۪��ˮm����K;b;J�2u�^]S��mbjD<O �!�${ח� �v�ߕ��"#$7�h���UM���\ww{�i��v��֌�i���e�P��$I8YN�޽:9�y�����j�QAQ��qغ�k�0��:�-X�Ϥ4�yO P&˲ȒC�� ������:��Se@U�Wswg@��ڳ <Ӽ7��{����D}��&�i��:���N�OQ��m�<�a��e�i�f�6�瘗�ns<'��1wW}���x��0�Z0y����T�L��N��S���t=O0����.)��"j욉���4�ـy�{�i��v�����&�C�'� r��o;�4� �;f��F�N��T�]���]�]���w�o�� �u�0z��@f,ϳ�nؒII %�RH  ��i�m��v��﾿V^���]�n��%0m���p	87nKn�ے   [Cm�sm����j�]�On�$u�� �H巉�f6x�̀�84[XGd���J�՝�ܷ�8���63ͳ�:��7	�I���ݹ���p��M{��۫]g�oAgmX�F�a����̲-��1ɗs
�hv]٘�b ��o3,*����.V�@C�Rev��М�ۈy���ciB��ڣ�b�6�Hd�D$�����zt���?���9Hi�@j�\PTi%\d]I5�h�� ��{�i���V���ؑ��WPx�fG"�΁��� �j��g�;g@�m��{�բ�x�"8��ǉ�ހ~�g ��)�w�р{�=���6O�d]�ww�o�� �u� �4�@<Ӽ~���U�����홞y��k�see�L�F5�z��f���5êLx�>���<5Mm��l�7�=�4� �+f��f�1�bq�"!�;���o�a���"����_���{ϳ�ԓ�=�MI=?�k���D�FI;��l��vz~�9;�t��"&}�<�q�T��IE�Ėwx�jp�Z0sOt�;��8�IWs5���.V���� �N�T��xU~��f_mhl�ӧl��Z�χ:��\�k����0��1��q\e�JY헴�*4_���4� �MN��F��:*�,Dq8���@?]��w]��=��N�yj��2=)�l�M�\wfff��v��jI��&��kd��&�0���0��/�B⛂bJ�.�����r�`�{�i���G�O�[s�z��b#D�� r�۷����*Jz��Ӡ=�"K����a��.Km�@e�i2�tʻn�"N�o8#;Xe�qSv1;\��Wm]U��n�~�^�����4��8��j$�FO�'' �{��{ޚp]�ޞH������q�Έs9�$��.���`�{�m������9U0x��H�� �ݽ��l����I��� �
��tꒆ��ȈV΀��]LėE��]r��0ͻ�5�S�wu� �݀�r9~��ʈ`��j�l��uצ��֎y��.2��i$���wNT����	uw�k�� ��F�'����ǲ�T�b#����)�=woz`���v���?n{49���8���ٓ�Ǻ����DG�>�M� ��tf�Suw3wwwy��%V�X�Ss�L�u� �ܞ�8� ꦮf�./깚��5�S�yu� ��W�|��feϷ]���rH�o���   m��&�I�r@t�92��QEr�[[hd��,��l-�m8  F��٫e�e�X�ꎩw]cZ�� ��g#r����j�χ�g;v�;vF
�Y��tmhgk���L�%S�J�����w�q��×��|�C��2f�㱇��;�fz뱶p��s� �ۮ�W\f�N
u�L0�30��Ԑ(��	 �S^o�ⴗ	I����HJl
�6:��Y�4Lq�,����n�];^�4��\\���f�75��^���0�{�)�� r�V�����<���$RC�m�{�O7X�ʰ.�`�҉u3]uu�U��
y���U�yu� M���JSd�l�૲���9ȗKUt-�tkV`�&T�u����7�Li���}=vS�m�{�5z��*�k�����RE���A��ևl
Sc;4��b�;n���u&x+�\P���&)>q��n��^��
�����N�]aq��9��$���;^����1�dY@�d�IE�D$Y$T ��I�	 
���wz�w��֤���{�����k&O�I��*�k����	��@s�� �	ĸ���&�2&��'2��9�i�盬��������<���!��m�� ���k�`V�����@��6e��&�+�c���+\ʱ�@����۸���d$ɗ@���{r8��N�U���7X�ʰ]\� M����2�/�brH� �}��n���6ݽ�z��/��~�`����^���';�wu��Q��
���
�u���hs&'qaws�r�O�η]J��A�#��Jٵp���a����Q�D���z���mt��-�� I���Uv�b3�ֆ�=!�;��*��.�0��FGh�Ƴ��9Wq˷J0']v�X�ʰԔ�	4�@r����q�Όs9���s��]v�~�1#v���U��U���g�g��WPx��B7 ���w�U��U���{��w�墭,D� �7'z��33�v�k�9z��o�vz��" �. )!"An����4�^���w\��$�e�k%5�L*�˛��
W����g��G92�O07����j֝��<28ǎc��S�"���2oV9k� 9Ғq1ё��M���c�1�S��]v��v��U��W���7s١�Dh��ɬ��n�Y�&Kt���[]�7ջ=��Cj9s&9'z[k�_k�纸��ހf�Рۑ5�'�$��8��z��-���n�Y�����)ݷ]��qAXr��U5����-����DG&j�i��9Nlw�_@���^#�j��  ��A ��w��"����*���qB �7
isxU� �B�U�DBAE� �#TD�  E� Q��� � H*�"B

"�7 *n%�P�aT A.
1@YT�U5t �D$T�Z��n ��]$UDU�(�@� �2*�ddE�* ������P����EPdTQd$@�@DoQS���/����������_�����������.��������?��������������ʯ������ ��D�z�<����O���� �D�� �2�'���G��H�?��8�?��?�?��D@ >?䘟�����_��g?���R@�7���������O�_���A�G��������AAu�I)R	AH)0 $H�Q $TH!! R#R) ED�H�@�@� R�D�Q"1Q ��D�D������Q �0 ��D�# R$H�"Q#1Q"0 $H�TH�TH @��$H�@��Q"�Q �Q �H� RAH�TH!
�D��H� R"�"	R*� R�TH0 �ED�� �H�Q (@�!(,H
�Q ��Q"�H �TH*H�H1Q  AD�$H� �D�Q $TH	�Q �H� ��Q"� �AH�$H ,TH��H�D��D��ED�# R �AH�AD��Q$H�@��Q"$HH,@�(D"�B D",B*D"�A"  A �D ��� ��B"�*A!��H�@H�@ ,*� ��B("� �� ,B 0H� B"E��B
A"	"�@ � ��@�0� @��@�BDE1BB@�dV"	 �B*D���B�P#" ��A�@��@�BD	!`DD�@�EQ@*"��)�� ���"(�*$��D �@F �QF �A���)G����HM���w��� � 
?����������� �W�!��������Q 
�ۆ_��<��������?���'�  �l=�?��}J � �ȉ����  ?��c~�*  ���V�?���f&Ɖ��QG��?�r�χ��뱿G�  �Co����������� ���@Y�����`�����)D@ <���?���D ���#�5�=2����c
%��������]Cx<y���: 3���0��P�?��4���RE�=�~p���O���!���E �?�?����Q  ��(5�g�	��-�������'I��S����PVI��N�����=�` ������\�� 	
�J�@%B�@ ((��� �

 +� ��      ��$��E���(�� *�E	%U )PH *�T  
`   1 �  Q,c
�ѝ�A���;�{��X0 �%��O�i˧kq]� ������� i�a͹�j� ת��<WZ�=��a��Ў�{���Uz]^*�۠9����b���E�R <@T
  b�(�P�p #��
b  P/ ܥ)K�
]�t�Q�QL���� +( G`(�  �b)� bh 0 �c4��� �� ���q�:
Jb4s�(@H(    (�0�:
&���޷����n'J�^˞Ͼ�_�����﷐��P.�7a� ��=>���{�����99��A�����������[�r>�����}��� |<@	@!@ K0�	�=���6�ƺrj}�������W;>o��{����q ��:S'���ݼ��7g>�wq +���ﳧ˫����������g=�{ܾ�O���q�z��� @   
R�H�O���s��9{�� о���s�z�/N�wxƗÀ�d�]�� /����7ʊ��cں8��rh�r��� {x�]�^N{z{��_�}��    ��j)�*�� hhz�f�R� d O��&Ҕ����R�z)*1 M1O�BSmT�*   �LҔU A�/���/��(���w�y`�*j;n�$�B�Wл���*�*�������ࢊ��"�*�PUN�O�		��2�@��B���D�������?�����k����,	 ZSy�[ҹd��վV������"��BK΄ Pt:I$ �X�ѯ)��q�h�Pӡ`�`�0#],0%B2!]����y5V�ߖ�6��I�^�~K�WՓ�L�Qa yU~흴�IT�A	X�%b�#ʸ�mf�2�!�y"o-��-ל5��3�1�:U�E�ă�M9��2ћ0����)�X�8`�����#]8�`F�01���DtL4F(�x�$M�e��癞\1 P�]f�pd��?�ٰ�<�JK�h������r5#���1ƚƆ�"�F4*jE�F��d�t4"CFN�������R�O)[��J�z�|�-
b��(�͈�-,�Ty�D
l^�Ψ��H�xT�5��,H`A��%1hh�p������R6K� ��a]0͜���4Ȅ$�K���٣���^MRSXv�
�JHIJ�[�����Zuaԣał�HT4�!t��h��
��jcM4!�����h�n%�ސ�<.�3�s|<SF���6��W4�)du��*�M!���H��.��X4!���"� Cg�%Ma�0����s~���1��a�pZ�PJ�E�<��ܥ�����SQ����0Extm�SZ$�.�;������!$���t������8���ĕюE"!a	@�G��m+	vc�kV�ȄBֻ��veR��b���R)ZŒ��h4�p"��b@��ftpr����]��R��J�yF�.�T�*���ط�v��j�,}i���BQZH��SF?�]Xa��@UJW�{)�EZ�oڈW�Չz�j���sgƍ6w?>��4�Y]C6,it��nf��7|��G�K���
\|��;�"4B��CDR)��h6�`WI���4��l1�� WA���)� ���6bƎ�p��u��s�U#���G�2�$�Q�Q�׃�మ�Ǆi�6xp�3rf��d]A����B�YÔ�l XI@��x�"��ќ,ش��l�RA�B%�Hf���0����x�	����
'௩
�;x	k���i���h�	 S�a6L�b;S��͋��V����)bKГC���i�5�Iv�so�S��j0 ��p?@��6����)�� l��� U�R)I��)DH��6sF����rnl�ќ�����SCŅ]�c�a��?g��V_0�y�4Ƒ*i�g����� �FCi���2?�'�!M16���4�����į!
r��Y���Yʒ&�E�y�4]�*��ol�n|��.7׵>\��%4�o�?aMh���DX�`¤+�!5R�;Io�		ʕb�����������I �a
h����� ��!�4�hA � ���o���7��V�m sV�p�Ӳ2:6�p�4-'�Y���5'U�^F�J�����h��X�'��L$��8$$��q�GA�ќ̈́� 0b@�8�!i�H��k��6k\64@���Y���
uF���!J�"B:1��F�Iv���$ �4c���$3{�ф6�16p���`]9�~=�������~ �I��8~y����)t~�N
`x���k�Cs �\4�\�!��8x~�5�8�p Ĉth0��d�4�L��E�~9�$��(����SX�V%�t�(��/^Q��j��"b���J^��d��-;v���"B���Y���,˨k!��\���xqk�aG\<��$x��`D�5$�<9��X�3���������6��~S�����$]a���4ћ8~�E�������pY,�*z$����R0'�p'���_�k��q��E��h��Rsjf�$Jk1p2%`�X�d	B��M�P!�HB�dA�$RB	d�B���CMbWi�@��҄���B4�h�1�k��&@�����a�1"]1��5�l`WEcLi��0��
d�RJ�R�jFb���gBJj�It"%W�h�du�d��ٶ�?l���"IP��
��`WF~3�����ؿ��WK�r'�ėf�D�"�"���[$H�|xp?i.��.�P�o��č�g��o�l���r�Z��^/���J��)��
I�R�aM����p�pa!SYt�����oF���kg2�"j����	��¾>8k"a
h�x�F~!*��e�r+r�bB�Ji{:��,�?C��82o�1?�:CaI+nr������o�����}�|79)H������F��B�5�
xI��tf�p���a�%���a���HQ�|O!dt9��SK��B�7�9�ᣎ,��kZt�E�@� �`B4�\����F���w勲�{*Q܉ׅ�̇�w~o~<]l#H�,�#B�V%IA���X�����R!'pW�ݩj\��Q�?y'+�������B���$FU|Vڴ	�����vt��~hѷ�ǁ��(J���0)���	�6H6A�r�
��P���WZ3#@�ҙ$a
�B�aL6��D���#M��ܒx��hH�E�q%t�ˣ��=,��x�NoG�������^�	��HX2G�����H�bؕԦ�tz��$"�@����j��mH R
�?�dnt�	  @X�X4q���4����B�4a��WA�
Ƶ�4��D4~?«Z	Md��y��0)ui,���
����8n��eѡÏ��)�#!])$
�4��	�%�ݥ�I�B'�)p6�6 T4�A�����yMo���^^��=x8$`h`ة��f~��5a�3.�h�Bf�]hƚS�{@��
�B��`F�F�R_64c�q?�����:��ݬG���H�=4��E_���nc@�3PĹ���Φ9��ƛ���͡5�8o^r�l��
���Ƒ��
a���i0,B� kA�]p�"e����~�egme"qdZ!���r}�MRBԪT�iѩ 0Hu0��c࿰��n�C�x],H��Ձ��2E��<��3��ԑ�¡ �xĀ����s��a��1�~�k��,,�c �5L��[5!!���V p+B6<��z� 9R����RZ�5h���7\X�A�$M�X�W�j��G�i�ºH]�peMXc�SXH���J�p����P��h�?<3��)�P�~?E�@ZOKyy8�)�| ;75�$#$`��4l��
I	�kxBK#�B���W�G_��1ך)41"m�D ����L�q�4��@���HSF48�����	Ml�y��ь��9\<��3\5���7R'�"E�$Hid�*������6"I[�=�2=R�	t1(��)��"�?{�fffffff`                 �                                �                         6�p�z�v�٣�Λnm�m����� 6���|ۚ۰    �ᵬ�.�Ŵ�m��lI�Y@  ��8�` $ [��mm� �N��ʗ��5=T�:�\7b���P 6ؓ����*�tL�[�"�`m�G�o��ݖ��^j�8�^j��V�Z,�Ҏ�
���r�K��4�M���+a���"�6�7Pn�f�m�Q[r��J��� h   m��V�� �8�Kj�6�aā%(� ��%��6̲�!,��kv䴜:.`                                 m                                 �                     ��|                 mU�                        h          |                                 l��                 ���>                         $  p                                      @ ��                     ��    :��Y��G^��	bj���XhV�Z�^;\e� ��K[i l��v�l   � ���UJ�h� �"���d*���]���LWV�M�l<�  �m��J��nl	8��m���6��u���t�
�VS�B��ni vd�����`�ŝzA���  ��A�8�'RF M�ճ_K�u�B@x�yP��U�MK=��@������&�lgkj�Wi�I'\m��;gk5 j۷I� 崛\�u�9P���K�UPT�	�W2����UTm�	%�l�  P�beUj���
� �F��[P ;H@LT�ְ$����mp$� R�km��i��G�d9�IP�,5T���\��5*�P��幪U�`b�V�W��yh
���U{`[@�M�zp�V�U��I�Z���^vK��CnĶ�.�&�mm �d�z�Lְl��m�� [J�KT �Z�U������%��I��jۀ "CF�ݛe�N kn��@I�Xն�pP+�a�ZT�В��_ N�Iŵ��,�6�j�-�m6��At���UҭXv�*�U�9]<y���ޢ�����������W�Fw8s�dZi5�ּ�^�l���h��)�AUUV�a&m�)uV Ԙ���bmdknĀ �@�^�-�kpt�6ٶ�m�mv�4P�d�8ڥ[�Ԥ�U*�U�J����e6@� ��8�lsi66��j�`s���5]R�E0UR��*�-��  ��HeT
Wf�Z�e$꫞A4�sr˰뀨�Q��u��|��ר[�Ö^Z�A�h�m�������ڪ�@ۥ���a�PY[�i!܇0�r�[[u���vr��Um[����^J�9��9ڪ���0Z��3!�ضAS3U��<����U@I��.K�tS~�_:@�kg��4�-u����f��[ٶ�<�m�3P
�L%ڕ@j�r�Q����}�}��m�8H�ζ�m�m�Z�V�@	-�����ll ���^����1��RU�P%{nc��  �����ZӒ:��#iP�UU�vV��m�(E�V�6�m�*e��`��rP��jP����۰�R��bC�����hU��r�!��Q��m2�[&���v�� m�]�En���b�n�� �u� -�	a�:��$fٷk8��E��  Ά����"eٴ� ;m�R�`���ݶ m�� �(���*��W�4������7U@NH6�|| �m����Rt�Mkt�Y�b�EH��-m�  ���� 6�D�I���6�n�I����C�Y]ڥZ�	�����m����Ik���Z�UW��^S�؞b��We�*���K�+�;�kvscj�RYWc����皭���y�\��8wg@��g�g��<[��ɗ@.�֫Hf�։������K*˼[a�},����H5� �۴��_^��r�`������UWGT� μ�UV���2ݳVͶ�$2�V�{e� �Q�]I�z��k@�� �J��������v�����&��vZ\\6��� ͳl ;�۰[ӥ��Jp-�m�6�.���� sf�M��Am �cl�kd���ہ&�8���-�R��̖� U�M-Í� @ ��H��8�fZ ��U˷ks������*����p��UR�l�8������  ��2��Y�� �[t��t�[pH l�6�%��h
�s�l[ۭ[v�H׫� � -� .�Wiki~�[~H	��l�kA�  ^��Z� �L/@mJ��*�˰�.�6U����� s�	-2:�[��l۶�[h��$�
�*���+pu  ��H'gm�����,��آ��  �۶�[��fW�]�j�ɀj�Ș��� ��۪+��P媱��+[\�J�mv^�"m4ms��e�FJ����E�XrƦ-ڻ�=6hj�-�v���[z];�l��8b�yc�����]�x���k�:��bb��nE�x�gC�1θ����㤳uQ�nP`+�	gv �Q��"�J�箪�;=��k��[U�P�%�8�fmA�pJ�Uq�J��v��j[md��hon�9��Pz�Iڧ���-J�W UYD����H�v�,�-��m��m�Q�3�wEU��J���qT�Hl�  ��)�h��&i蝪ѝ�' �p ��m��m���ʡ�$6��5�i7l���6�D����S/��* @�[UP@v��    ۶���ݶ�i:g^� [@[G[CZ�%�IĎj�m-�l �e�W����V��k;]���e����  �Ud�l�m&�m���  9g�� �l�p����o��um�M�� 6Z  [\<�j���} ��*�l�����<��U�H �n�٬��re�lJK�m��.�M��t�-�٭�Cz�A�K��$6���R��a�'M�Y/	8�m��Hn� ��]sod�t(�6�A㝣 J�O�c��k������� ��n-�  ������<�]2�զ�X�Ҁ���ԒG��*m�����ul��H,s���H��{\�`8,��|OM��hd�I�{t�N�@ kX����^��jL�	:�l��H
��*�4�_	�A*���Lf�rm�l�=%��Zͷ]R-)���������"��`9&�^�`�`p�8�s��+m��K)�@-�@���h ں���s���}�hu&�b@ m��m�`8� p �k3 קM3� 8	$[@�B��Z��]�絇;7'<�ɭ�9���M�y���i�/���C��:lm�`�-��I 9m��I�  u�	�6�  H�l�܋m�6� -�m�iX���(�[�����6� [A     6���:���b�6�1����2����UC���T [����:W��Z��a4� 늺��aB�����Z��?��|���AW�bLT��[�c�sUR�/*V1v���R�kiz ,00�;kd-�`H �[�-���\M�$$ll(b�,�Zm�F�I��k3�m-�Ӧm�[CE�z��6Ĳ�       ��AmYm�$�6��m�kkm�$�h  l  ����@�*��ELa�_2��kl����d�h �\�` m��   pEl�7Z���H�j���� JԫV�+j����l�� 7m���  mU��      ���?B�ٶ   �`m��  9�K-�eh	W�Wq������/H�m�q�$��A#e��[I)�] �	����UO�CB�_�
i3H����O�P?��P�-":D>�U<P�(��S��ب�����B(���������c �F(��	 �ł�A�A���Oh@���N >�?�(�@>��P�(�@���
"��/�H�@�H B"��� �D�<���z�zJiTt�*�4���O�8���(�~��4P"@ة�G����X ��*< /�h
��&�\@`5�(���� ���HH�@�� E�Ab�! RH@�BbF!�����<G�I��b�`�X���BJ�0�B0`B�@T(�T�!"A`�0��,"��!�C���c�v) �V(AS�K	 B2F$	 �-@���%�?�
	ૂ*qD����	$~�ڪ:POЩ��O���()���P�((E?C�<UҪ�O�� ��v�,D=A����(��AE����mh�v �D"��T ��bF��*���*(� !�(�QV #j#_���              ٧-�֛Q��J�x�2�槅�[K�l�f��L3+*����̓@J���ufN�,�$լ�             $    m�  �@   �Ѷ��      'M�   m�    6ٶ�      $    6�$ޅ�����8��:@�Y�e�Ai
v��EgI�'(`�j��*�JX9�2ͷW�2�����s�:R��|�6��m:$0�\s� �<v8�6%������.�@.S�(+��Aa��2t1�:�ܑH�#D�ܗ�ܱz�q�Ld�6vT::L��T�w�q�[p�@r�JND���9B{v�6q���ѱ#��x�6+'&��[�e�]��܆�6�u\���#q�:w����v�j����q�A���NSڣg��F7^҉�L��z�:$������!��'N�`��R;f��`.N��ܕM����sÃ�ݓ���n6�v��˱n�áX��W�-�X�]�kv
�M�����'+s��l��b�T��>��J�q�±����l��v����U]�ä���Wr�ֆ;^T�NS�� "�:q�4�v�Sun'vW�8#��n$#uTz�2�[j|n�<u��v{m��q�[����e�Tn(��5T�Λ� £���:
�j�nѥ�9IW���bn\�0I�(g��v�VŹ�ݗ��0g@�@��!Op6���#�Ҧp�"ٹ���=˛lW$νr���,�8v�YM���<�.6�p�!�ٖ�7\��e¨ѱn۴&�뚧�F��&�$� �U�s��t)��*��Q�u$�C�f�ǰ�S	��R2�K$u���B/Jh�,KT����6�5 �B��lcR�6����c��.%�J�hV�8\�SS.fd�:$�3�P6�&' ES�uE�|
 @�	�6��)���޹�&ffffff`Xkv�:i��KL ��l�7j��p �C[.�,I�=�5Wkvm�M�;R�{��iη���{aM��K��i�,0w=P�u9ϴp�	�-�R���d.��l��nNN��3�����$���v���;�"�R궴��r��{q:��`B�nC��z[�ѷ\�k�^X/'�8�ժI�z���������{ǟ{���pw�'`A �x><&�ʊ�S*�)۳����lX��ٟ6��}�)�w�s�o@;�f��|�
��%0�Hh�S@��o@/����hu�:��a��Wkz ���<ݳ }��T�N����*�	�����@��M�Jh]����,�&D�EȚrh[)�^�M��� ��h�\1�)$,�l��ݫtK��\���ԓ�ç]��"n�e�����:���"r[��'��4����٠}l���w\1�Ě��5.���=��w����U!R�Rw�RJ�7&��٧ �za�<����?�2�� ��h[)���[?��~o@��x���E�mI4���/�S@��oC�f%���{��,܆�}ҚWkz}�h[)�z�tocPr�Z��N^�>L�ܑ�$�I�S��ҝ l�ܱ�<�&!cq%��20p�:�[��� �v��[0[L�MU�Jc�'�N7��f�����Jh]����c�"1�D�&����`zم(��(�%D(�wM�`����5x+�Q+��p5U'��|`��� {��7l�<��T�œ���p�:�[��@��M��4/b�������o�r/gϧf�A���.��L�M	,��:�-bM�����2�L��$o@/���e4��:�[�/\�=0�"mI4���/�S@��o@/����<(X(���ZWkzm*l�f��vi�;��ym�"Y,
���9�uX ���nف�%�h���q���a?�q� ��h[)�_;V���ށ�ⵑ%#��Cb�(�\豎m%]�휩�D�/$��^nv:\"�s/6�]\�F�D��o�e4�j�:��������@?Z��1�d̓!�I�@�v���ހ^�4�Jhgu�[��aYR-��ހ^�4�Jh�ՠr��fA�)�X����@����|�ZWս��x���h�jI�}zS@�v���� ��h�oĀ�H���Kԓkli�Y�� -���t� � �z�7,�W1�� [z��hq�s�n�v��������m��`��`gnG��A���z��ݻk�q�Re��f�yx3�bz�8^x\��pu.��Z�tu�]<���'s�,���X��wgv����6�Ȕ��f�z�N�ٞ�����ﯠg�Dj�����M������u�g��+�U#"�-v������6��[77�vZ{N�v�F�8��Y��Gb�7!�?W����� ��h[)�}�B��,F��Ӌ@��o@/u���h�տ��xb��(���	����M�e4�j�:�[�z�s"�̊%�4��>�S@�v���� ��h����L�2�4�j�:�[��f����/b��Лq���	#X���[(Z��u�ڢ�:�v�x5���W;.��)v,�EF��@��o@/u���~�IWXo�u�y��2�N(4����<�7�
$ �[V$��UR���IA
aPKw� }M�Νo@��^,za0D�mI4���/��@��o@/u���x*<�48�C��O}7_ ͽ۾ g��@��M���20qh]���@��M�ڴ��,Q��yS���q��v��tG..�Ϋ/-��j.<�39�CŹ�p�I�3��e��� �v��78:n� 7Z�dS"�D�&����hϪ�=��w����UUI��X��HʑAA�� �f�pe�]������J��f���M��cks(�4�X:n� ���0��`��!�d��Hހ_u���h�)�uv��}���7���M1�8}	σ�����YB�ّ�����c=�x
�y����x��	� <�jI�}l��}Қ��.��%��6p�yvKR�G����/�S@��o@/���e4�����L�4����;�<ݳ {��V��u1e�	Qܻ�j�o}�8�٧ �ޘp
."S��u�V�m\�+��V�rh[)�_t��k�= ��47����<w�VH��r��6���㇛�&d6�؀���x��
�x�y9�5Ր�$�_t��k�= ��4���=��p��2,���p�-vǠ�f�����Jhs댘�24b��$z}�h[)�_t��k�=���c�"@yԓC�g�'�w�p�o ̼�|���{���=���_���E����/��h���;�<ݳ �P�O�]�����Z�iYqu��	�+r@n�0 [@k� �8 -�:U���{*�mָic(��'����<q!���!��{X��۱�8�ǄJ6��F��F\I��^"�Nْ�eܗm�k����,k@g&������|b���Y�t��˷�5���q���^��ɗ��Zonw7���%�s�u�h��]-(؀�O�����/�N
YTଥ�\����eۈV�0w������s��d���&��c85�
2 �8����=�x��`y��5m!O*wST��� g�d��%J�?n�8�7�@���}�̊dC2(�Dӓ@�v��<X��w�y� y��X+�2�PPn��ڪI�z���ـy�����hUX��
��u5v�=�� �u�0��`�������I�C���=�R��p]'U��*�K#�,�:G�X�s:�������Jɛ��� {���l����Q���������=2 D�mI4z�9�T�MR���'x�6���ד�m�=)5$��9<G�
���%z]F�����H�)5$��_��K�DG�F���Ȁ�DjI*�;>�$�ғRIz��>�$�K�Ԓ_gL1v;�MD����$^���Kׯ���%z]F�����J��blm��R�3�y^�3��^�,v��ۉ�c9k�j��Msg���.��:���~������%z]F�����H�)5$����:c�#�L�B73�J���I%]瓽m�=0�m��=�]��*���,z���E��Yr#RI~��>�$�ғm��;=�%h��$R<	T�#i����2j����et�	F�i�C5��5�MWYB���]	���FU�2���(�.��0�i�-�s6f�4�H�#2�%�˦$tD!$�
=3��a��9!��~���8��6��,)Wd�BSI.���Oދ��#��5�M\�d\4i@$��6��|)ȟ�	F �$B,HR%ԅ ���*��7EB�J��a�!B��1`�e�Rc����T.* GU��LC�.��.�
��J1�#@ͩr8��a�\<�j�4n����Ȱ.��#Ɉd!�)t�$E�"���*cv(	���p?* x�� �LT���V��(��y���9�m���ٻm�Ӯ8����%r}�K�_��&�����w�����q��]�ܽ��m�����Y1b <�jBjI/z߳�K�t���|�K���|�Gt�ԒK��^
YTଧN�v�v��O�-&�O-tt.e��ù����o��秵��7�������6����'z�g�0�R��I~���o�]�m��2Z��m�IrY��U�v}����-���$����}�Iy��o��^�0�q�Q4�	�H���:��Ԓ^��g�/;���RI~v���H��\Ȧ�D�&�&��7߯�g�$�\��ݶ�u��9�n?�7>ผE���*�k�;Ϧn�m��/ӳ3,u�L�5z��3��m���
U�߯�m�6|MI%�v��Ir鍣�cJG�%�-�oM����n�B�5�v�r����g���DE?���]|B��Q�������׻N���ޘN6���3��UU/�$$�8�ߧ�������ct����k������>��%$o3ﺻ�����6����'{����)#��}l�Ƣi�-B��N6�������{9��|��I>���w��_��MI%��G�0P#Ng�$�bU������m��v���m��0�m�w�~������Dx�k�IL&�RIW�^N�������+�����o3ﺻ������>���{�߯N��߿�@���YwD�k=��K}m` m�@6� �< �$�lI*I9��	꫙�
N��Å��Kq$!��*�kW���cj�^�J���<�>��ix4������;7�n3
g�񀃭W!�q&CO]r<8X\��0����e�U�l�����t��}<�X�k�sg%l�<���9	�-�r-�]i�K�7���{��w�������,Q*�;�{�}}��r���:�i�0u�-��dx�7�\���痷?���M������� ��3��m���p6���oo2�w��e�6���a�e�r��&n�o���Ü�UO�RG��8m����ӽm�����]�o�ʱ�1��&C ����%���jI*���޽J����4�m��n�w���/<F7��`5B9�/ٙ������H�N6���3��m꤯���8�o��Qn�qu�M~~ o���u���{���K3］��͟q�m���^N����<�~��
YUyk(k���R8����zӄuif�I��{8��v�_�{��;��k���nnBu�߽��޶��L�8�o/޼���%����d�q�߽5=���%�	�浬9�m��{�7�=��1D�����E���r�����[l�����m���xs�ʧȂ"T\���2Z��m�DK�3����~���[l��{3v�D~`.f{�~��[o�϶o���.��������~~�;��O��`��;��零����Ü���fq�m�R���{/gz�f^#n+qX��uu�7m���{Ü���S�����y$�����O�I#�)5$�zb�8%#�B�XԽ��օz��&␤�N^�B�O/��f.�ƙ���vn���vx��l���%���jI*�]�|�G�R~��ϛIvf�w���^-!]�"n5	$�������꫻g�i8�oٛ�޶��L�9�3i^����Ddh�2����$u��ݶ��y�r���	 AD8) ���Z*�A�G����'����vn�o�{�w9�[�x�[-��!l�ې�m�T�/�䐊��7￱w���O�3����e��[ʪ�}�R\����q�������v�h�#���m�ޙ�q���_K�g����l͟�jI/w_��H���j&4��[]a��v�ɮ�;E�R�lv�䃃j��uŮ��u��oG0�e�	��fe�����~���[l��{3v�y�:��EB0P�RG�2��s�ٻm�����]K����fs��?y���� ȑcJ���7�}��޶��?��6��������_"�VC{ݟk�k\2�C.[�WY3v�{���9�m��{�7oȟ�1�g���}���{�Lݶ��O)�a�̱�L�Lְ�-�D�H��HU3{��q��ן_ӽm������*�J�ȥT!W9���w���k�
��.Fq��o�^N��������7��I/�����K�.�RIy�\�+	�)U^Z�n�v�e��Ӻ�*�N�t�8�7H�֝\��Z���
5��p���ˆBF��I"���jI.��}�I{����3?��\�����$���cCֱAh�nBq�߿g0�~T��$y��3���y��;��?za9�_ԕ/�s��Ͽ��vZ���n�޶��?��6�����޿�J��R���pߧ�8�o?��Ͻm�����"�Cn""\��m�T���̽��m�ɤ�m�繇z����*�\߿y�m���Yͺ����rw��~��q���%_{����$��?ڍI%�����Y��Gl�$�T�Tb��'��=s[V% �� �7��	���z�7k��!gf��qͷ����,Yl���;���;��)ٺ��ݎ��5�^[�{=�۶��W=��VѮ6�с�]V�2�cmk�����x[�#��tm�:�%I����Yz��q�;`;nŋ�۴#�5�,�t��Ґv���H����;Nr�.
�sn 6����֛�˩��k*"x��@y��Ԁ��خ�&�Z�8��S�9.���Kn�8W�Wb�]fe���2kF����A" GF��sQ��ȢQ4�<�K��������K��m����>T�`�B ��̶�{�LԒK���c��&c�2!8}�I{��s�T��)#y{���[l͟������ԕ/���Z�B��DB.
�gm���ӽm������$�RO}���[o6��K��/��"1A
d	��_�ʥ�}�N6���~}�m��8�6�I%��~���%_�?����PD �s&���{�w���*���~��Ͷ��o�޶����� ?_���+����Җ����K�܏X���u�e�PoK�a��gb�����~~9�i��a%$�rI~�?ڍA����;�3��U��a�~|3F}k��M�ra3Y�w$�|�^��Cj�P0 �]i|���)%�Ͼ���>8���|�UU�+�SX��_ͺ���;�' �}� �za���R���̽��{���^�#.[�2�n;�ꯕUU_���p�ߟ �������/�%T	U_��. {�_¹��
2�>��� �UT��2�t������>��p{�ˀVV\c��/g�#4�2����ڣ�&6����.��s��I�L�#�@�^ָa0��!��U���M�[��}_U�U%�H����ߟ ��>�),Np�35���9��vo�@�P�F(fO����������y9��_UP���/���������������߯��5I%@_�S�?3Y{�}��y��l�߯�^[�-K�q��|��J�Uy�ߟ ǻN�ٜ\�_QI_����f���%��r�"\���޼����U{>�������߯����Ndr�ۥ�N
�-����WDs�r�n�G��P��6��S��hz��۾︜��N�C5����hW�h�ՠyw;4��#.[�2�n\wܿc��J�UWf�����o��?fL9�I�����D�Q�q���|���'�I�n�Ɓ���Z�����`�ZJ�~����=�4���>$�\��"K-������;w$�����&�n(]��?fL8�T����_��@��vh�]�o���p��z4��k��kۙ��=��t��oZ#�m�$�sf�Y�j��rj̖�������=��|���'�T��J�TP��UHI!Q��>�|p��/�wv�d�K��f]�<�^�w�~"	��Db1Z���_f���}7$��ۿ��1!��UU BT�ٻ�ϭr+t7,"%� ��������>���;��@�Y�W�^�]\֬�WY������"��RRE$��U��w�{�޼��>_�� X� ׹���ܓ�oQ��qF+#�ˎ��;��p���*_�*UB���?���pٓ ����[	�sSO(��)�d�D�o
��e��!�,� TԘlN��e42댺!MZћ��0!Y�WA5��̓���F)-ͻѽ������Ju����E�.�t�ᭋ"HhSȐ=`�	4�	 �M�Gqd]��C`�aIq	t]o�Ӹb��Qx~d*�#���YR������j!m��1h����t�E&��'�@eD5[��M*jqO�I!Bd�0�r�Y����            �� ��(�b�]e�%��e�A�*4�d��hL�lT%q|���m%�H��UZ� u���t��#ol�            	        �P   �$m�       �l        6ۛl      �m     :n�u�{;E�9U��5����� j;���w�Ԭ��KMV�.	1@��.ڶ:����5l3NݔIҔ�I1�l���$X��.��k�ấa8Z�TΩel�jT˺������V�������:wGdOJp[x)��s���o/qq��;8�I�2���d;n�3c�b��#��;6r����)3r���ӛ]z���"��A|���z�z�oQ䒸�,�p�N�*�M�b�z�E.�����&�[��v
UF+)�F��n��oR&Mf�qă��n��i4���Lʄ�H�W\�rF��vSoF�����Yri�ݽ�p�P���]���jr�+-�����$��b���Ŗ�i����v��SN��`zqt�kjx�܄;�JVxs�p�P�/.PB�+��5m8\�fw]n�7Tc]aL�iN:sU;��c�[�۱P�iwl�kvQ](磅+����K�떌�ΰZ�k��Tr�x盧��{
d�ۂ�U�k��r�ː�@k��s��a�M�����<�V�ͪ�"R�\n)V�Ѡi��[<p:����v��u�£�F��틜��#�'d��O=n":�ph�z��}���vkuY�v�6�cm�8�1.��z���>(���Έ2�5�d�����m�c�9xl���5@U�ʖm�;N����X|t5�3ܔm\n��sI����NrŶ� 6[d�.�[���nۤ�`R�6ښֵ
/r�l�mJ�F�*�Kʼ�h�\tݷF�{�����ނ���+�S� mB���x �v���|A�.
=A6��'���䙙����kY��՗6�=�:�J�S5A�h � �$  �u�
��R��Ɏ�ƶ�N5��.^z�G�=�wn���g�Q�ܲh�݀܍��HmAxT���[���\r��(v��n�kl�`�%rkۚ��\�K�rr��@�� �\p*�5���p�c�A�É�=���ژ�s]�v��Sp�Z�޺p��wwz��8G��²D3�xy�Ԛ+�8z�PfCf���0��b�z�ن�����@�6n��5�05�!�[��ݿ�� �����?fL>J�]a�ri�*��7�0��A�˹ٿ�eR�U%�UT��O�g�����L8s.�	�3D��7&��e4�JpڪI�͚p<���??رFIm8�-�m�p5%�W﷿w���??z�p6�S��4��嗶��R�4�l��ɇ ڪ^����n��Δ��]f
1)���)���M�uN�ưӸ7�\��NĦg(�?�{�����X��&���k�4�٠}{=��Kı=����r%�bX��<-��]\֬�WY�ͧ"X�%�|�{�NC��H��!ZU.�R\ �A���j����Mb����4`��!�b���R
|��ED�K��7��r%�bX�{���ӑ,K��^���ӑ �U5���t�k5p�L�nMf�6��bX�'�wM�"X�%���fӑ,PlK��{��r%�bX������Kı/z{Mv̘3)�]d�r%�`b{�wٴ�Kı<�w���"X�%�|�{�ND�,�
�����iȖ%�b^��־	��Y��ɴ�Kı<�w���"X�%�|�{�ND�,K��}�ND�,K�{�ͧ"X�<ow���o��Lz4��D��0����K���7��$
�z���c�ꚗ�������u��5�B�m�2�k35��%�bX����ٴ�Kı;�wٴ�Kı=������
�DȖ%�����/��Re&Re-��_�2Ki��l�kZ��r%�bX����r*ED5Q,N���6��bX�'�g�f���bX�%��m9ı,O��u5�]h�,#M��!�])2�)2�f�NR�%�by��s[ND��hPt��ɠ~T@�A,!D��ER�P
�b�a�7���fӑ,K����㔺Re&Re,����7,"%��ӑ,K?�?�D�VW"w���٭�"X�%�{����ND�,K��{v��bX,EXDHQ;߾��BE:�����m��wnU��|T�R
_�2R�E���AD�D������bX�'�siȖ%�bw��u��"X������o䨬Q*�9���i:�u<Iԛ����:��WMb�y�ܜ�-[MLֳWSY�ͧ"X�%��罻ND�,K�{�m9ı,N���	�&�X�%��ͧ"X�%�~��5�5�04fS,ֲ�9ı,O}�y��D> :���'�Ͼֶ��bX�%��ͧ"X�%��罻NEO���T�K�s���0�hɓY��r%�bX�w>�Z�r%�bX������K�U��j'�g~�ND�,K���m9ı,O��JM�L��u�fk[ND�,�b'��B�����ͧ"X�%����]�"X�%���6��bX�@$�	�1UpW>T�:�����kiȖ{��7�������Rq�ZV��~oqı;���iȖ%�a���H H������%�bX��g�����Kı/��siȖ%�b_�/�'rh�U8+(F]�ck��ڀՉ�1v����fy��c��\ȩ�h��4}���bX�'��{v��bX�'}��Z�r%�bX������X)	�&�X�'�g~�ND�,K��Y��f�-��0��̻ND�,K��{�m9 �b:���%��ͧ"X�%���߮ӑ,K����nӑ��&�X�;�M}�Rc�.��ˬֶ��bX�%��ͧ"X�%��罻ND�,K�s��ND�,K��{�m9�7����n����Y�}����x�U�;���iȖ%�b{�w�iȖ%�bw��u��"X� 6%��m9ı,Kޞ�]��&��e��]�"X�%���u��Kı��{�m9ı,K�{��r%�bX��{۴�Kı?!�{��33335�k3)�Ճ=p��rn�8t�G -���  $  ��f�z�%V����8֦^3
�%��`�>І�P�y����웨7N�OYۜZ�ㅸ��d��On�?�]�	��Ɍ�5�:�<pڎX7�u!��lqM����j��y�F'�x@Sl��:����i5�ݶ�6^����v���P6M#��R��Hu�����S|k��	%n({zcj�j��s���=9MN8�{n��uuQK���H�P��/�/�I��K�O�ֶ��bX�%��m9ı,N�=��Ȗ%�b{�{�m9ı,W��M��&�r���w�])2�)8������,K��s�ݧ"X�%���u��Kı;�w��ӑ,JRe/_�j���q�[!.�NR�I��K��{v��bX�'����ӑ,�*���w>�Z�r%�bX�߾�r�JL��L��fY{n��,7.e�r%�`���u��Kı;�w��ӑ,Kľw�ͧ"X�*X�ٚ�K�&Re&R�ћk�ƛr�)����r%�bX��;�kiȖ%�b_;��ӑ,K��s�ݧ"X�%���v�K�&Re&R���؝ڗlwq̒�:Խ�'������>�oi�im���5�x�V��3����w�\��k�B7���w����bX�߾�6��bX�'{���9ı,Ou�{��r%�bX��;�kiȌ��L��Z�۽�mإܷe˓��QbX�'{���9��: mWl���'u���ӑ,K����[ND�,K���6����uQ,K��i���Ɂ�2�f��iȖ%�bw_}����bX�'}��Z�r%��Q�MD���iȖ%�b}�w��Kı/���5��adѓ%��m9ĳ��}������Kı/~���r%�bX��{۴�K�K�w��ӑL��L��wSE�퉨ܲ��w�]�bX�%���m9ı,;���iȖ%�b{����r%�bX��;�k��Re&Re/׉�T�7%ܻ��Wd�غ�H���p��3��3s8�ql���Yh�2=u���ҵ���{��7������m9ı,Ou��[ND�,K��{�l�Kı/��siȖ%��_�e������q�Hr�JL��,Ou��[NC�����'�Ͼֶ��bX�%��}�ND�,K��}�WJL��L���6���Cq�D�%�D�,K��{�m9ı,K�{��r%� �a�*�	��!�ؠr%���}�ND�,K���ӑ,K���M^�uu�]f���Kψ
��~���r%�bX�}��6��bX�'����ӑ,K��&��)t��L��_��-��F݊^�WSY�ͧ"X�%����ͧ"X�%�)��u��Kı;�w��ӑ,Kľw�ͧ"X�%����/~5d�Ƴ�*ƥ�v�j�6]^
�k��e'���vZ��M~w{��|s�����]d�~�bX�'u߾�ӑ,K����[ND�,K���6�Q,K﻿�ӑ,KĽ;~!�|Ʌ�FL�Z�m9ı,N���>.�j%�|��iȖ%�b}�w��r%�bX����[ND�	���b���&���F吗nK�R�I��Iľ��ٴ�Kı;�wٴ�Kı=׽�bX�'}��Z�r%�b2��ڵD�15�d%���])2�'{��6��bX�'����iȖ%�bw��u��"X����X�M�&�M�����fӑ,K�_��e�n��7$�)t��LK�{�u��Kı;�w��ӑ,KĿ���ӑ,K��}�fӑ,K�����Ï�^{�A!�=emt��/]�&�M��R�pٙק/C���+�s�>����붛r����JL��L��7n�K�,Kľw�ͧ"X�%����̀r%�bX����[ND�,K��=5{�Lte��9u��ӑ,Kľw�ͧ!�$uQ,O����ND�,K���kiȖ%�bw��u��"|
,�������߽�_�_K#���ߑ,K������Kı=׽�bX�'}��Z�r%�bX������Kı/z{Mv̘3)�]d�r%�`�'����ӑ,K����[ND�,K���6��bX$Q>��~6��bX�%���k�L,�2d���ӑ,K����[ND�,K���6��bX�'{�xm9ı,Ou�{��"X�%�ơ�}�߮������ߟ����  c���N�t�{e��� �m��6 m�@ ց�Y�ě��sUv�6D�ku	ڗ�s�n
Xtm읫e�ön�ƞi�Y�8�;��';��l���vS�t��WV��#q��-����mtCf�z���P��*�h�9�p�v��bÝ����ۙ�:��:3�vDݘv��z�tm�.֬���n^��M6�$�X������p��θ
Yq�Z��y�����V�y1�:+�H�֝\�����w���L�8�	�+K���oq�������m9ı,N����r%�bX����[ND�,K��{�m9ı,{�����gq�)�+_{�7���{�����?�X'�L��,O�������bX�'�����m9ı,K�{��r'�#�&DȖ'�������Fh�d�-��6��bX�'����[ND�,K��{�m9ı,K�{��r%�bX����Kı=����֩m�I����m9ĳ�@��'���k[ND�,K���fӑ,K��}��"X��DD�wﵴ�Kı:w��juu�]f���Kı/��siȖ%�bw���ӑ,K��^���r%�bX��;�kiȖ%�bw�����L!�]�y�Y�V".�亮wi,Q��;�]��F������=ݹ���������K�n˗')~)2�)2��o>9K�X�%���u��Kı;�w����'蚉bX�߾�6��bX�%�����d�љL��&ӑ,K����nӐ�!���U�7DA������~P���V	������浴�Kı/~���r%�bX����r*��E�MD�/N߈k_2adѓ&��v��bX�'�Ͼֶ��bX�%��m9��!�������iȖ%�bw���iȖ%��_�u5l���7,��ܗ|�ғ)0P�@����~���r%�bX�}��6��bX�'��{v��bX�'}��|�ғ)2�){&j�˖&�r��k3iȖ%�bw��iȖ%�b��C���]��%�b}���kiȖ%�b_;��ӑ,K����]�e��P���z�Yںs�=u�nx������%�p�r�qANLY�۵�V��"X�%���ݧ"X�%��s�ֶ��bX�%��m���j%�b}�w��r%�bX���Ϯ�kT��$�f��9ı,N���� &�j%�}��iȖ%�b}�w��r%�bX�����r%�bX����z�te��9u��ӑ,Kľw�ͧ"X�%����ͧ"X�1!3����1_d�!b�F�����"��&	�p%%�0bIV��,P	bR�`� :��Č��bH`��J�i�tI�iHH��Dp�"	H�P`Հ�I���BQR4����HQ �	$	R4`B����A 1H�@�ǊB�;k	v�q�R~^@�"�"���P��F-@��! F<�$�$XJ�C�MB0FC��"{�J�#b�Uj	�x����"~D�x�*z�ET|P=<U^(����.
���T��P��0D�O<�>�ND�,K�7�R�I��I��+^[w��ݨ9w	��fӑ,K?������iȖ%�bw�߮ӑ,K����[ND�,� �kϾ�6��bX�%�����d�љL�Z˴�Kı=�=��r%�bX��;�kiȖ%�b_��siȖ%�bw��nӑ,K���C���²���vy��d��-nL��6����i�bZ�u����n�.��ܿ��4\�5�e�~�bX�'�Ͼֶ��bX�%���6��bX�'{���?���|��,K����Kı=���L�8�	�+K���{��7�����w���Kı;���iȖ%�b{�{۴�Kı;�w��Ӑ~b������˖&�r����.��I�X�}���9ı,O}�{v��bX�'}��Z�r%�bX��{��r%�e&R��,�=-KA��r>R�I��~b���]�"X�%��sﵭ�"X�%�w�ͧ"X���r+�i)l���_@J	D��4�����4�Ō u�KB��"� D !�ɶ���@
"��L�{��9ı,O��룚�e�d�3Y�v��bX�'}��Z�r%�bX�� ן}�m?D�,Kﳿ]�"X�%���nӑ,K���K��%�U8+7���ƈ�G.��u\��.{m���0̉Z4=?w{�?w�ｯ]�ˬֶ��bX�%���6��bX�'{���9ı,O}�{v��bX�&�ݻ�.��I��K�ז��#wj[�k5���Kı;���i�#�D�K���v��bX�'�Ͼֶ��bX�%���6��bX�%�Oi��Y�Fe2�k.ӑ,K�����iȖ%�bw��u��"X |�Q5���fӑ,K�����iȖ%�b_O^�]�L�����])2�)2����[ND�,K��{�ND�,K��}�ND�,E�������ӑ,K���)��p�e���u�fk[ND�,K���6��bX�'{��6��bX�'��{v��bX�'}��Z�r%�bX���X�+ ��gy���gD���t��,ۖv�L���m:l R� p �hc.MNSv�d�֤ꎴw�O;m��Qwez�qJ�t�����mJ3��N����Ө:D�ݮc�ND :�׫��s`2��Gҳq�+i���g=>zr����t]�n£�gY��r��3͓�6�^����un�s[99��Sp��n�Qݪ��{���=�}�����ղB9��#���q`.���nH��xz��v�oD�0������w����3;��ԙ3Z�fӱ,K������ӑ,K�����iȖ%�bw��u����O�5ı/�}�m9ı,O>��j��њ��-�fk.ӑ,K�����i�DMD�K���k[ND�,K���fӑ,K�����iȡ�WQ5��~�}tsZ��,�&k3.ӑ,K�����ӑ,KĿ���ӑ,K�����iȖ%�b{�{۴�Kı:w��f8e��9s5��"X��T�My��fӑ,K�����iȖ%�b{�{۴�Kı?{��Z�r)��I���ym��7v�帋�')tKı<�=��r%�bX?A�{����X�%��s�k[ND�,K��vr�JL��L�����z]���[�6����͹(2*Q�f���m\qm��E�u=,j��'W4�u�u٣�w���oq�{�}�bX�'�s��[ND�,K��{��Kı<�=��r%�b2�ŏP�����pwr�K�&Re'�s��[NB��yBAX�X!!�I��0�*X��B�V� �D B�h#E�6ؚ�b_9��ӑ,K����nӑ,K��^��m9�T�K�~����njf]j�ͧ"X�%�|��iȖ%�by�{۴�Kı=׾�[ND�,K�f��JL��L��&j�˖&�r�L�Y�ND�,� !GQ=��bn	 �_���$�H���n&��'�/{��R�I��I��l�OKR��˴�Kı;���m9ı,>G߾��m<�bX�%����6��bX���L��])2�)2��Omm�wN
�Fy[�[����%[v:�ؿ��Iпq�]�-IP�=N1�Ҟ�[UO����{��'}���ӑ,KĽ�ͧ"X�%���nӑ,K���u��Kı:w��f8e��35�ND�,K���6��bX�'�g��ND�,K���ӑ,K���{�m9 �,K�G�u��[5�%�\&\��r%�bX�y���9ı,N��[ND��@����3�����"X�%�{�{�ND�,K���;��5q�5��k2�9İ���ӑ,K�������"X�%�{�{�ND�,K�3�ݧ"X�%�zv��C4f�MkY��"X�%���s[ND�,K��ͧ"X�%���nӑ,K���u��Kı0�w�՗�N�r l�.�9n��ne��G�tN�9($�
���5.��<:�A�P+Z�~�bX�%�{��r%�bX�y��6��bX�'u�{����bX�'�L�|�ғ)2�)~ɚ�2Ki�8�n�6��bX�'�{�ͧ"X�%��w��iȖ%�b{�{��ӑ,KĽ�ͧ"
�$!���by�|kR_��Ԅ�nS.d�r%�bX�k����"X�%���s[ND�,K���6��bX�'�{�ͧ"X�%���Yۢ�Q��$���m9İ ~Bj'}�~�m9ı,K���6��bX�'�{�ͧ"X��� �j���j'���kiȖ%�b|y�ƾ�Lp˗Xd����"X�%�{�{�ND�,K ����i�%�bX�}���9ı,O|�{��r%�bX����_⨬Q*�9g��.g�<�g�h�[mu!�&�b�Js$]��N��[6�]2�fӑ,K���wٴ�Kı;���iȖ%�b{�{����~���%�~��fӑ,Kľ�;O��f�9&��L̛ND�,K��{v��bX�'�g��m9ı,K����r%�bX�y��6��}���b_���5��,њ�.��iȖ%�bw����ӑ,KĽ�ͧ"X�%���iȖ%�bw��nӑ,K��ޔ�u8\�L�̷Z��m9ĳ�B�k��m9ı,Ou����"X�%��罻ND�,K�3�涜�bX�'�sޚ�Im5��ܜ�ғ)2�){3�r�D�,K��{v��bX�'�g��m9ı,K����r%�bX�y��&���j�Y�ہ�U���v�� [@k� �8 -�m�2��Z`�z�ք����ƃ����n8�mm�mn��&ӑ��܆�Ic��"d������ʏn-���c?�.����[�����.����V�.C˧�]��Z���t9M�<<�{cF֜��VSF��\�Gm$�A}���k�K�qv�;O���;���:u�;����O`��N
�Y㫷l:��;1�lԝ�-���Wi���AF�ȃ˱g�n�ڭ��ı,O���v��bX�'�g��m9ı,K����r%�bX�{��r�JL��L���5�}��� K�]�"X�%���s[ND�,K���6��bX�'���ͧ"X�%��罻NA,K�����c�\��%�f���bX�%�}�m9ı,O<�}�ND�,K��{v��bX�'�fl�R�I��I���ym��5w.Ȍ����Kű<���m9ı,N�=��r%�bX����5��K��j&���fӑ,KĽ�v�a�ɬrK�̷2m9ı,N�=��r%�bX��g��m9ı,K����r%)2�){��9K�&Re&R����Ȁ�	%n({z��NM�g�\����Ɲ����n��")zܷmpQac�w�Kı=�=�kiȖ%�b^���ӑ,K���wٴ�Kı;���iȖ%�b~�ҝi�L�53-ֳ3[ND�,K���6��TN����n�r%����M�"X�%��罻ND�,K�3�涜�򁪚�by��Ʋ��R�njL�n�6��bX�'��M�"X�%��罻ND������;�kiȖ%�b_��ٴ�K��K��W`��,�#��.��E�bw��nӑ,K�������"X�%�{�{�ND�,K�=�fӑ,��L���5�;e� K�>R�I�bX����5��Kı/{�siȖ%�by���r%�bX��{۴�K�����������ҘX�K��y=qX������穧bм���
�L��y��8eˬfk.���bX�%�}�m9ı,O<�}�ND�,K��{v��bX�'�{�n���bX�'���]����dDrNR�I��I���朥�,K��s�ݧ"X�%��^�ۭ�"X�%�{�{�ND�,K���;��&d2K�̷2m9ı,N��[ND�,K����[ND��p Sj'e�ȗ�����Kı;���t��L��OV�Wz�&�Kv]ܾQȖ%�b~׾��iȖ%�b^���ӑ,K���wٴ�Kı;����r%�bX����Zk��l�L˫�˭�"X�%�{��6��bX�'�{�ͧ"X�%��w��ӑ,K���{�|�ғ)2�)~�'��Nr]˻��x�[f󝙚Q����']L����%��4s���ԜtJk@�����7���{����m9ı,N��[ND�,K���n���bX�%�}�m9ı,W횮��jX"�G!�])2�)1;���m9ı,O�����r%�bX������Kı=���m9 �,FR�њ흲��d	$��])2�)X���{u��Kı/{�siȖ%�b~�=��r%�bX��}�bX�'�p��&9��33.���bY� �M}�~ͧ"X�%��߮ӑ,K���u��K�� ��@4���D����iȖ%�bxh����K��kS	�36��bX�'�3�ݧ"X�%���>���~�bX�'���]m9ı,K����r%�bX����R	M�gT��Dq�;^BuKL���a#�z�@�̼�::�Zw[Ԛ̻ND�,K���ӑ,KĽ�����Kı/{�siȖ%�b��u�JL��L��n؅w�"nԻ��k5��Kı/}��m9������b_��ٴ�Kı=�}��r%�bX��}�bX�'�{Қ.�2ٚ��[�3iȖ%�b^���ӑ,K����nӑ,ı;���m9ı,K�{{�ND�,K���Mas-)��ɖ�3iȖ%�by�w�iȖ%�bw]���r%�bX����6��bX�%�}�m9ı,O<Ζ�z�K@p���K�&Re&R���m9ı,>UB:��_�i�%�bX���m9ı,O=���9ı,O��G���@�� H�"6 @�E�h�U��FQ` h��
���BBF�����l8*HUMÒ�����80U�):w^��==��w{�~��              EJ�9�����Z����	��4�����f�1��ek#��qX �K(�U��d������                    �l    ql�m�       $�`  �    m�l      �m     9]�k|��Ҹ�
�D��Uۯppt�I�6K�s\�ɠp�R�鋀��i:��G�v�]�����X�N�N�>�]m�"ɑ�"�:;{*��
@��g�L�LbY�΍�������m�b\u>ʹ��.�{NY3��͆
���X�)�l�73��89vۖ��n��/v��V۱�Xm��G �=�qՎ���!��=v��=��R힇��f������r¹�� �P��笤l���h��Y1�qX�3ڇ�G
l�Tl�{V�
��[U֠�W8��v����i�MtMn:÷�Ȭ H�M�vݙwq�*gu�_;�-�՛4 G�G�<a Z�\����=���`6+�v��`��,�U���y����7SFw�sK�Gkr9�ݛGUP
�P�l��.6t:�
�;6Ț�;uI �M�є凎�cZx�Z��؃T�[\��v8�oGZѲ��C֣�1��:��u�v�B��8���6�F*�Z�8!el���u�p!N,L�]�Tv8��L� �F�]�e����U,��@7.Z�q�8�݇�5�l�1x����Wv�f펎D�.��4=nu���L�Y�۲֍�'lغ��sq�Vɡ�]�;t#*���s ��khց��m�7`.1)�Γl�H%鬹YX� �N��Zӱ�:��݂����F�j@ȳ�Au�X����ӹݛhJ�ۖ�� �7U�M4 �f�J�W"�NUtQhԫTҭT��d�Lɭf\�m֮i�!�(�0� =�@J����-Ƞ>!�L} �P=��B@������I�Y���m� l ְm� 	 p [@��Ē�I�]��8�@i��^�6���m��"1�V�ַ=�c�I�����s��̻��m*ԛ�[�n�qcb�9�P�͓���:5��][7G����g��3��s>�M���YG����\��%�.���C�3N+��ћM�X,����7�?ezPHr�-t����6�ͭ��h�:皆�n�8n.[�(��Dӽ�v��S��ı,K��osiȖ%�b^���ӑ,K����nǑ,K���o��Re&Re/b�+��Fڸܷ$��ND�,K���6��bX�'��{v��bX�'u�{��"X�%�{�osiȟ�j%����k��K�L��L����Kı=�}��r%�bX��}�bX�%ｽͧ"X�%)=���])2�)2����d��@yL�Y�iȖ%�
D�>���r%�bX���~ͧ"X�%�{�{�ND�,K�s��ND�,K����$��2��5��Kı/}��m9ı,K����r%�bX�{���r%�bX��}�bX�'���Ѫ�9�,��-e�qӳ/%����kvxb6������=4Ku�<s�7m�F
�m9ı,K����r%�bX�{���r%�bX��}�bX�%��r�JL��L��&j��-��r��fm9ı,O=���9 p�E�"���d�z�T �RA=U����D<uQ,N��|�ӑ,KĿ����r%�bX������Kı<�:]��I&&L�]�"X�%��w��iȖ%�b^����r%�bX������Kı<�;۴�Kı;��;�[�FL�e�����"X�%�{�osiȖ%�b^���ӑ,K����nӑ,K���o��Re&Re/b�+��j6���I.fӑ,KĽ�ͧ"X�%���ݧ"X�%��罻ND�,K��{9K�&Re&R�b|��ܗ��n]�y��9��v�%�s�	Z���;&�Ĥ��z�9̈́�Kˣ��ߩ��g�����nӑ,K����nӑ,K-��_�� /��h�U��$#2�&G�<��|�RI6��p76p{&�y�2I���q�uVhI�{���Є*B"�>����p�,z�`>w�n��R�X�#$BQI��3���[�~4�Y���ĭ��M����$kD�"�'&��e4�Y��Y�z�����������r��3�Js����幮�����-ɶ-��X�<����y��p�C���a�C�����U�׬�|����_߄~m-g�#x�$�M �'>�T����36i�g�s�l������D�8�jE&�_���;����H����_���Y���E�2 �N��7�p=�8�c����*�D(�
u|� 7�JwE�t+	�S	!��f�wUf�z��u��o�www���q���p��c�vy�4�rQ�n��_G!��i���=[.�������$�y"Drx����M ��4u����@��q����Ab�"�N ~�d檤��٧�Tٹ�Ӏ��M�>��)ő(Ȳ	ɠ{���w��z�4׬�=�q<J��`""r����n� nk����4u��:����̍∑�4�x����ـ��q���������$ m�Xƭ.v��n��WR�t� m���� 6��8 /��j��$M:cg�2�ˣ@+�R�6��[����r�,�V�.�ݜh�lA�I�u��.`ݝ�q�m�6��-���ݴ6�*˱Gm��k^^���{�vq�h^��o ���<wn�N�̚�Y:�u5´�YvϮ^�ї/f���`���_3fc�w��������wo�8��%�U8+^K�����Iɬ�q=f�].�h��l3#1�u������$rt7vp��qp߳'�U��M������X�YL��>�����$�l3۳��{8�=����2H��
,�)3@;�� �r��DL��X�x�WO!U**�dwp5UU&���' =���w�����7�ݜ}��Zj��8�cq��|� �%
7��^ }�׀�.��o����I	�2�7h�k`�K^ݩ����7���{Ȼ�;:��Z�y.>�{y���� ;z]��w�n�SJe�)��Y77f v�x�(���I- ��E�Ԛ���nI=�{��s�Jhh�ص�ȉ�"G$��+8�=���$��dӀ���;�Zo,���8�jE&�z����� �[4����g��d)DɁ$�����>���~ߧ��N {=��}�w����>;��� 9���F3Z�Vm�ɛgZn���:�&-h���\�5���uB��#m���M �r�@:����� ��$�$��D�$���Nj���~ߧ Ϳ�| �{' ��b�x�$�,S!1(���f��v���$�%��%IB �%+h�(Pv	.��$F1�Q�)��B��LL�0R�l��l�`Ą�@�")Id%��%����uVhs�b�,Y�� ����~������^�� ��h�%S�02 �#�@:��z�4�Y�{��@:�ciH�m��H6�廛��b�5,�!I��x{��AջZ�� z�cK�g�"b��I> �/�@:����%U�nl����56���I� �{'5*I��{������y4b�en�,R,��I4s�h^�@/Uf�u�4��Yc$#2� 9�u�4�Vh^�C��� ���=��I<=�^���D�H���z�4ٟ�����u�- ��h.��X%țm4�2]�Aks�r�v�j蜚�i����it9��"H��2�M ��h�j�g�jI$���׳�~��W���nY��8�^c��a��8��g :�4y�O��`dAG�u�h������ZZ"�-g�"b��94�Vh[f��v� �l�=���\Ic"�BH��fd�J��n��f�� g��������v�/n��[�I�}n H ��i6 /H  6ڪ�3��R�̣@q������bH�1�nۨ�u�� �6�yO8۸�,q�N�[�v�����L�:����+H��r�0f�]��^%���o�r9O\I�Ǐ^���փ��<=��d� ���V�\#(�������ƺ�7Fp���N��[�k�=���󻻻�|��WJ��Y짧3۞v3�X��l]9�d0v+��uvMzu��^�y�t������@:�4�Vh[f�}��,d��@Qd"��f�^�� ��h�j����L �c��@/Uf�u�4s�h^�@��q�FƑ��Rh^�@�;V�u�4�Vhs�b�2%B	ɠ{��@:��z�4�Y�������{'�Rʧe:���m1��gvtn�{R��x;<u�;vc�5b�����.�D�q|_�@/Uf�u�4s�hh�ص����"I$��\ߣ�B*�M ��,�����v� ��h�	sk.$�����I�z���Z׬��Y�{{+vAcp��I���u��- �����@:���g,����(��h^�@/Uf�u�4s�h���VLIH�Q��#y�^�Q�[<I�r3�ɓ3,��������aUsnl��,X�D�$��Y�z���Z׬�=�cH�
d�J)4�Y�{��@:��z�4���Ha�(�NM��Z׬ӿ���
��ެթ5YMiXGaCG�@� � "��(:e5�P�`�˚!i�MZE�I�v��#�+R扢�5�Z!� k+a�h҉f!�A��"B�%��V1Na��톁 `�ae�9��	�Z%֒j�п�2"��,`@��4�� 5"G� ��0�e5��I!s0֖-$C�0 �F1Y9O�QQ��A�}E�R�� �舞 ~M*�58(b����P<U *�Tɬ�|��'�{�nI��.īf)��!Z׬��Y�z����:��k�D�I�j�@:���)�z�������zSIy���~����ok;t��FT4q�_f�!`���\�`T��j$�O�/��h���u�4�VhŞ�ݐX��Q��$�[)����M�nl��^� {=����Y,���$�ɑHh^�@=�Y�z�������L �<�!I4y˼ ���nف$B�j"DB_���u�u���cH�
d�&���Y�[e4�Y�Uԯ@��*����)eU�����[5Ke�
tb�#2����6�����e�vY	�,i	ɠ[e4�Y�Uԯ@:��˱v%[1L�!����f�WR� ��h�M�QV��3�&(�$�@��^�u�4l��w���`߮���V[���K�mU7�͚�ߧ�@;����zb�en�%r&K��I8fL8�'�ݝ^i�`�w�bV�IJ)�O[۰��UT*@����xqy�c �� ְ  � ��[^Dʫ���Kd9`����p]<���t��k�G���M�I�z6�n�+q�;P���lB]�5��v�u���&u*-kaC.���㶹�7f$l\n�+�����v�:ݸ��q���UY��nk������kPr�A����f�0�4�]3Z�֭�%�[f��A������	M�l�/ע�\!6Bu�ڭ�Qc�n���6��n��/�ڼ뛳�[��1� k�%��>��������I0�@�D���*�W��f�m����@�[�64���BA�= ��4l��w��]J����$0�#A94l��w��]J�׬�>]��*�&�E��� ;[��1� k�z�S@��<tm�m&�cIbѴ��z�i�I��d��N��j���݀�b��9¤��Lq9&�z�f�z��̘j�K�������Z�j�q3Ys7$�����Q
mh�_Tٯ�~4����uVh�=�� �Ɉ��	$�:�M �[4�U���hݜ��HO�QdȤ4�l�uVh�Y�u���{�#�$H�M �Uf�z��[)��f�U�^:��JF�b7 �o��t���i��an��4�a�k�#���-m0c�MM"bB�"�M ��4�S@;���� :�_���w�8�C"�F�rpfL9�$�6���f�� ����J�g�jm���V�"Hp=�0y˼IRQ���ϭ�4ǖ�����.I�ڪT߳^� {��4�S@;������_���E&�z��[)��f�{���o�����#0I�]�]zn���\^Û��1L��vM��P<��g�u�KV9�"70$�@�e4�l�uVh�Y�vr�$FB",���w������z[)����28�D���uVhW��:�M �[4�.4liJd�I�45$�O׹��3vi�~̜�����?����N ���{��~�^t�Y$2,Da�Ǡu��޶h��4+���ֈ��bm,O�4|��\�;6.z�[\�\iQ[�G��a�y��a�l�B-M��� ;[� �r� �|��U��4��3n��(;.2K�py˼e���`kw�"dr�6�&�;�.˸���������bGz٠/�@�Y���LDnG�u��޶h��4+��wX�	�Ȉ�dR޶h��x��87l�=�@�`%�I*D!+Ł�A!D����F :"�	g�ߟ���Āl�ڴ��I6�˲զ�@ [@t��� p m�ܺ����;�^L�QC���r���S�n��hVrk���-�:ä��錽�A�L�Q�m��OF�}�]ۥ�<$H����a&oTnY��(��Y���
kq�W����=M�nwnYy|�fs�fn':�۞y�%ƻ^A������j�xc�~w{����S
�1�����ٮ\-l��卲��4!�8���ĵӮ8y�t�u�z�#��>�Vh���:�M �[4�.4=b  �"jM��z7l��� 7��ϔ(S&�?�\�أL�Qܾ��N {�dᴛ=��M����\9*���#�I��T�{vpٯg ���|ٓֈ��X��c���4?fb]/�@���Z[)��f���jF��QF}��㛺��H6��#�[��$�r'WK��a��u�*u�x���������@�e4�l�uVh�=��"F���ֱ˙w$��sټ�A��(*��� =�]����D$��4����"!�dȤ4���@=�Y�z��@�e4��;�G&!�ɠ��=_U�u��޶h�ȇ�2D$Ԛ���S@;�� �Uf������ɑ��y��_g���u�u��^ݮ�n�<^x�of�:��8)1�E��!�qhl��w������Z�J��4�0�C@;����u��M�;�hl�6�USfn�۱��(;.2K�p���ܓ���۸�H�AB�CP�E(I+9����� �A3�R��$����@�}V���hz٠Գ@�Y���(���E�u��޶hu,�=_U�}݊W�%^g,�э�Fʓn�<��`�6�buOE<�a�5�ݷ���������s���ݳ 99he�2ENM �3�#�;�h������@�n\&51L�d����S@;�� �}q�E��!�qhl��w�� �c��"!\$��U�Z:g�V���AC���8�<�6t���u���α��n6��VR�[�<�q��t۫��W��s�>�OGit�fN�z\�F���c���> ���h���:�M �[4�Ļ.	E1!&���������@;�f�س�[��91���@�e4�l��Y�z��@;;��d��Y2) �[4��h���:�M ��� &"d�4���K4u�pnـ��P�\B��LD���� M���I�]b	���R��MhBPXQ!R	@L�6] � -\F$!�RB$ Č!B0�P�%��i(B��fʋ͂ �bA�9���� ���*�&p��c$�FBd�)�6�"a�)ti�!VRi�t�JV���5<aY�l0�m�X`@�$��*�����dX�F�jB�\q��kZ)c!S��H$I�����Čh�@8��u�J�(@"A D�DHN� ,B0d����!���q<���Cg}��=��N�wwK��O���               h��6v��tM�#hj�nV�a�]m-j�%[X�ЖHL�7�1��r5Vq$�yW��C�m�                   6�    �z�        y��  l     l      �m�    �Ch�6��[-U@�g�1����$l�n��c�v8��)�e�:9"L��4��oc�QN��[m�`Ȯ�4��h͜q�Έ�ݒPü""�N�5A U���)�U���6�:!�G8�8�2�]�l�����NJ�t�ȱ���X��;z`��4�C%� a^�3���b�g�E���\�s��Ru�l^�!���ݗ2�q�(�&��H��7M��ۃ���:R��**P:�q���������#xu	{�{���{v�:�m���::�x��p��ke$ٕ���d��y�q��������L�q�[�ҰS��5�[[9�Y�]s�&�/ۍm>]�V�m�R�S� ۅg\\��X�]p �<����l��ʞ�M]�j�B���s����.뗷Q�b��);�[�9B�)���n^�k8�c���m��SZ�m��]�����t��i���c�v�[c��61�]��a�N��l�����1
gr��ʈ<��e�e*���½��gg�p%���f�i�� �9Ƅ��[{5d^׭�:h��'����g\vёUL���S�mp�۸��iu�����o6؛t����t0�
n�9 �d���^{Gn7W8��TX��n�&�q^������ֱؐ#�R�5�8����R����n�˽���k�-pnԷ=�Q���qT=���l� �m�와��.��,��� 
H�Mn�ҋl��j�j��V�85��I)5�)lˢ\��*����E�?�t��X�� ��PP�N�w�ww�������+��L�}�]5�ݵ� pm p�`�H��@�����M����]YɄ�u��7l���v���Ar�G/9�CN���$��sՒЪ����{s��9t�h�����s�eySٛ�q���n�˭y4�gm�EƎ4cm�9ǥ���n�.���03K���=���LN27\�<��V�)��Tv�Qg������{���倫�Z$�U6uyr�u�g%������vt,-҆�M*Qz�6�����&H�2M��hl��w���K4�����C��:�M �[4�U�����OLx,�0�C@;�� �Uf�������:�
����&8��@=�Y�z��@�e4�l�:�K9�q%��L$�M��Z[l�|� 7���?�$��u5_U��%^g,�s�s=��c>E�-�agr*��]np���:u��[�9��_ԓ7f� �{' ?{M�I%�����2�Y$eH������9)�T+aBQI(HP�Aa<���M���4���, ���(�rh��4���:�M �[4V��cS1�	�����:�M �[4?b�UO/4���y�����%��9�f v�xO1���� n�oo�����YN+qs�][�y�舓;u+�<cuv�j:�h�v�&;!��wkq$4�l�9u+�=_U�u��Z!V����#�h������:�M �[4�sj�?�0-TݗX��87l�脕�P�P���@�ߏ�@�Y��D������E���I��4�{vp?a��?e� >��2BfHd�ȴ�l�<������;��@���f���ĢJ]��o�Tvz#<Y��BrY����n�T$8�E0d�D�4���R���Zs�hz٠�.���"�d��/����U$ٙ{���٠yu+�>�� s�$b�C��=��| ����j�o�4����|��7��+CI�AIq�5$��n�睝�䟽מ���dD"�A4�(�.�Z^�KX�bc���4.�|U%U홯�f^���fN�ފ�nz$9%��+]n���[�籛GgT�oeڞ<�p���7Mrf��.��\���w������ �n��c����݄I��F��R-�ڷ���^��h����=_U���c$�fHd�ȴ�l�<������;��@;*�2�	�"ENM˩^��� ��1�6�y���<�V�+q2&!2=��Zs�hz٠yu���$�{������� l+�Y��n���ʓoZ�8m $ � �H  -�.Ň��j��d�q���ј�G�nIםbI�t�[%d}��9�S�'��NOC��v�R�;�웜������ݺ���lX.��Nv�c�c�e�O;������A��y^Ò��8�W�'��o9���zPD��vr�x�K��ny�r����u7[�8t� w{����wG�|���`��W�Lm5�N$�r��&�N����Z�fB��Vv�RG1�D�Sa\y����l������X{o5�ڌo]�V�)�!�8��l�<������;���J�$ٛ���e�Nˌ����?=��Zs�hz٠z�H�V�b�cR����;��@;�'j�$�y�� �ז��wq�.�E"�;��@;��˩^������x��l���qPR�[I]-�*�l��Zx�u]�`YznvΗ	�gf�,���d�ȴ�l�<������;��@;*�1�b��F��@��W��@:��B�!P�4`�@��ҧ��$D4[ �h7�(uT�4�" D�@�R� &0T��=/��>��5�߳'5$�纵
+q2&X�d�繷�=��|5RI�;��r���@�Ϯ8��葊a�ǀwSs�����u�l�u�y����#�#�@;��˩^�����ڴ��tm�m&�cIp�R�h8zr۳n�ۯ6�q\k�j[�����k���LBm(�CD�I�yu+�=_U�w;V�w���g2���LjB=��Zs�hz٠yu+�;{+w$q,���Zs�h���74X �@�t�$��!(U�Jg��� �M� r�N�DJ@�D\���Sy���<�M��U�w;V�vUF;�?�JENM˩^�����ڴ�l�*�U�駰Rˌr�Yy|�Ù�Ԉ��x�8�Mb���=,C[L���.5��;��X��8u78���
��K���s������8��jۚ�R_�B��͸=��<�y�9�<�'�<X�Sd�- �~�@��[�U7���3/u�{��匃-8��@��W�z��@�v����(S	��Α �u2�Ձj�������ڴ�l�<���������$��.�7Hui.np�p���)5˶N3��U��x�]t�VE�?��h�ՠ�f��ԯ@�}V�vwe��"?��`�Z/Z�.�z���j�ʨ�C	�R(�rh]J�W�h�ՠ�f��n\2cS1�a�����ڴ�l�<���y��Hd�C��;��@;��˩^����s?�����i��InI&D9��rɻY�-������ kX6� �8 -�	U�:m˥��U���fC����`�L�-����й�&Ƅ#;�l����]�3n�_k���Gf�x���<c��]ϳm�4�L�'d^gv.]9�^3�t�n��mv�S��B�IAHpC�e��ڭ�EOG����.�=����)+�m�T�sb'c{��3N^֌��(p���Ӎ5��t�KZW9����v^a2��6�F)�2G�?[�h]J�W�h�ՠu�ik4�)�@��:�5�9�;�����?	%'}HAY����cR����@�v� �[4.���=��H&Ƞ��j�p�np�n��n�u�pWvX�2#�@�&E�r��@��^������Z��,�m	��9�6\�[.�l=pu�n^�n� ��ô�1-t�%9�O�ґA���ֽ��Z�ڴ^��V��&51Lp���䟽מ��ȂC�Ɣm$P+A�
�UB�.t(�0꧳�l�� ���>JL�]�� ��/�0�Šu�-���.��_U�}h���<X��!�8�W��<�נu}V��v���KX��4�'#�@��^������fk���|�=��6��Y���e�JYT�awj���swRs�#c����v���[,�LƇ��ce��v�%O����ӀoSs�t�u�l�u�j��ӄ�l�	��Z�ڴW��<���e�6���yf-�H�*@�D]��~V����ޤ��*+ə	k.��5�㰩a0�%B]ڡ"@  $�������xC�� BEB18@�`AS��a������#?0`��F]
�)"�2B!��P_ʥ�N �C�?��!�� ��x�������%('��P4"
�������9�s.d�������ۏ@��^���Z�ڴW��[�x��LA1�G���Z�ڴW��<�נr��cy��D8���v��n�.������&y����#{5��-�x)1����8�s�h�W�yu�@����D=1��da�Šr�^��ֽ��s�hh�Z��"XӘ��=˭zW�h�j�9^�@�x#��k1H��M��ι��M�������f@
bE�S3�%�+�>Ş���16E��R-��Z��_��9u�����;݊3?d²D����9�l�6�&k��k��7pF��9�òk�n49g��0�W��<���_U�}�j��T�p	�R(6��<����������@��-���.�pɍLD����_U�{�ՠr�^���^��>��	��SaZ��Z+��^��_U�w\AS�,FF�qh�W�yzנu}V����I?h� BA��)Idc�I������?_�����V��I8]��K�;i �P l �7m�l� ��n��j���:c���ˣՑ�R칏.�Y,o�t��M�y�"n�X�Y�l���Gh�N����ݵ�>3TkB�/on:�հ�0GOcYr�7�N���zE�N��=�;m�ݬoo8d�᫱θغTݮl��7\�,���,c�9�I�X�Ik��}�����|�B�U8+)pg��q�:X��[.�#~�N���.�r��L6d��˜bICA�ܜ�>�=����Z+������#���)���Z�v����/uz�g��16E��R-�;V���z�������e��"?��`�Z+��^�����>�hT�C���)q�^�����>�h�W����S~�AЪ l��ۍ��TJ�s��h��R�i����4n�Μ�]c���E]�ι��� �|��
zC�_�@�w�8�C ���G����|@qV(Q 0U� S!�������=��|�UTٙ�����,FF�Z_��y{��:��@��ՠu�k[H�s�ǡ�!DB��V �����np�ΰu�9��$�&4�zW�hyڴW��<���[2�M��&�Fי�=��][����լ:Ӹ��Ю{`���Z�s�a�#s��H���H���Z+�����{T�u�m� ~^Ų�b�DY0r-����bG.���;�h�y���U&�to[6�-�.�_ ���`��	BS���؄�*��uh�W�y[����LA1�9���I����7�4�y��T���z������/�0�b�-��4W��*�W�u}V�{�W����nU8+(f�s��n��AXۦs@𻈀�1]45ƉƆ�N�b20�I������=��z��}�N�����dn�w%���{/�UUJ�3o5�������^�:�̒�ґ���zـt�u�9�u�j���q�M��s���}Қ+��~��n@7 B��E�a�AF��XDLQ	W;�8�ZwEڹ�%ʻ&��:_:��:�9�9��� �v���h�LJ]����;=�,��Y��]���v���	��5�פ(���{��:��@��M���
�ˆLjb& ���&���Z�Қ+��޶hs댑E_�a�Z�ҚoY�z٠Z��ۋ
l�x�@$��[�h޶h��|�J����p���.� �Nb�94�[4_U�}Ϫ�z��O;����>H �`�a�[ۥ��[����n H ��i�`�D� �@��"�mf���
wO�Il�D�|��:I齉�������)�����Xѓ�9�v^���ޗX��;sq/Kv�j�s��2n9�g"8��4֚�k�������{gun����v�PtogviAK�[g"���\j�r]��L4=��yvn�Z�B@b{n��s���6$9%��+]˛��=l����u�p���Ovn�X:�t�&l��L��uYI8����-�}V�[�h��hŞ�vbo�9�ԋ@��U����u������X�2#!K&
E�[Қ�u����>��hT*�a���)I8h��h��@��U�[Қ��p���LA1��M��hs�zS@>����������������i{<��&3�6I/
%ɴ��ZI�a·W��ذ�Ъ�N\|��c���p��O�UK�7o5��MkW�Zi�XAIq��ٞ�	b��興,.�� ����}V�ֈU�MӘ�R�{' ̿cᴒ��e���N��Cʚ̑��$����>��h���}�f��Y��`�&���O�Z���ޔ����-}V����[65�T����v6յv-t�g�,��]s��m�ٷd�q��9oZ&�p�ـ�w�7\寢[Aߟ� _�_�?C	�R(�p�{������>��_U�y[�ɍLD�Tuw�7\� =��J:%
A�(P�j E@�g��=��O?{�hW�"����%�8���h/����N�{�5��Mk\�i�da�@��Z������{��>��Ѷ%ډ�%��F�&=r1bm����ƺ夻8ݦ�6�F�8q�!1�&�Ĝqh׬�-}V�}�f�k�V#��$b&�h�s��w�7\� =�� �+WS��&���O�Z�u������bG��4ߝ����2L��EȒ�h�9�>w�7\�В��"JH�B+��*T(�AE^|��4�B�����R&�qh׬�-}V�w����h�yQK.0��Ng�r�Mhx���p4�vq9��=EF�=v�.5��;3_m�]s� ��xu�~�����x�O��P���,QŠ�@��Z��4_U�[qeY����da�@��4��h��@>�@�D*֦�"M9�5!�wY�Z�� ��d�jUI��4���cNֱ)jۘI�Z�� �u��)�^�Bp�}� �aI`�!F��������<#a<�c	�8t:d#!!U8�4bĕ�x�T�F���d��D���V$E4i��������#t����c ��$�T?���Z��d� ��(��$�2+`1���?�π  �      8    ���rQ�8j����SU��ڙeq\�)��n��;[�@��]&莀�*���h
�z�N�m�      8             l�    ����        �6�        ��      ,�    M&��n����%kX��+ӹ�ڇm![ӯTݮ�`��	P��a�S%�8`,��b�l�#=���u��]��
�v^.5��魘@E�ۃn�C�����VR�f�
�nqq��݁��Z�nx�a�ϻb3��9�"���ŵ��]n�&Ѵ�/<q�'aN#�vy�ݫlc-T;��"#]�N�-�ak�r�s�j�`��o���8��b�CI=��Q�&��;H��}u��U=��f��ڱ�=e҇�����X6����>v})�U�{f���7�k���	�tP��m�YR�l�5m�n��SvB1^�c�3t �rn�]��1�a�,m0��ɮ^��������z��/�6Yx.�ۊ]�aJ������P:�o� ,�=v7ee��9�d�O"�[�o[Q�pC�C�ս]��s�gi�%y-�������|�v��6�+];n��ڰC�t�<Z�tcl���A����Q��49]Vm���s�lê4�	f�5�`����1m琪6X6�r���X����Vqؠ*��m����sS)�1��.tO�iCD���[A��N�Kgc	ٓOiW�m��Kiؤ���vW����ڨ{Z5��ү���tn��ݐ�c�6�G�"�A�D�����!\�AaS��5�y��;=$zn��&�#�v��d9�]�[ݬ���՗e$�5� %՝�N
U���[�jsL�R�5�ڤ$��e � "[Ͷ�]'$���&.�Ըk��?�Q z��P |vb�@��x��@؞��{����w������ m�[�d�Ñ��M�9]UUp� H� � ��ܮItT��-Ӑ��Y�3XG���@�m�V�Z�wo�؊8���pu`��$L�b�&bm���M�FFq�v��ۭ��ܨ˵�'!���V�������Xg����ۢ�w]�z;;�a�(�{-���b�����������d��]-(q�po{��wz~���
`������ ���<\7=��Vx��a���T.nx�ź��H&��a?��~ ���4zS@>�f�k���2L'�"�dII4zS@>�f�k���hT*�a�ђ&�p��Y�Z�� �u��)�yr፩���c�����Y�[Қ��4�댑E�,QŠ�@��4��h��@��;��j$�6��9�{]8�Ӭ9���\�ܮ{'f�/0��X�I��b� �rh���}z���h{��:�
���ȓNbNn� ��yq	)���8��x}l�ʒl�dvZv��KV�A$�v�^ v���`�;�5J���&lW,%G#�jUT��6pܚp��N���ݙ���j�d��HF�b�h���}�f�k���4�~���� 9���3v�QX�]��^[�8k����5�7`Ě�F��&�p����-}V�}�f�oJh�ܸcjb&,&0QɠZ�� �s���`����	)�~����l�Sh��7W8��x}l�EQ��(��Š��ƃ?$�	FIU����pڔ�e�)Sr� ���-�M �����h��hh�G�A�&�Ě�����-}V�}�f�oJh�{MH�U8*]ɫz���&�Q��t���#<�a���D�#Lx�DfG�)�$����w;��gТ�o��9J���$f8�E"����ؑ���� ����k���2L����dB�h���}�f�k���4�h�Ɉ��I8h��h��@>�=���6R�"��D��$ 
�5(0]k�7�ܒx^ˆ6�"b�c����?g�b�f΁��N w���6��Ko6�Yv��B9㫰��P���oob���V��q���U-�خuIgn.�q1������4zS@>�@��Z�l���E�drh���}�@��Z������h2$Ә�R�����h��4zS@���<�̏S�4_U�{��-�M�uz�g����L�O�Z}�h���W����h�,�$��j�K8����Օ��%�-��� H�  � �@ܐFwO3�nj���\�C>�(8v�U�݃��c��gd�w!�pK(���ZH�I6�/Z1��%�����9� A�9)1$�w%����Cf�a;c��+�j�e9ܬ�Щ���A�n#Z�n֮�͹iM��<�o(9	��Y|�ձK<0-ỻ��s�eY"U�r�녝lD6�Fl;��1�s힝UqWK�f���&2B%�
I��Y����N�~��UWX��8��vlL�2E�$�z٠Z�� ���ޔ�e�mLA1�2NM��h��h���}�f��}q�F���,QŠ�Y�[Қ���UUT�fk��OF�����B�r`�� =�� �s� ��x�Ky߼�Rʧe,�ܻ��z�,���}��ܜ�.��d��˜b͓n�������^ �s� ��x}l�6�Lx�Tf(4�rh��f/��1BB!D�P���x޶`���=�=��$�n ��H���4zS��I���g ݼ����,�H����dB�h���}�f�k���4�Q�1�H���4�[4�In���{6p�L8^b�f\d�����o�A��A����4�fK<�SLӁ�����Gj����'�}V�{�f�oJh޶hW�$j���,QŠ�Y�[Қ������/�*,zdŊ,h�#�@����n�$TB�R�D����7]V�{�f�ֈTz4i�I� ��xu�pw���� ��4<O*3F)�ܚ���?fb�~�g�@>��@���17��&�Fי�=��.gp�s���j�p�$L�nFM���UӞ��,�BA/��	��@=�@��4��&�*]a�y��^ղ�q,�RMޔ�>W��-}V�w�� �Te�LF)�,i'�����8����ـ�h����h�dq�|UT���3_ 3ٳ�fzdܟ�N�H�@!H(���?�h���d��c�S �G�w�� �[0:�8u�p�(��K�}��)eU嬡�[\����V�z�KR�\��	V:�hk�2�c�[G&���0~�g�@���@�ڴ��h_&*<S$Ә��-��������h�ՠz�L<��A��N-�s� ��x�np:�8�Z��I��0��q�{��/��@���@��� ���&!�D�!I4���%����}-�X���U����������o���%u��.�&;i�� [@�� � �z�.��A-D���כnc`ں��[j�۲oIw��'U�RD�Wm��|�Ξ�h�!��ݵ����lF�{$)�[�w\l;{^6LO9
��sq�z9-/\�'�l/N���f���7g�a�ٻWc��y����Np���9�6⒐B�j;�C���w����履��[0I)vʽ���jN�zs�It�u(��Ӹ�e�E��4U�J��gVH���\~��*�@;�f�|�Z�ۃ���F��ŠU�^�w���ڴ���댎2����z��4�j�>���*�@��TX�E�drh�ՠ}_U�U�^�w����1Q�&�ĜqhW�hwW��@�v�g��D��Lj7�Crd�Nn���ϞG^gq�b���B�ڳpݮzAG<6"&��I��?+�@}�y� ���}�?g;�A�d@��#��Y�O�	JS��B��T;�� �m� ��>���^ղ�dq��}�-�z������h�e�D�⑫�����I?�����6���f�_[4e�o�	��D'����������������??��^߶x
YUyk4��>��nZ�Ӝ(��I�I�5�����k9ذ��[ɽ\���}�@���˺����n*,{#X�G&�}e4�uz]����hWɊ����J���==ΰ=ΰ݈�q�W;	4��$aBX��.���H�J���tJ�.�1f�U����H�HV!�ABCj�im�(hV�LHM��T�"T�?
9�6��I4�+i�FK?_ʄ���	 ��l6�\Rc6�)
����� �0�	���8�`���@�Łi����h��4�h_�_D� �+��.P��W[@"A��:P<��@)��4��	 $?"?�R��	)�ƫ�6SDY�{�2H$V"E����Y(�W�����
���L���qC�+��pC��B(�@-��ޚ^��=z&4:5���S��=�kz�u�^��>]��{9ܓ#1�0��8ހ}�f�ץ4�uzs�����Ȓ��@�̣�\�X�On;V�;��aX��%�z�Yy���&H�0��%�
I�u�M��o�{יw��X�6p|'��"�cĜ4�uzs�� ����Jh�n��	�r=��ހ{���Jh.���ێ'��d)#z�u�^��>^��>���k���qZ�,B%ЌW8
�e��]nI��/e5���5��drhzS@�{��;�����4ٙ�zV��6�j&4�'�V�h����4�6��[\W��0ɍƆw�����({x�dHS)!�]=��ހ_u�^��>��A���zu7U�y�ϭ��n��j�rL��8�D�z{��/���W�z�����2L��EȚrh�S@�ֽ�kz{����ɘL�cI8h�ՠZ�o@/u����?�?�<��I$����ˮ9퍂g�}�p� H: (�����M�A��h&��<��.'up��Tr��x���E%��k{s�u��s�{FA��g�
��i7�lu�j�0 ��y5ͅ�m�����4��&�z��W�<Y��t�<q�Se]x�y�5uZ��x�4"x�s��XЌ�)r���C���(k�����:�n�w��Ѥ�Rˌs�5�ܳdڲ�n����c�w'F2;OE��
a����a#YR/�����ހ^�8~ɇԕ%���|^j�e�.��,�D��Y�_YM�ڴ]˾j�l�jz5|�Kj�ےp��Ɓ|�Z����Y�}_'���Ģ��/��@��ހ^�4�)�}�B�(��"i@ƜZ����Y�_YM�ڴ�b�(�Lq'a7M8�.����s��9�.���oc���n��Ź�t�S����e��� z��n~J�>���� ;;�~��"!�D�&����������HQp�D.�����p麬 }�h�Xd�&H���4�j�3/2�����?n�8W��Wo�L$k"JE�uv�����e4�j�9u�P�2�L��$o@/u���h�ՠuv��{ϝ�o�l�/*>��������YB�ٖ��w+u �� ݧ�d������9u���岚�h����@��OG�)�5!�_YM��= ��h[)�}�B�(��"iL�4��� >�xB�J�D$�g��0�ՠ{<���I��D�z{��;�0���U$��u� <��b�2!�K"iɠ}l��|�Z+jz{��-�Q<Y[BmƢ�,q��7n�\����-�r�:1���r<OEW<\�2C&a2E�I�@�v���= ��h[)�}��mnbɄ�dIH���.���6���~ݚp�y��r��q1L��$o@/u���h�ՠuv��_\TX�5��mI4���/��@��oCs3���P�E�Ps��3rO|ו� SjC@�v���� ��h[)�{݊X�i����*�F��ůT;E����g��g��3%36��X��DM)�Ӌ@��o@/u���0������5wtEU�\D�z{��>�S@�v���� �z匓"!�D�&����h�1�ԛͽ۾ nf� g�?dH�F�n��Ԓ{��m���=��e4��፭�Y0�,�)�շU�������8DBJzy� m�9�$ݹdݥ��tζ��8 �`�  �8 -�8�*6����$�^��i9�e����Bstz^�\<tr�7k�r	��z뺁z��x�㙫<=����V�nz�1�q�٨�[
���2'v�9�ŸWں:���"����Z��}��G@�#��u�(N���,���.�;n��O/3t�6E盵��<����W�ӗ�I�C���=�0���s]m�n�������)3A�6�vu�9���Cz���}l��}ҚWkz늋�1dk ڒh[)�_t����ހ_u���x*<P2$)�5!�_u��:�[��@��M���9�i��8�䋁򪧛7n��?� �v��<X�Z�5weL7O�o@/���e4W��~�~����ar��*�9g���ζv�b�-h���4�k�],f͞.xz���fEȚrh[)�_u��:�[��@/�\2�&a2E�I�@����� A�QO��O{��Zܒw��4���>��6�1d�(�4���7U�y����x��j��,P�qA�r;�|���{���?n�Ɓ}�s@�mO@�qQc�&,�c�nI�;�0����f�t{���f�}qsʣbJF�m�JA�;r�v�"�P������$�<K���:z��=�<P �LQ����~4V�����>�S@����Q,FDҘ8h麬 {��7l��� �+S���b��..j��;�<ݳDB z
x
/�
nf����{�w���>�\��̊%�4��>�S@���\�y�|�J�7�͜ �	�f�&a2E�I�@�빠uv���f����V�h��qģII�T=����3��>�ⶸ�홴�z�E�i�S'�mfbɄQdiɚWkz}�h[)�_u��9u�P�2�L�ŒE�y���0��`�79�(�������,zdA��6����~4\v� ��4���Q�
)���С)}O�Ss�[�	�Q)� Qee>�#�"�J�-Q�CY�](�1�@�(A �G�@CZ���ܓ�{�:��a��\v� ��hl��{�4��f&�)�n)j�9g���N�}��un�ͺ��EMdd�n��sea�#�$�N?�q� ��h[)�^�M��� �:��ȚȢYNM�e4�)�uv�����USa��͂�H��p̚pt�V =n�7l�<��T�R�ƥ��8�O6n��}�8s&��I$�3�py���,P�qA�$��~̜6�$��J�n�O�n^��k�5��?���*�QU��EU�Uh(���H������*���*��
�
�*@��`�AR
�Q �EF�*�UX*H
�
�D�� �E��@��R
�T
�`�ER
��� �EB
�@ *��H*"�*��DB
�R
���@�B�`�D
�@����U �A ��@@�� B�
�"*H*H
�F
�R� ����@`**
�H��
����  *F"�`�EA��@��EE��@
�D��E *���
�����"*F�H
�`*T��@F
�E��AX
�P��E
� *��H��
�`*b*��A *T`*R"���
��* *��@"��B�
�
�V(��* Ȉ�W��QEW�tQEW�QEY�QEV�*�E_�EU�QU��QEW�QE_�EU�QEW�(�����
�2�Ωyh�#)������9�>�y� ���     T Р 
 �� ��       % )QR)R�PT� J @�QR�T����B��  �QH�� �   6     
Y� }�F[�Zrk��β�gK۞ ���퇼YC.���˙�g^�qu�ru�  g�Y^�=�V�< �s��s�s��j����š_�z�q5֕�;���b�ۉ]̶�� "��� ��� ��X����Q��jMx�c�����J��ul�W3*��om|�(��s;�(�:��g�x����Wǀ(�׫�����ǻ��.�V;�ko� �==9o�{^.�ӗuF�ݥx{�   �
 �c U}�ڜs�;/o7�@0 �)J�('J�bP �Δ
S@E)NpP�:R�((,�t  ��)J1���PH�R���JR� ҖYJPX�)Jp gJR��JR��J)K1�)�M(  �(  � ���3�)Ll�(�vtN<���t��Fw����=�y���۟7:�����g*e�������y4�7�K� yR����Y�u���=|x 7�,�sMv˞���w��u���(    dW>���m�'_-95;9:U�������m�=�*������s�Y���_.-Jd׀ NZW^�g���B�{�O.�ܧ�U��Û��������A�����ק���;��G� 4�%)P  "��i���J��  O��J=F�� ��T��)J0  S�BQ�R�M � DHCRT� �x�ȟ������X�����_����>�K�}�k�PU~e��@U�**��PU�����"�QT�����H�ptA�F�����2�g	�4]f�]oi����x���a
bL��S��.k�0��7�
p�!2XB3�r�S!��.���
>nBz�$I����Z�i	L����S�Լ��{��akG>���y_�3\p�K�8g=w��$|#B5�X8E�� �A
��Z�#Z8��
����6BZ8Ė� ¤	"k�BH��
aT����d���P����Hd�Y�)cH�V[������eˢf��r���ܸ�Zn7AlRi��!۪i���0H% �"�au��d+�(H�z�:� ;'�]}>��f�E��!a�9�v꣠�Wf��tl�qS=u�n�x:��<�c#�J$M�xH�k��"B;a`��Ƹh�e,bT%H�Hi����ܦy�e��S�����=e���^y��<
f��\K��CF����<�ad��e8L޶z�Fy����>=���=��B4���wxn@��֌yFQ���
���B8bJ�K�2HH�3V�h20$�_X"�Q4ui6����x�>Sq$�I'��M*(����jje�x�浤�h P��@�#�2˨kR���L�oCL�.B�Hl5�!p��l��$�!8o�7�SEޡq5Ł
��c@��0�˧e�߼7�>���P�$E�DȐ�}u?GE%�+4�>;�+$�
a���Kb�2��$JB�`F1��,%�Cd0��]�lی&��u��34r p@��ٰ  SDJ���Qs�PL9�qЂ���8��A)p��q�H0�pB�I�E�`H�F�������\%57k)N9䘔�̆K�:���!��
]቗ZJVd2d,�����ʊ`�]�4$hd�AHƤ�-�!n2������b�X�H�`կ�	�$f$da)"B���	32�AIF�澘$�O�� P!dCkBCQI +��� F��,���+D�P��J�B�������)��f���|>H�jo�s���}�1D�	Ps_Cxo�̅s#R�hU	���ŗ.��ī�Qq$�PƎ.�377H�j�����6{�a�3~r�0�y�Á�p���$BH�����S��6y�s
���o�:
m��J�Ɛ��b8�rA��ja�4.A�\%1��e)�P�bƮi�8$k���B���`��QOj�l�S�wϾ�h�f���b_�P������4�9���?�p�Ǉ�{�1����a	��S5�q�<�ۣ�>!~G���H�XHB1�����)�tC�x�#s5�k��Ѿ�NG6]���05�$��.��ˠ�\8B�S$.$"GLB+,�RsX��[�8rf���伐�-4<&eV�d�i0h�T0�J��d� @��Ӻa�^M��ph�4L`CE�l�aP1��8B��C+�6L	p���2_P�G�"F(a��EC5y���9��7�&za��!�4z�!Lt�x��|g��m���
da ��0a$ �`�,���U�u�<=ܷ��J�цs���<����,w�؞� G��F"��M@��'tv뼮K��bDCUw�3���|�M0�$i����'��\����N�ᣎx�� ���^`Ȑ�4���h�i�7����N�:N$��h6��
��� #��c<�����0H��{�5�Lk\HP D��c�p�ԗh�m0��)��,
шHHF�"�HV��bP�Y+��jU�1�U�:�+��>�w��|�:H�����R��J�v�Ԑ��?qq8&�g�B��O�HA���P�K$.:���0�LRE���h��\�sA멆ѧiL0�$HK�5�&����t�L�=�~R�t\ɩ�9|a���MU�WBX�5�H~ƪA��W�鞮|�y����TH���3����vS0���2�2��bW�Z0"�@Ʊ�̦M�C����q)�S�
y�7�5ͻ��y�)Q�t�#
SS#S�H��4i' c�D��$I�&� y$i7�ǉ�����3 >ICi�L�x.�l��8��ܤ����$X���]��5�igz[�!;�mO��p�Q	E�>�q0!�)��`o��>�lӴր��|<O��>���8r�1�y�k7�1�t��!��'���i<q�T���,)��Qs�I���_P���ԈsV.}�F��Д�XN<6y���.z���HD�$�F)H��sĀFr�ӽp�=��<>�@˜�yy�{�g�|��0��<$��O�J0�B��)G58y����7��x|����h�����H�ŀD�0bE�R(�Àd��������aCN��Ă�x9��6k�FF-�F�E�F�1�{�| &��"@0�Y��\SA����!kf�$��C��0H�"b���G��$�!��D���0��V:)@��H�X��Vbd3߃F�	V@���R�d�	 ��8���-���R�aSi�])��"����x�!@�5�#���z�s�s�y��))�D#)��$ƞl-a��#A0R#S�)s(h��4�$��J�Ú5L5�ہ�$R��p�a|���6a�� ��Tم��L�����i�]nÎ�2%4l�����<�l�kf��F�H�!�p*F	�����F�^bƸSF5sg�Ӱ�b��@"5J�
BB�RL�BB����}8'�����!���0<������9<X��9�zJf~<��P����2�|�{d����L� ��HŰ��b�<C�ͮ��H%\XID49p�ӋBAjڸ����H�Z3~���2�$+��
'����RD���/�Έ1.U�e�&�A֥kiJ0��[H2����p��eفHjR�9$n�xesg\Y���35��l B��B�J@�fn�Ԓݛ3xpHS�!Ln��s�
�/��#Y�Yvġ
����&��ڛ8{
2��k�s�6�p�܁������<߄��ta��D�t���D���H�Y��F���#F\]M�iXS��՛;k�*�?fת�6�'�T����7����SR)k��9�f��uϟ1�����}������+��LIR"�O"25�N�:x8�.��8pB5�FÆ��c�.q6��ӵ �c�C0���� B2h������+�}�.k�,.H��
K7��㞅�`��
�I�J��1!�)4�)�"��4�I����0�Ri���9Y͞C���ٞG�XIy��4B�l�|s=͹�SA��s�y`���9�4a��4D$m����{�i��盫H��䅋 R�B�RB040�8i���j����]k��RJ�t�b�` �_��$�M� k2�. h��5��� �л`��m��$HI���H�ץ���se�$��                          �                                                 �`                     �                                      �>           $    h                                                  �                �� m�  $�@                                                          H        ���                 �                         	m�����@ ��  ���a�`	m��m��:ؖ�ջ	2	 u�  ֹ����`i6]6�`$�U  K[�5�u��sWCm�v؜c���3��`ؔ�۞��ۊ�ܐ8��&۬�m2q�l]L6���5��@
�UUR�����,��S���`jU��		9����[%։m<�򓈓m��ꪪ�$YPZ�ꫫ�,2� 6ٶ�ٛ�f� H� �[pZt��L�֠��L ���}��6�  H$-��:5�np��-�m��      	-�)D�	�-� 8 ���m-�׉�PWl�����U۝ Ā A��6�m6��� ��tٶŴ� ���m�  �l�  �`��^���,�*Q_+�o�m�nצ��lf� �[�� %�l��Լ�h�.��v���Ŷ�"@����޶�$VyM
�^��L�4UQ
�Bـ��l�cNIxuJ[�c��\Q�V�gNKm� 6���[m�S��)��n"�3,WWn  �`ږ�� ��W�cE:D䍵�q��Uj�]���6�q��:���`x}:KD6�Xt�ԫUT�R�����՜�.   �d.��,7k����]�f�e6�ew@⮣efu;(�I�Vݳn.ݍ� �@*�^YVW�UR����i���-��Y�.�+)��L�@6��"���*�*	V��*�l���}��pthQ�U�펖r�U(���]�|��gm�*���n{,��5l�6�1,�d���RC���Un�]mJ��PlY�mm l�mkZF@P���m��V�B����Z��x�Cc�(�c����j�VS���cnZ�ej���媍9`�8�V�@@�y@j m�n �4��Z�r�m���ԫmm+� $�Eu����n�*�iĀ�d�n	;*�R���P@��a`�����&��*
��Z�,��:)W/ ��9�|~I�l��P "Z����:��`H8H-�ͭ��i%\�L�mm�4II	i����6�`v�p-�:%�"i�6�m[Rf�6�꺕@�j�!ګhqm�&��-`Mz� `��z�>b}���$86�p����$�s�$�%��i��}��|�ʭ]U��L���W �[*�U-�lʵl�rNjU�� d��zG1��VԫT�0L�w-+UR��v�@o,n�|��u��݌s����=�:�]�!��(��/Vt�rn�)��v%���c�un��M,�t�=3d�r6e ��IӮ�Ƶ�iS]$oA�ϕ��U�*�kivZ�8*U3펻R��im�M�6݃�WM����d-���(!ͫj ȰAN��e��-���b�8�m�$&�kY��m�[�5(�i� �Iv��jm���{M���n�d	n뱲� 	ڶ��I�F��[V�h���ٶ�m��6���ѣ���kf�: �m���ԅ�mm��� 21a�6�  m�%�[I�j�gm�j]�N�YYP�8��   [�� sm��   �F^6輫V�� m�K� /[��   C�p
�U��u*��(�V�"�@��h��TD��L��m�lm�A�l��[v��m�/$� �a��`X��I�b�n[�n��l�����v�N�ɧKp }����t�;v� �c�i�n�7m@Up�P6�u��v�E�P�-�FӦ�ۢ����`.�`�(�T%KfV9�lsR�Sӈ
��m�
����U�~j��ap^�l�Uz��,{��� ��V�������*���H;U9�A�ۍU���gC�U���fNN��E�6���
���/!�`f�
q���6Cf$wϜw��h�i�(�UAㄙb�u���k��8�)Yf��]����I۩����z{*VO�Z���&�Y3e�M�����\��<�֣�ojj��T��r�Q�e!�&�ml��Ov�Y� Z�k��X�nnͶF�m���@��ai�@Uh֑e�7WnI�����E� q��I�����-�65dC��6X
�RY{`n�k׭	8[�m�Lr�m���KgT��5([M����f��	���q�ְq]�I��uHp*� �Y',n��k�-�  gĵT�a���\n%al�t�K�nBF�Xa5��ϴ.����=*�V�[��e�ٹ� u�RUJ��/-�E����Ib�av���V�;[�q�P;ས���6���i;I� nv����Ivi0 zƢKM��m�vµD�rU[V8f�۞�mPPd�Z����lP2q5UR���l�jvu���x8��[�HMQ��Ԭ�J��m�m�lΐ6Yғ���+[�YFٶ$�`pH �ʭW]J�*�*�:��S� ���m�f��փm��M��� $�I�-��|[d����a��m���  �Kd7X���!�Dr��0m��ѕ,K��3Pn�U�8[nA���V�jU����]�e`6�*�
vdSJ��El�\� �]�4.܎P�V���U"�Z�h]�8 m��HS�\���B����J�\�=/l�iWjĠQnl՛` ۶�f�6��8$l�$������-���A! �ؐog[( I&�&�c �U.�;J�U�Ab�n8� �F� �ʴjjU�ԡ����$���-�m�:	�3i�U�F�x���RZ�k�l�6��Lg*��٩�Z^ZU�z��ʚe@ݚ8݊��re\�j�RZS%J��U*��m  8@88 -�"Kn�)%	-�$��� kn��:�    6�  Lݷ$)�ֳ��Ѧ�ڶ-��m�۶�  6� $$6� m ��H �ؐkjͷj�I����m�띰6�8_,�r�  ���t��� ��d� ��>>�6�]3�j(]��I0�����ZIm�A���m���Ѳ�qm  � l���'f�,@49j�4]ɤ�ֶ�6إj�6���p���` ��m��� I����-���h6�km���  �m�  �\m��ݰ�j�ۦ2C�  p7�l-�e��'6�ml���	��iWH(-c�D�ݔXi$X���V��i6�8 �����yU��C�)-UU�=����뀩r� g�6�Ɛ�H�m��on��K�j9G7Ͱ[x�F�NQ�5D��۞�ݠX��jXe[g���u0mYv�@�]ڶn�M�%$����[~ N����km�Ie��7M�{M��]Si@[TѮ- �8  �'N��6Qw^�D��Yp.�]�A��moWʹ�6Y+v��� �`����
�  �[[V�L�UK�U��r�]*��4�j��m5 ��t�m�Ò�����m�`$�B��*�*��i".�m��I�|Z�/Z;!�v��4P   ��l�ڶ:�&V"Y�4Fy���Nמ�j��
�E8���<��:�Lv ��    �  $ �`�h  �`i�Yv�l�t�   m�e�mp֛0 ll�v6؃[%�R-��Cil [B鰽m���e�  6݀8�'A�H�[B@ ֱ }��|��p�m� M&� ���kZ��
���(
	���h�A����/�"�ࡰ�G��>"��C�Zo��SJ��� *|"��'�ڠk��I$bb����W�>1U��F���T<R��h��� �X��Ra�W�h��-�U�('�@Z"���#��OGH4t�s�Q���TÊ؉A� }����� pa���Bx���}d�HD",���"$�āc	,���`A���"���E>TN$@��
(B�!�IA"��cTj�A@�A�X�"�`� ����1`H		$)��"���0Ă�1I��D���@#Q *D��F
1B "�� 0��b�X� ���.��B+�b��(�Jʎ�`AVP��V A$����Sׂ�l *#�5O@������!�'����
�G�_p|P�Z(D@��T}AN����hA���5�vl`@?���G�P^QH���{�����o֝�W���P��n�\�Z�    $     �    8    m�      �� 6�-�            m��      �     X`m�  h    ��S�r���zaj�<��[����zրѕP1���l��\[<�s����i�v���UɹmRHi�9MUP
F@.zy�m
��,�	�n�j�ħl�8na3���=�2��r��lci�ԙ��[	�ݰ�����m��X��U�{@k(ymΪ��d�v�����-�1=�0�i�b�������v0��
��t���\���70��K*V��R��,��� A��	��p�F��Į6��ن�M�4R�m�z�ͭ�s�5iۑv��:J�NK�qk��
X�n[I���8g���xՋ��c���[�Qs�������<�X�;��8+۰������Q�t���� �S��������CM��15�Z�fp��:3/����=m7g�#�az�۶�/[�8܉��E֋���s��Li�<�s�n��nKlaڌ��]i\=]�0ꬮn�TLv�A.��xsK]r�V/%ۢۛ����u��{��m�����[G=���Lt�+�9<��Q���6���o�8�p�B��� �{5�!Ӷ����͌�qnʆ��)�gnQ�گMa\�x��j�nN��nJ�D9�KN��&�W+<Z�;!�ţum�c���n:������j�XQț�UgYi�q��g���Z�$����p�e��eAˢ�b7kg�s�=T��wQk��	�`H�2t����9�+�;m=w�k����q!�js]��=�ݬ6\�j6�<�Ƣ�/TJ���i�p \窂�l��^v�����]ӯ\f�:Jhշ`&�t�t��M�-�2D�e��܆��TN���{����w��Hd~|G�Z �zA�"mV
5F�����kZֵ&��kZ�� �sl�ΐ �lp	9�9]�A��÷Jn��Fg�ë�
4v����n3c��5k�H��[���s8S^^��qv��<�g
e͸��mX�0����{\��5˴Im�m�I4V���:�ч�����m9�rK�'�7��ct�@�[�Ԓl\[��EN0�/3�����������=��|�����;�=��y�^rvq�.^yN�L>�˓)�	�&�ưi�V�yW��;9�n�p��&T����K-,��=��h�)�r���mz�z6���S!s'��4V����BGLoRH��Ī����4Vנx��@��s@��M���FF�'1�����٠Z[��wt�����:�S��	�Dk3����\t����GZ:h���9���T\�7�I��F��18�@��q���\�0I1��J]%+,XM��4�������DB�߾z�w�@��s@�PV$�S&BJLuE�י�`�ʳa��vՁ���@/u���HF����@<��BGL��0:䉁�)B�%)R��I4Kw4��9[^�_m��TJD��~2G�S�<�J�7ڕ��j�m�
��f���cdmAG�3��L�I�`���Jh��@/����� �{f\LP���8h���/dL		0'vA��TJ�G�8э�$�@��^�in�����	$NWk�3&�#牘����)��UM��n�X�ZXy�6/mz���n��&(��Nf�{�rD���&���t��0�0�@5���Uϐʝ&�p�Y�j�f�:z$YM�ܼ�P=��θ�o�:䉁/dL		0'vA�N(��Iӟ���{k�--��/t���ڴˎ��y"jȔ�`f���k5$�l� ��Ձ{�Y)��9���^�M����1���\���oRH��`���K�K`K�BGL	�)�{x���l�5���0S!�lp���C�vʹ�	��}$���b��ƈ���m��Q,m�$^��z\�s@�ҚWj�����.8FLDM�#�:Ԏ�� �褶��07�K��LN
0qbs4�)�uv��mz\����bLɌd�)����D����wd��9*�UL�D�S�1��6�%���[>4�ՠ{z����$� 8� $m��6 t��۵y ۘ鎜��7Z�&.:�{' [�]MvH��Q��J7�thN/���x��N���k#t�v�:ͳ��Z��Q��a�99���9n��h���vɮ#&ix�N.^�k:���mq%��3���Xٸ���ke�z��
�kvq��e7dc��H�SKܑp5[]V��/O�߽��|��"H�rI\l�SNCc\�m���e^9;y�n���Y(箎J�P�q�*�m�?w������:�V�_m���D1\�T�R���`g{X_�l͝�`�ڰ--�����a��҂�xㆁ�Ill�����wd��Y"j%���@/������Jh]�@3�ޫ���19$�@���wd��&Ɍ	)t�1#lmV�l�bS=:�n����TlS$n:�ڬB֥9Z��[�h��J�����;���>̭���0�7mh���_D�)�ɈRWj����j�BI-%4�
"B#���.��aܵ`g{)��:���&F۟��h�٠Z[��^�M��h�U�X�"q���@��s@�ҚWj��@���+�)iI���^�E%�	�cBGL�pV���%�/h�C��ή1ky�n^�L\)�p$��-+�L����Y��6�������������ER�k"�MD����h�٠Z[��wt���ڴ<�긋���I�		0;� �����������@��Ս܈ps�d���ҚWj�-�@�����&
@c&!Hh[^�ym�R�h�)�w�%J&���D�R'�HdF�^;>א�w)��"��:�g����2��N�P��&Fۘڑ��٠r�٠wt��B�0׻�`b�+\��USsJ�L��`u˓ݐ`K�&�&0;��*�HcJLi'&��ҚVנ[f�ʫf�_{f���ǓSE������`n�X�y�a�Qp�~|�i�{^uy"h�nI�������	rD��˺�ClhnCf�l��W��&����u�mxwm��K���3��u�x�6�q�*�ʹ��������.H��"`l�.����`��@�빠Umz����Z�9�
�����s9L	rD��������8Gr��(�T��*�U6P��wvl�{�`w��V�{;�6-R��h��)	��=�V��빠Umz��z���~�Ƕ�
d�I�2I�L��$ @� ݶ �� ��I���9�N4&D���H��M֞1wew��Xs��
S��%7 �W����H��6��<�Ç���[��Wc�v���k�藞˽��dyɡ*K����H�r��@�+o�v�[���l�7�t��Yg*��j�3�mv�4���*]�[45�Ϯ�ߏ{޷[���e�%�dMcbÜ�ۤ�t'd��`ȱ��<a�n(�-�˜��&r�D�4��$��:߷4
��@�u�@�կ@/�f\CPjc�$�fM�$��盳`f�ݛ��-XW�+kp"ƛ�G�x�נuw"`ott��$L���\�a��*�����ԡCͧ�6s6Ձ�3&��u�@�����CH�z���\�0=}"`tW"`+�ܼ�-A	Cӹ�y�+�����`�\9r����۔�W[]�^�C����u����%���&Er&�GL	�-5*QT���UN�l>�M��!RP�:+�0;z:`K�&T�TDJ�˹"�$zV�z��s@���Z���D1\IHcJLbN=�빠K�&��L��Ll��EE�5S9&h[^���^�ի^��u��=첉H�Cj9��f)�!len���װ�n�Χ����9y�b-M��8)	�nI���^�ի^��u��*�� �?{X�#"2&���[̛��-X�2l>�M�B���i��!����8�����k����lN'��L��� A�dP�XAebWec`���j°BB4�
A�X<7IM!�'��چ̄�3#�$� ��/��pK��u��
ń*�F�4���bFѠE-� C=!0�
,P�A��:7�f�RR5�c@�.	��VcPj�c"U��D�VcR4X-4��W	��i�B�	��0�Z,+
��3F�P�ѩq�����B.!���(c�(0�I�3Z!%�yLX�XPaHPr5$0!�*,1��3���aM�P4 kkD!2��VaLB1"���A���	.h@a���s1T�H�Z��#ʔ�Tę��4��,�b@�
$h��U��} ���E���A�D�̸1�	`Bp�3���s
��0�,B�1L�0��e�\H�XZ �U�p]�N*��"&����Q��}O�8pT6�JJ���d�d����V�r�)��`'3@���Z��Z�{��xî�Ǐ	2	��)�����{���"`I�)3����nxg�S��q:�uzM
�[�w:s��=�U�D棷�])���S�c��{���"�U�UW�6��Ɂu�b�Rғ��@���h[^���^�ի^�_n7�2���K*�fe0%���&Er&�GZ�����LL �rH�Z�~��ٹ'�����N&���T�_���5O&]�D\�R�ؕ��L��L	]#��"`ܰ�íe�jH��[�����!#�j�%j��D^ώ��]�5�ݗ��I�hͫkvu6��Z�1�d�}̝���3e�́�<�>po�1���h[^�����{��⎎��*3+K)e�&��L��L�0%��s��+��G�G�ujנv��.H�s�`w��b.U���ۚ$njl��j��I$�����{��U[4s��~���[�4�q�$� 8�[@ @6ؖP6�  	8�V�s*F=�7��wk���lru�۳d��mĜ�!���o3,�.�tk�en��v�x^<��es�#m8Gq��t=#pg<�vh�G͵�Ѹu�XL�N�n�vc^���GQ���m��K�4&Z-^��s٣������g,�[+y)XS$5��Q����Z��35t�2�w]sz�ln%]���n��Y��9��w=3�;fb�H��CQ�19�]�=�z��V���s@�[H��I����;��w�f={�`wwmX[^�g����#Ɉ��-�Vcd��䉁ܤ��R�(Rd��rh�w4
��@�v��V���po�1���h�d�2�_ ǯv��2Ձ���<��F�c�>j:ɈJy��l����mΜ^��/� �Σ�鎽�C���`w)-��.L`l��\�0%oұNKeSu46�ꝁ׏2�a/�BQ�vf�-X�ݛ���{	%ٝ0��̂I����}�ۚVנw;V�ʫf�u��0�F(�s%�M+P�$���́�;���ǙV����>�Z��i�1�)˙������`yyHK����]~�j�Ǚ�`}���!j8���e�^n�^Mؼ�kY�����˪t52u %Uly	qLs�>2h�T�S)���~~�Xfe�fO��+��w��X��2L�!�NM�m���������;�eX����1�����k�;��M�F~�/$! �X�"�*$D +F �B� �X l"T%<��~���ڰ3�;���ER�fi:uSa�	BJ<�v��`k�����3-XzD/O����Y����T�f�i���x�*���� ׻�`w��h���MH�CqHa�GJf&9�w,�u���՝��S<����l��+��o����%M$����4
��@�v���|��h��m�|�b��܎f��3&��&�������U��fZ�BK�L���/9M:�:ARL�UM��z�Xx�*�owvՁ�wf�����EJ�ʙTXl<�{�`n�ڰ1�d�Ll��4�>�:�΅*�T"I�5Vfe�V��� �����ǙV�Hw
,�%c5��Uϐ�x��c[P�K��JzzLh��e7~����77�ip{�6fV^<�����V�����0� ۘ����M��E_=ڰ7wmX�2oT6j�J�;-�N�h��\�`c׻Vfe�<��Jg������Ł߄v�&A4�n�����b����wf�����b#��y��`��m�5���j)3@����м��o<|�?z���}��D�n�	 Xa�[@�l�Ĳ� ]6 I�+���[��f�A��t=�br뗒�:��=	6�6�rs�&�g�L�]VN��sm�{S;`1��؆ݚ#v8ܻ�UҳX��.�5�{�t���l����6��֠���n��a+U�=@����=nsv��	��ΪQw\CF��T�6�k��v&�_o�}E� 5���;�^��~�{����?�u�p����v8r��z�6��́F���N��n���5�S[���H@ BpѾdx&LO1�$��O�h��h�~��O�H�B$b�`0�<��M�.���4*�&dQ`{~�}�����F,L���lܓ���6gk؈�� ��DDɞS�W�*�T"I�5V���`c�ɳa%�I!$@�&}��?z��+��5.�Վi�4nN��R��_�zl{kŁ׏2�6!x��!O���X���9
�D��t����a`jIFN������y�6_Lo�u.�lQ�%�=�v�g�r-�G�6�M��e�j�hƹdo��w���~!�F#�m���ڲ[y��.q��r�^�(I}T����s��f�Ӗz����rۚ�n�~�߸s���(i���~�.���y_��m�߽�q��8�)ި�Q3-���O��Q�<Ƣ�<�$�O�ԒV���=���g']m;m�����6�J�Y:0�4]k&f��eݷ�?�P����{~��6�ϝz�������{�B�$D*���Im��ůS�&��Rd�Iu��[o���ڻ���C�@F���������%����Üm�⬶2�"�m���9ױ�<��ۮy��f�d���v-B֥9[���������_���뛫hD�Nj�Ͷ��{��m��˒�m�e��!DB�i���^�m��)o��&�S"j�.q��s.K��K�
"����~9����S��y��\�Jf^����I�m�Q8�I%��oǞ$�:��R@���D?���9��������o���z��CT�GH����{��Z�i�m���.q��s.Km�DL��4�H낉��A$IGI9����3�m�н
=~��|�o����o����������G���������v�>ru��8O�h�r���ԆT:�
����������c�~5��5#�ܒG���SRI[v�x�\ꔚ�J�|�<I*��c�Ɋ`I$�����y�xs��&e��ZU������m��T��Jf[k�'��
�LS2��o�ҭ��fg8�D̽���$��}�x�J㩏.Ls$`��V�Ԕ/	*�{���o�޵6�o;]����	$E$dE�EH�0�"h�XA�ZPB�B �R �����jI.�/�8)�L��s�ng�$�<�Sm��J7/5��m��ZU��Ͼ��������_)PBE�nz5��]�ܾ��P9��q�C��nu٬��D��?��w{ݽ�䢤G/�NB�Q34�9�?6�����׎��m��fqyyDB�	DG{M�?{�? �}����j���4~~ O�aW�!B�!$�US~�{��m�����ݿ{�~��TE?TZտt�W,�d�A!���&������g�$�mܚ�J���$�U)5$��n�Q��Nd����6�Q��B����m����o�aV�؄�<�"QU�������Y����x�1L�$s&���:�<I_��	�������^�m����r��̵V�n��0"i&�8���量/�@�!��J�9[�)��������=$# �����`0�`��z��0�C�C#σ�)� �X,�a�c�\�(�$D�ѫ)H�#��m<;0dIZ�J����Xx�ͼ���`fU%|29��7���%t|R����	p	Lf8\�Ӣ�^.��Q�l
�,.�.2��&m���Ed��!�©�!4��Jh�X�)JJT9���`{͡!���f�aq%��HA���K���������v?���m�6�yP.RP��v     $     �    8    m�         l�             �     �     6�     [@    9��%��t�N]�R��-����������5ɗ�2�M��$�뫖�Щks�{u�5E�G]l���� �l�.݀��m,�����T�-%��M�UU)�<�EAܦ�D�=�K�[u+�w	����N�;G1�dګj�p�L����L���8�M�&,6쁬Yvс�r:�0v�����^7d�u�϶P���{,M,�c��k=��3���L�}Q�:�&��8KU���Jb|���:(pnv%�چ�m�Cc;kh[lV\{#vu6^�s0�i��g�<[uj�8�Q�4�b�۱��zc���r[��I�]C6�M�1��t��x����@ݰ�� M�/ �BG5l��\k(�@�m䯫>I 2Y��-W����I"�<;���������g��&�M�ݏS0�P��٨��nv���ɚ���c���;�.�ײ�#E/=�����t�9;t m��hWx�v�۶)s+i��ʅ�BMp86�y'�zqA�%�'����m�Z]N���٪�Z窃k���Bל�u���� <���"��'N�G;�P.Y��xys�@��<v�g�n�\�lvr�v��t��۱Y�쭆D됭�&̡�J�^5����m�X6�Ի�׭��v�m�{`k�h]ȫUYKK� ��ɫ$��������q�W�p�<J��g�j�c)jK��{gDc+;���=��eA��EJ���<C67[9�ݭ�+���3�œ��C��6��\FN�(6�9Kl�OW��eԆ���ш�G�v�k��vF��ZM�[G�f�uX�v�R�IZ8���`x�sY��2D�m����V	�se�;���u�_
�8�gAh�mQOPW��X�@<?(,Q�����{���~�?Z�`8�[@ �@ .� � v��/Q7	��բMiS.L��Ϸ$w>�	z曄.m��%a]gx-����3�9,���rj ���S�6�k��f��gWO<�Wwnqg�u����� �<��u�8�涳m�a�uRd��]�s������]�Ls���b����Cq��œ��Q{#�i�e�`��kLm��wﻮ�����z�(c)��.=�u��8z�	8>.9����Ŷ�kM]=�9�������9.>	z�+�������� �����l��U�"!re��Y��m��u�+U)�T"i�4M��ϳ8���P�UT�{֪�m�k|���̒��m����s���L��s�ng�$�mܚ�J���jP�fwd�&�m�wx�����hNB�Q34�\ҫm�Q
gk3g�m��+I��y�g8�؈R�w����څKQ������'N�y��̒��m���7��/�I#�ܚ�J����$��P�GӉ��󣵅9�I��]��q�µ�<a��Ө�����k���o�b|;Z�fܙ�� }�}�y�I�ɩ$���J�J=I$�ۂ�%TDo�Ԏg�$�mܛ���"$��#�<�p '"��� ��"��஀̦ݛkFR,�RVP.L.�8�(��(@da�A#�v��!�6�lqR�CP�󜷙�?g9m��&�Lݶ��3���D$�	%UO�ʽ4�5%'H*I���V�oӻ��o2J�m���L��w��m�wmU��k����˦T�L����y�ި�S�E�6�o{���6ٙ���z�(�����o����*�M*�SDӃ�ԒW�|�<I"۹5$�}���I_���� ?��C�HZ� �[�f眯��m�6\�A���/Oju�ݗ�}���nm7Ht�1MC���Ͷn��y=�O8�}x�
�Q	yD(_U6���8�~��M9
�D�Ңf�[m���'�Ԕ%�%UO�μU���{�\�m�̵V�KˆL�Q�#S$Ț���IUT��m�y��9���x�� l���倈�H ���* @"* ��� ���" �b�7�M���[���}���[kΧN^���Mۚ*��%�$�����o�ع��=�����y=�O8���Q
<�D$B��s��m���5#g�+0��.��9�m���5m��A�1{����[o�μU��ϳ8���}YX7T昤���qz�Z�E�6{��y��x9͝OY�HJ�ev��Z�WSs�:��37_ �{��6�<u���}�ű	B��6���E��k�O�j[�T�3%MT󍷓���ԔB�����\�m��j���O{����wwr�������]]���m|��w��m������$����l󍷳�������t�TSP�is�����BU[�}E�����y����YN�p�F�W�^��y�{��[ol'{��$֍3J����m���<�m�G�%�>z��$������$�݆����jQ�4�.�ysB��]��-�WvL���]� n����8��q̍m��W"S����_i�m��3��m��ˣRJ92�����h�.(��H�pi'"ԒW�|�<�""f[�ۢ�m��l󍷓���ꄔ�I^���L��s���ĒW��J����$��X�$���3�J����5%'H*I���-��Q	Uz�}<�m�|����;���z��3����m��ߧ��!=q��O����}��R�_fo��m���m��=�O8�bJ#ߝ_�e��   $m��`   E']t��N�5������ݫcoon9�^�����=�m\WeoZ]ml�u�{aN뭷T����M�WJ�v�VI{#׷Y��bVr���x;rU�������WK۲��qPb�D�ۥ��� aXȱ�۳`�0
�i�xb9#iCl�n��C\be�7.�f��}����:H֢�֥$\k��cW:�8t��m��5�.S=�L�rpN;l�1G/WWV���?��f�s����t[m�O{��?(P��(Df[o��u��=�����:�b�NfiX��W��y(I
d�����:�`y�w4F�ŉ��nc��x��nI��]}7?�O��)`)
A��{����~�`q|�fK��)�)U*su�ܝ �1E��b���ן�����nI��}�ru�� !dP����X���o��i�4Jnh�=�0;�t���D�ړ �&��1�/S�ճz�wmu�t�t�iu�]ɜ��8���d�5���ֵ��F@bGY�&�䔪�9�5N�|�j���rl�ea�xP�����;��Vo�ziJjJN�T�USJ���rm/�DB�D(�%fVٙj��s-_�K��B��$(BJ����?�j[�T�3%MTܓ�������߶n!����X����~�`c��M�uf<*�ҪUH����`s��V{�j���rl=䈈"AH���s���~��}{���fM�*��f����Z�=	/D	@	"�R*{���y$���_��<��>�mƠӉ���d�X�:����.��ҭ��^�t��7<V�8�U���!&F���s4uz�l���u���$E�H �  �������z\�!MM2UQ.�l��k��S��H@  �"�BJTg��Ձ�~�j���rl��M2�"�'�p�<����*B(�@�D��� �� ��� "����$(Q7׻�;�u��;�&ɔ�&�k֦k.�nO��?� "����P �A�����U����6َ��9����.i4�i�����V{�`yDD%��$QH��P��AH�1 ���<|w}j��̵`~�ӎi�tU4BDa��v��r�s�ю��ڵ`w�w.`�.�3��2f����ʐD��  �@)  0��̹�[�4Y��Y�����:�X�rՁ��j���rl�1�T��R�E4I4���Z��?(��`�@���(�S����V?{��f:��%�B_�B$(�`�R�S�����ff���b�NfiX�~�j���rl�a`s��VX����!UB��U.iX{�"0V$R ���f�~�u�nI�}�f��l����} �?�����_~����)_�K��)��J�%�Kd�����I0=}�06�������K�1l=�8��r���s�hv�L�ls\cdmD��������˿8��;%:m�ۚ>���`ffZ�8�ܝ^B��{μX�d�zJ��:�j]R�33-_興I�癳`wu֖;ܵz�B�%2o��sLM"�T�USJ������%�H�WT���"J�#��}�}�ߍ�~��33-XjI�9�6�u�T��R�E:��wGL	$t���D��VB����!iG˽3�&����*���� �`��%� m�N!�s]lN��*h�mN:xh��9�v�	nKmd����ڼ�l�}�9A.ۛ6������pa+�a�����;��C���kpӂ��"�z,����mc/�7�;�ܸ���K�h��G��-���8��6ŮvɈSmfݮna�E���x��q!q���t�K%��Ҧ�ur�
�<ӷ!��n�'']C�\��1Ls��O]0������E���LN2LM���}���x���-�)�y�w4F�ŉ�����ӊ���ro�(J?��*�߿*�X�~�`ffZ��%�~�U�J��\�!MU7*��U6�ߕ~,w2Ձ��j����6��<r�R��nh	SE��x�$B���=�zՁ��rl?B_�?!	!$������`�ɲG���u)�SSJ��#��tL	%d�0;��-`���H��rV�8 m�Z�j�r�✧;&PL��:o�R���"BPW)s�LM"��UM.����6f*���s-X۹��WeiȒ��6��z��lC��� �E�)���`�TC���! "�au9���=������ߔ%�BJ�BJd7���iU*�SD�J�,�j��̵g�%
}y�6������S2�\Ԗ�r����T�V(g��|�{��3aa�ٻ�`c��Ӑ��I�S.iX>�&���G��P��P(^��<|w޵`w������H�1�!��v:��4����s`�9�U�Nݝ-b�,P�,�s�R5ۙ��D���>�U����Z�;��^J#�BHBP$���}6��.|��N�s@J�,w2��#�!	&�j�����@�ܔ���Cj8�� ㎕���Z�>}�M��BN�@8��I$BB$&��h�q�+$׊���
�%��`T�D�$�CA{� �P��(��UaQ�|#e�Qp�IY$B�J��+,�M���$�f���@ F0�&���7�"%�B(`��(�>x:3� U�_�@�T��x���
Gx,E���$;��f���훒w1e�&�M"���M+СB}�͛����9��V��"w}-^�<ӑ%	�m���m�Mηs@����=]��庄�N(�M8�o%���F^jۋ&B]��sO'G-[j��[������Ds�|*��R�
3R�����֬��j����?�D{����_�_�7?�J��aw�eZ���ޑ�o�&�����s-^�^DɬFo�d���35S_����ޕ�`{�t�ޑ�W�Vd��!:�������l%�BA9�\�`w}�V�̵a)GRI�4�}p�uD"����]�Z%%�R�i�"Q�1`�.Z��BKn����;�ܒp���\�Jt�d����̵`~��o���{��@��Jh��u71��ɍ��'�A�GL�O*m]���+ɝ9��d������EW-6H�.���uD�����zՁ��zVA������U������njiX>�&�	/D(�3|�Ł�����=�w4;/2��IBbdr;��,w2՞Q�"!"&s}�V_}�����#�$"!�qㆁ�fZ�>�e�����y%"!	No�<X}���cy1H�14�h�����ɰ>�*���s-X�)�!V�����o~� �À�-��$m��` M��x��ۻ,��2g�8t�xuGr�;맩1�FK/*�.��댕��	֍��n�Dc�i���9Nle旬t�����c��9ʘN+K������v�)�`�j�wj7N:��P]aN\nk!%�A����P@Jo3��4px�5X6p��,���N�βr��k5�ן����Ǥ>��z��X^�N�Ϯ,�l�;E�<�c�ze��������ݻ�������ʪ��:�_���6��XX�e��$��;�����[�3T��2U���������ݵ`w7mX>�&�DG����eϘS�S&��4X�����Ҳ�Qt���әN���T�<�zs}׻�=뒚��s@�.��~s	��I������P�����fm���Z�<�*�%"q��c�5�2?	�Bo�?>O�����h�x�֞Tq�i�9�h��Y�#b�?V~�:�}U��6���L>���I�`�x�y�vn�GqH� X�$X�# �	 AY!HD��%䒉Wd�2Ձϧ1�waȅ	z!*�~�3+�s@�T��Ұ7߿Z�9��;?7��ZXfm��G���.�P��C��aſ�m���^,w��{ݹ�g���܀(� G��qV�����~���߭X������	��%�NM���|�
B{%�;F�@��75�]3�O7*s]��Q��4g T�`{�:`oH��]/����?{�1|�q�r5&h���;=�`}�U����-^�f-շ4�IJ��v�e06)��Ҳ_}��#W]�ηs@3��V��(DclRE������ၲ~t�ޑ�ܺ[ �0���G2"78hw]��ٙ��� ����=뒚�g4���	 �z�㜙,�+Ս�v^�p㱞ݸqm@����q��9����d��s4�mX����b�6!.0�3mX�w7�Cs��}V��)�ww-X�e��J!��V�˪Ժ&���Z}�O�����n��v��򞱣�e9t�T�a�$�fo���j��Nc��I�%d"�K�30���h��,b��F�h�f���Z�5(�ku�����{���߿pP�Rnuv��[:�*�)�V�v�ux͝U����6�y�b-M���;%��8Ye0=���+ �����}�	?~t�3�3有(DclRE�{nJh��V{�j���X_�L��G�5SI�*����R��?�����:`ṽd�M��wp���nf�ح��)���~%d�0:���BӪ��ʚV;�����W� �fڰ;���g�ݭA<�I$�$�d�G   $ �` l 	5׎����|����l�ck`�|v�z9�wa���y2:��v�v��)�"[�=p���;v3��Q��u3n���N١z4.ݞH�&qq��L��^3v��v^��2nR�Ӷ��vg���lv'ppӰ�������f���Ú��ss��vǧ]Ԅ��;h�M�9�ꜷ>�WQ����]x3�jB��]��=t#�6m���ms�bώ��9kv�J�q5 Ӈ�w�d��=u��� ��>4���#�"#`��@��:`wH���Y�(�E��#xH4I3@�s@󬦁�)�{�w4�r�c�?���h}������,�ܵa�BI'���`�_��ND�&!�7!�{nJh�o�g�[�ۚ�e4z��M(H�I����G{J)�Y܌5oX�s��s�&yA{l�G!r9�L�/�qㆁ�u��;��V;���wUi`c��t*��%��e�ѹ'���������j!/�0�r�����,�ܵ~�l�eW�<�ۘ��hߧƁ�)f�Q����w޵`quJ�9��3-,�Z���VA�����GL?~^߷�@��B>Cc�8h�GL�0=� ��+ �&�p��c,^����\޻;��t!���t���<#\��i�9ݘ�S~�/ϝ�q�3C�d�w���Θ�`N��`ott��F�6�uPL�f�����az�f����~��/[��s�+ND�&!�9�,�*�����VL+!���N�s��nh�>4�'�L�/�q<p�7�:`t���2������H@FI�73@�n��g������>4{��s�v���N&�[��χZ��l�Ϟ[8!�b{Q��$�6�;,��&$�M̍9��e4�V��Z����V���.�%e��+X0:J�07�:`t���+�l�uN��S�L�3MMs6��GLt�0:J�0�E�.
���U��+/$�}�|��Ł��XXq%�	@�B��Q
�Y+��\�mH�&��UM+�ea`yyF�˞>߿�4�w4)���iBE�&����ё{ u�zwn��X�c��-XN�'�&sS���"J���=�%4}���#��dZ�̬Yiʚ,��Z�Pٙ�j���ZXf)M�b�Ĥ	 #$�ۙ�w[��s�,��wUi`w���b��"B�U	�Ңf���O���`wuV��u��;���<�q婩&�M�4�`}��a%�������}���A}�V�H|C��Cj�=я
����%�P�R�I%5"�1��1X�F����`(2�@��-|�p?(ePY�[l4s:��    @    �   �   �         hH         �   $(     l     m[     H    �m�Mm�"t6�N�/k����)�V�{m�.�3���[��\͹�\��z���X( �:v���Ňm"�G�����q��R^��p�Uҗ,��UUW����dx�}��[Wl�nz�8��[��oh�V�rT\.4�����\@@U]�{���u��a:ܱrv@NE���su-m��=���Wq�mhY��ض�'d8l��W�6�뙀9�y�Զp�d2��N�ܽ���#e�u����Y�jkcr�pAG6��lqI�dx��r5jD^���k1ʰ7dBc����ܵ˸�iL9� 8[o9�z�7lPV��^��$�0�F=gD�q�p����nԣ���`���50�Sͭ��q;)K�l�xLbh���qڳ�uG.OnݷQ��q�<�ZgK��m�ݶ.�F����.�N8�2�������מN�ݓu�to�>�/6���Ocmzݪ�!�n���f��mȽh�6��\�h�K�NF"�QnCGV���mu8�K�v��!�c���I\n��dD���6�I*[;I[Q��tɲg��0Q�h����%L�q�c�ն#zrFݔP�s��J�n�*�JHs���O�&�{v�p��E�%['^)΍wm��e�`Y]%	�V��ͣO+�v����
%@�wO5�Zx6�g<�m�������s��[��$�nx灁�ִ�,��綷PX,`�aq�7[dq=�0�V�lr�k������dL�r6n�� ;�F)��V�lh�cV%��B�3���o*Z�u���L��Ut�W�"��IN:��E��V�K�T겴�@
� z>��QVx����R�� T4���>>��zjڠ�H�  $m��m�  ��!�:V���ٵ���Ojl��m�
c�o.W댳Kٷ=qE�.�2�ݨ;Z�&x����e��]DdCu�p���L��\�ny1�kv�O����K���Ħ�\�زq���[�4ݍr�n$6��
[;k��q��㴽n+v{V��uҐ$e�b��6�#������-��ˣ,V�/L[��<�`��y29ʺIe�6��U�r܏Tͼ��q�X�:?�oϲ:`wH��Ʉ��(�E��"a �Rf��n��S@��c�>��j�zd���Mĺ�PL�u4�����Ʉ��GL�0
��L�5M�)2fI��a�Q����;����:`{���6H�#3+���,�0;�t��)-��VC����v��0Qda+���\��'v�v�mt��ZV+s·�y�e3����V�@FI�73�-����v��rS@����*8]pɎnc��{���`�Ȑ
D����0�(�)��� A�
%X A A�1�,H@��H 0$�@#�`� �	�c !�@�H#B� ��E�W�4��t���xd�~t���k�WKK0.�X% ۋ@�ܔ�=�w4��}������=��:�e�C���8h���t���K`l����E�Yxd���.�X�e�c2�_ ��i`}m��/5�N'2E�E1�I��f�z��h<�X�#�"8���wꈦ��P�	�U3J��g1�̬,5&B����<�bX�'�w�6��bX�%>=�4��m�I�2MU;��!2!wv�6��� �DȖ'{���"X�%��߿p�r%�bX��]��r%�b2��52UR�(C�s4\.�	�X�}���r%�bX�w���K��@�>1G��`�H(E�G`�=)�MD��iȖ%�b{߷ٴ�Kı>ϻnv��I�,5�e�ND�,��"w���ND�,K�����9ı,O���m9ılO��xm9ı,N�>�t�&ֲ��3.h�r%�bX��]��r%�bX�w���r%�bX�}���r%�bX�w���KĤ/$�#��o�]:�Le9t�tITP���s`��\��"�z��S�Φ�R�k�j��0����h�j\�^'�,K�����6��bX�'�w�6��bX�'��xlD�,K�뽻ND�,K��]��鬺�2��ӑ,K�����Ӑ��r&D�;���ND�,K�����9ı,O���m9�,K�{�\��j��ɬ�\֍�"X�%��{�ND�,K�뽻ND�,K��}�ND�,K��ND�,K��y�-fi�feֳ4m9İK�뽻ND�,K��}�ND�,K��ND�,��3q5���iȖ%!2_,�4��m�1�2MU;��!X�'���6��bX�'�w�6��bX�'��xm9ı,O{���9�7������}������(b(F�	׆�^�ZJ�\�.7%���(��h�֧p7�ώ���L�T�i����!2!n��W�,K�����"X�%��u�ݧ"X�%��{�ͧ"X�%��}gs�]PUP�U"\Ҹ\!2!2n���ı,O{���9ı,O���m9ı,O~�xm9ı,N��_�ESjf�˚W�&Bd&B�V�\�bX�'���6��bX�'�w�6��bX�'��xm9ı,OO��T6�ʩ�Nfi�.�	�&B���ӑ,K�����ӑ,K�����"X�%����nӑ,K����i,:k.������r%�bX�����r%�bX�w���Kı=�]��r%�bX�w]��r%�bX�[������{��߻��޼ 	 �-� �	 �bY@ .��-�<���9�.z;l7!،�gsv�-]�q���k��*��ŋ�����(	uq�y9=�::N�.�eK4�D�]S����&3�v���Ѫ ݲ�;+ �����ū�n��e�n�3!	��s�Z�%�m��dx9�gQT�ݺ��l�<��G��;[.��Qp�k���c��`�_��Dn�9l˞\�fL�ˣF=`�D���v�zw..��/aʝ9�u���g��t�Y�eӓ5�=���7���{������Kı=�]��r%�bX�w���O"dK����p�r%�bX�{���n	�*	�U3W�&Bd&B�W{v��!bX�'���6��bX�'�w�6��bX�'��y��Kı�ݓQ3ASLd̓UN�p��L��>�wٴ�Kı=����K,ZB�ݨV(A	w'u�B!wfKO2ܬ�.i7�W�=����Kı>�{ͧ"X�%����nӑ,K�
L������9ı,O��?g�Z�ZԵ֌�4m9ı,O���iȖ%�b}��۴�Kı>�۴�Kı=�{�iȖ%�byӲv�2�V4$8�m�F��`]�I��p��!��wL��Wb�Azl���5'-�7�w��ŉb{��۴�Kı>�۴�Kı=����Kı>���ӑ,C{����޻��J%s0�|�~oq�X�'��{v��� �uC�D6�'"X��<��Kı>����Kı>�]��r%�bX�>��%�Me�a�T���ND�,K���6��bX�'�w�6��bX�'�k��ND�,K��}�ND�,K�{��5�k2k&Y�Ѵ�Kı>����Kı>����r%�bX��]��r%�bX�����Kı;�����L�4�e��h�r%�bX�}��m9ı,O{���9ı,O{���r%�bX�}���r%�bX��>�w��[�\Y�d���ڥ�����Ź�}����x���׋j�\M�g=�9��\.�-��2�k=���ı,N�k���9ı,O~�xm9ı,O��xm9ı,O~��6��d&Bd&��7e�3Jd�i��p�%�bX�����r�r&D�;�߸m9ı,O���ND�,K�뽻WL��L���ou˪
���-�+��,K�����ӑ,K��߻�iȖ;�)$H��ǸcJ�DR��ұ�$"����XJ B���j�C"8`U\z�'��{��~ݧ"X�%�����"X�%�܇��D�����iI3J�p��L𔐳7�ND�,K�����9ı,O=�xm9İ?ȝ���ND�,K媼x�T�%�"j���p�Bd&Bd/{���9ı,O=�xm9ı,O��xm9ı,O}��6��bX�'������&r0�Y<�G�|��NG79�uǰ�R97=	�BX�<ܩ�n��kc3͔���ND�,K�{�ND�,K��ND�,K�~���'�2%!2z��p�Bd&Bd'վ�(�4�N�&�e��ND�,K��NC���,O���ND�,K�����9ı,O=�xm9ı,N���h��4�32��4m9ı,O}��6��bX�'��{v��bX�'���ND�,K��ND�,K�>�N�3Rk5e��&f��"X�%��u�ݧ"X�%��w�ӑ,K�����ӑ,K���.�g���"X�%�O{	��.f��V\չ���Kı<����r%�bX�}���r%�bX�{�xm9ı,O{���9ı,C���~���!"׫i�w&Kn˷Z �G�m�W=�pq�S#��v^�����֌��6��bX�'�w�6��bX�'���ND�,K�{�͇�D�D�!2s}�p�Bd&Bd/I����a�k.L�ff��"X�%��w�Ӑ�ș�����6��bX�'�w��"X�%����"X�%��񮝲�d� sELҸ\!2!2{���Ȗ%�by����r%�bX�����r%�bX�{�xm9ı,O��]�f�&�J�U5E��	��	���^�"X�%����"X�%��w�ӑ,K����iȖ%�b_���4�ML�$�����!2!w��V��bX�������%�bX�}��ӑ,K��߷ٴ�Kı=>��~6��sm�m @	  ��� j����986y�d�d� �&�n�h�o>B�S:��[�8z�ْ9��OV��ch{"��[v��xro#d=���=������ׯ��αlwL�i]��у6�,r�Kd�.5�#:��tq�xmק��t� ��nNM�������v��g=�����%�!�ܓ�������_���6WZczz�뱕����ny�A:k͜�&7/>�E��Cۍ��ײ�7~{���oq�������"X�%���fӑ,K��߷ٴ�Kı=����KıMj͓Q3ASLd̄�+��!2�{�ͧ!�9"X�����ND�,K߿~��Kı<����r%��L���7f�MU)�p9����p��V%��o�iȖ%�by�{�iȖ%�by����Kı=���m9�d&B��ouӪ)��K���p��V*؞{���r%�bX�{�xm9ı,O}�}�ND�,K�~�fӑ,K��Oe�I�0ֵ�&i��6��bX�'���ND�,K�~�fӑ,K��߷ٴ�Kı<����K7���ߧ�hr0�^�͒�8���:�
gZ3tE���t%�X�Gp��{��q��n]Sl��9�nf���	��	��ܽ�ND�,K�~�fӑ,K�����ӑ,K��߻�iȖ%�bt=+Z�ɩ��UMQp�Bd&Bd/���i�P@ꫠ��Sn�r%��y�ND�,K߻�ND�,K�~�fӑQ�,K�}ܸw0х�d�L�����Kı<����Kı<����r%�bX����6��bX�B�2��\!2!2�[�&H
�f�k4m9ĳ�L��{��iȖ%�b}�w�m9ı,O>�}�ND�,K�{�ND�,K�;ܝ�0љ��d�Ѵ�Kı=���m9ı,O>�}�ND�,K�{�ND�	����+��!2!wsN9�-�T�qqun��xsa7k=�h�L��S��l��85�&�Ͻ���:>Ѻ��$��>�Ȗ%�by����r%�bX�{���r%�bX�}��6��bX�'���ͫ�&Bd&Bܬ�\�N�$UJfj�ND�,K�{�ND�,KϾ�fӑ,K��߷ٴ�Kı<���m9�,K�=��&��Z�f��h�r%�bX�}��6��bX�'���ͧ"X�tP��wܦ5
��e�a��C��xF�$D�p�����b6H�U���
E7E�H!	$I 0�A�U�y�1HDd!P�5MIh� @ �CHU	X�Y.��j˄Q`E�]h�K��j�ZLC@K�M\�L�s%���Ċ$�Tj�ȁb@h!4b,@9C�K)��{̄31"ā�tY5�A�s	���EH���R'X�� ��+�D4>�#D��M�*>�*��ȟDϷ�&ӑ,K����iȖ%�bxzk�n]j�34��[���r%�bX����6��bX�'�}�ͧ"X�%����"X���2��\!2!2��Z��UL�Xk5���Kı<���m9ı,O=�xm9ı,O>�}�ND�,K���p�Bd&Bd'�cѺ�4ɚuuv֋���͎-��!�W �w#I���Q���2&&ri4�|�~oq���<����Kı<���m9ı,O}�}�ND�,KϾ��"X�%!ne�Ba���&Fꦕ��	��	���ٴ�? �ș������r%�bX����m9ı,O=�xm9�L��MjݓBf��19�T\.��%��o�iȖ%�by����Kı<����Kı<���m9�L��Mwn��3Jd�sU3E��	ı,O>��6��bX�'���6��bX�'�}�ͧ"X�@G��U6B���\!2!2�X\���R�f�k34m9ı,O=�xm9ı,O>�}�ND�,K�~�fӑ,K����iȖ%�bt�����]LK��z�s�ַ=�p�Ņ�՝1�Mm"�p�6��dwq�WGg����������bX�}��6��bX�'���ͧ"X�%���w�ӑ,K�����ӑ,K����N��j[34��[���r%�bX����6��bX�'�}�ND�,K�{�ND�,KϾ�fӑ,S!2��Z��ULөUUE��	�X�'�}�ND�,K�{�ND��$.�ߋ��!2!fm��\!2!2�f˖=��mԲ�JuJ�p�bX����"X�%���o�iȖ%�b{����r%�bX�}�xm9�L��[�nP�m *	����p�AbX�'�}�ͧ"X�%��D#�����%�bX����m9ı,O=�xm9ı,Lv@!,�B{��������~�y�p� H ��7m�   u�%7^u'���Pw:v��N�;���λ�w!��Y뚞Wv9$�ĩ�I.�}dt���V݈�tyձ/"z-q��nq��h\j;��/l�CU��fIu÷i;vyq��&�`�n�n5�z�� ���v�l�"��lWh�N����785�f�:�˚�s^�1����ӛ��w���������H�6�Wt.���	g�֊�J��;<������{���;��-�4��XMQp���L��[�z\.��%���w�ӑ,K������� �"dK������Kı)�a=�&iL�j�h�\!2!2ٛŴ�Kı<����Kı<���m9ı,O}�}�NDı,N���fiӪR2�T�Ҹ\!2!2��xm9ı,O>�}�ND�,K�~�fӑ,K����iȖ%�bw�uSD��s*jM+��!2!}��ͧ"X�%���o�iȖ%�by����r%�bX�}�xm9ı,OMt��f��3Nfk.kSiȖ%�by����r%�bX�}��6��bX�'�}�ND�,KϾ�fӑ,KǏ���~�b��u���!�=���(9�L���扻���׶�fN���g:�WZ���r%�bX�}��6��bX�'�}�ND�,KϾ�f��$"dK������Kı=;�w)��[u,����p�Bd&Bd/�7��r1"!=Ν��K_�o�iȖ%�b{����r%�bX�}��6���L��]Ŗ�6���TҸ\!X�%���o�iȖ%�by����r%�%�by����r%�bX�}�xm8Bd&Bd&�nɡ3Jf�ə	�."X�%���o�iȖ%�by����r%�bX�}�xm9ı,O>�}�N�	��	����&iL�e��p�ı,O>��6��bX��)�{��i�Kı=�w�m9ı,O>���\!2!2ݠ�cuN�sN]P���\�l��z��<kk�giH��Z�u.��ı��X,�Es�]+w�w���oq�y����Kı<���m9ı,O>�}���"dK�����iȖ%�b}����e&��at�f��"X�%���o�i�~��2%��{��iȖ%�b{����Kı<����r%�bX���ۚ�Kff���\֦ӑ,K���ٴ�Kı<����r%�� x�Q5_}�ND�,K��}��&Bd&BԺ�Z��S�u5N��r%�bX�}�xm9ı,O>��6��bX�'�}�ͧ"X�%���o��p��L��_,�r��je�Rʙ)�ND�,KϾ��"X�%���o�iȖ%�by����r%�bX�}�x�L��L��ǜ��6*��Ӥ�u�J�)�*�=%�D��X{W"m���ftQ'��[�Ȥ��U *	�����.��	��?~���r%�bX�}��6��bX�'�}�ND�,KϾ��"X�%�V��4&iL��a5E��	��	�����m9ı,O>��6��bX�'�}�ND�,KϾ�fӑ,Kī�#vF��&J2�h�\!2!2��}�ND�,KϾ��"X�%��o�iȖ%�by����r%�bX����3SN�&*�u4�L���B����ӑ,K������r%�bX�}��6��bX^��|> ��"gw���Kı;��~�j�55u�]75���Kı=���iȖ%�by����r%�bX�{��m9�2!}���L��L��V7�]:�F4$:]z�x�l{q׊K[��[�N;:�
��1�Y�s��̓5��o����7���'�}�ͧ"X�%���fӑ,K��=�����&D�,O���m9Ĥ&BԱW���uN�S�.L��X�{���r%�bX�g�w6��bX�'���m9ı,O;��6���B_,ѡ�s,l&j�(X���A$Ny��M�?(��Ow�ӑ,K������Kı=��vPѴ����Ӛ��\!2!2���ӑ,K��o�iȖ%�by����Kı>�~�m9ı,Jt��hLҙ*�	��\!2!2ۗ��Ȗ%�by����Kı>�~�m9ı,O=���r%�bX��#�B0�eB�H�e��� !X�$�N��Ym�kZА�H� �� lK(l� 	8�vt�{H�g�E��'6�2K&��@O5{Q���km���9ɋ�����]�ug���(7�v&�U̱+�s�ŭ�����=��nQ=m��n�6�q�l��[��۬.�e�GL0����M����`,��i#nCd�r���o]B�k0q1��"�L&�2䄸�Ji�cn�~wts�� ������::�{6Vb�㋜C�B��l���k[��;��ݩ���u������oq���<����r%�bX�g�w6��bX�'���ND�,K���ͧ"X�%��e`5���*�LS53J�p��L��}����r%�bX�{�xm9ı,O;��6��bX�'���ND�9S$&B�0~򦉢�t����\!2������Kı<����r%��"{�w�m9ı,N����ND�L��_,U�fjhl��I��3J�p�ĳ�#"{���6��bX�'�w�ӑ,K��=����Kı<���ڸBd&Bd,K����U*T��:���Kı<�_v�9ı,O�߻�ND�,K�~��"X�%��~�f����{��7���[���2�뙌���<�l!�oE	�c/aʖ�xu���g�QВ��Y.�*dS�\!2!2OssiȖ%�by����Kı<����r%�bX�{��v��bX�'�m�6m �"dt�nL��L��sxm9 ���Ȝ�b{��ٴ�Kı=�]��r%�bX�g�w6�!2!2Z�dЙ�2Rd̄�+�Ȗ%�by߷ٴ�Kı<�]��r%�bX�g�w6��bX�'���N�	��	�Dn�R�M%�u4\�bX�'���ݧ"X�%��{�siȖ%�by����Kı<���ڸBd&Bd-��jvf���)�3UT�D�,K����ӑ,K��߻�iȖ%�by߷ٴ�Kı<�_v����7���{�߽���HZ�(|�s`��Ů7\�v�9I1ϐ�}�I��# OL�X�T�4Sn���U7�&Bd&B���[ND�,K���ͧ"X�%����iȖ%�b}����r%�bX��ٚ�*��sT�i\.�	����ٴ�Kı<�_v�9ı,O�߻�ND�,K�~��"~L��,��b�4?1UR�UN��\!2!1=�]�v��bX�'���ͧ"X��(aQ�H Da �@Ѹ���;��"X�%��{�ͧ"X�Bd/�m�h٢�˦�̄�;��ı>�~�m9ı,O=��6��bX�'��}�ND�,K�u�nӑ,��L��YnA��L�"�t�nN%�by����Kı<����r%�bX�{��v��bX�'���ͧ"R!2��=��9�L��4RU%���0�m�Anݗ�\����Έ�d�ܵ۶g9Z��ˣ2i��L�O"X�%������r%�bX�{��v��bX�'���ͧ"X�%��w�ӑ,Kħ���rkSD�@�UE��	��	���f���y�L�bw>���r%�bX����6��bX�'��}�ND�,K�k�);3SRU%3UT�L��L���ٸ9ı,O=��6��bX�'��}�ND�,K�u�nӑ,K��!��Q(�)�AI˪���!2!}��+��,K��o�iȖ%�by���r%�`pWQ>߿w6��bX�'�����Y�j��w�w���oq��w��m9ı,?G߷��i�Kı;�w�m9ı,O=��6��bX�{��w���3����ܙ�x�F�O�p�`݀M1J�<�&M	b��r�5�p��q��.��u���Kı<�_v�9ı,O�߻�ND�,K�~��"X�)��ܽ.L��L��ͷ-4T�uu�,��]�"X�%��{�siȖ%�by����Kı<����r%�d&B����L��L��YnA�RS�̗W5��r%�bX�{�xm9ı,O;��6��bX�'���ݧ"X�%��{�siȖ%�bS����34fM72ɚ��r%�bX�w��m9ı,O=�ݻND�,K����ӑ,K��߷ٴ�Kı)�a;ܚ��fMIl�jm9ı,O=�{v��bX�'���ͧ"X�%��o�iȖ%�by߷ٴ�Kı6�Q�N���6��HE�"�H��!(��gOf$�N��D 	�_��8���0����4aV[n*����$AbVI�Ra�l�n�h2���]��"�yp����$(*�H0���BM�ZB�P�(�"F$b��
YYBc ��[bA�2��mYy͒ ]�ڻ܀!�b��Q]�"�ܫ
�!6�bDV#'6&9����hd�
�,��6+��A�vB����.�r�Ē�j0>k�>e��N�h'[i�t     -�            �         �$          �         �`    �     H    �h+m��tn�9� %��(N��緈N��W���s<���a:.���;��F�-bۧ�ݱ���Yt�; 8�L�t�@��:�p�Qv,rҰvY7�&:��s²�n�)u:р��
vb�d[�Y'<V����r�p]]�]��^���b�ɝ�Ds���K�6��:��ݻ>y�{mm��q�n[qĘ��bރ�G�˸�!����dz��v�n��y8tWf�	݊!Ee�쌴��5Ŕ�w9�,@g��g�{k��[bl�茙��W<�뮠춱9�v�Gv6��"hPh�x�[Gv�`�GdY��6�/gv�C��l�Ksujm��+�$mbAJ�fp�ݖ��:v�5KP[۷���gU�����1���ʳd;f-.���k�XM�]��M�����y�\v�r����pm۶;1+Ŋ��ۨ�u�4k׎�>׭�駳�u�����&����гٝ�k���z\:�u(������կ;�/k$䷮o$�НN���[W�9õ�I������(�n�t�����S#�m�}>v`e�lER�i;,I�8/'vƶK�n-Խ�1fc'l�-�e{r�+�p�M�[�}�edu*ӹ�;�[�Z�\�7�\�-A.�6��W��8�T�+=�dJ
�H�[��E����G�] ��H�=<�κ��x:��vtg�;\b��]X�c��*q���!Q��Ff�y8Fn�r<Y#����h�Qͨ�g��A��ڶT���q�C�1ۮ����̀�\Y���h�tV7�rj�)�,�j9ƹi����r�P	�Vͳ��/R�4�svlhݩx����������������{���=@��#��x��|w����w��]���~d�my���� 0H��� .��$��0OF�e�U����&�^n��sp��^�8��[Y�uu;o�]��q�����ά{[�]��ǩ�ha��<uջN�VsrF�\ �|��r�P{FL��g5������rSv�vS^#�;�9&^�n���v��1`��ͩ��V������F��5�0���������|���R������v[��8�{v�b][��n;=�UZ.Ǯv�3�̳:�o-1����q�������ͧ"X�%��o�iȖ%�by߷ٴ�Kı<�]��r%�bX���Q4SmR���M��	��	��߷ٴ�Kı<����r%�bX�{���9ı,O�߻�ND�,K�n�5T6UQ$�S���p��L��_w��m9ı,O=�{v��bX�'���ͧ"X�%��o�iȖ%�b}U�vFU*D�Tꋅ�!2!}�۴�Kı>�~�m9ı,O}�}�ND�,K���ͧ"X�%��ͷ-iԹt�\���p�Bd&Bd/�߻�ND�,K�~�fӑ,K��o�iȖ%�by�۴�Kı?���{���~��1�.��}����^���c�m�5��z�*��hW�ؘ�W]C�f�"�t�y�!2!fm��\!1,K���ͧ"X�%���n��șı;�w�m9ı,J~>�'�f�d�ə	�.L��L�����r4���"�46�'"X�k\��r%�bX��w6��bX�����p�Bd&Bd&��3eԧR�f-��M�"X�%���nӑ,K��=����Kı=���m9ıL����p�Bd&Bd-��jvj��Tj�3Z�]�"X�%��{�siȖ%�b{����r%�bX�w��m9İ? �L������9ı,O����M�*��U7�&Bd&B�r��\�bX�'��}�ND�,K�u�ݧ"X�%��{�siȖ%�bw=����K#	u��6g]k��OZ������s�.:�)�މMt�ө6�5틉��Kı<����r%�bX�����9ı,O�߻�ND�,K�{�˅�!2!duV�9�T�GSTꍧ"X�%���nӑ,K��>����Kı=����r%�bX�w���r%�bX�ww)/uu�.���&f�ӑ,K��>����Kı=����r%�����"j'��o��r%�bX�{�߮ӑ,K����ܖ�3FMXL�uu�fӑ,K? @Ȟ��?M�"X�%�����6��bX�'���ݧ"X�����fӑ,K!2Z��x&�%C�j]Qp�Bd&%��{�ͧ"X�%�����iȖ%�b}�}��r%�bX�}��v��bY�7��߿��aPBE�k�pj�SÜ�i�vӧnҞ�x�gT3\v�]�ڒx�F̘��7�x~ċ���
���W�h[)�{ρc�G L��qh}�M�DBI6}����kK���r��P$"KLN8�9�Z��i����{]�h[��=��hܐH�5��9���M�}V��^�1��Uןo���8�gԗ>�uthn���,v{���J";;�<��`w�S@=�*%"q�?E�`BF)�vF8-��Nڱ\�Ru�geu�;;s��!�����F�ĕ��J���`m쉁�[vd����1*��D`آr=����0;WK`m쉀WV�@Y�$eX��y�vd�K`m�@����g�ëQ�#fLM��Il��06vA���[yp]*�q�rI���נ{zS@���h�h��դPo$�I2I$��H � t� � I�ڻ\<Úݾ��-nv�1';��G�s;�V�Ŵ��1�uK�0�xmmYYӻ���\Y�8�\�GH�L)��te�fR�u�r�nM�� A�ܙn��)����̎��6�k��T�:ۋژn�`F�x��mV�E��W��v�N���y�X�I��Ҕ�ؖp�����w����w\�|�ed�0�[a�c�����T:L��a�s���D9q�k��n*�L$"M�15#��Қ���@�]�@�{k�<ˎ�n8$I��y�07WK`v�-���gd��S�vGN�&骙�`ggu���06vA���[�;���bB�WV�-���gd����w��-���/��Ȱx�nG�{zA���[�Il^Ș�A��Wv��H�q��㮅ݝ���6�AM���6=�+:�::9s�n95�\.�)�[������;T���쉁���[
:+�N�Tȩ9��v~��|P�kQ
�D�A����]���HŜZ���0  <-B1HE$Q�bE��Sl�4�bDш��H�EEH5�$ !�Q������	����@�I�|�QdW��G��/|�7$���h����|r8���I"�8�̛��Z�TD7��k�3����V�@����bjG�{��h����v���@�.;F�QL"j�Sut�����07�t��7��%b�$��e^�7e:�:����!�����RD�˻#�d�����W:\+�`o)-������;/F�%G#M`�Z�۹�{�:`n����R[mvZ��%���%��)��#���l��}�V/��R�B��DP=E����rO�̵`|�,f�'2T9���+������)���0=$t�+aD���lɍG�����m��<��h������JD�DԂ���u�����{�n���ZXj��t]��3��[��Yfa�|�b�`{dt����uv=�ID%������vi�U�e:L��`s3-^-J%2fN�d���3�}�rA(�5I�����������Vۻj��|�X�$QL�(dn-��Z�۹�ym����Aֽ����I���̥�L�e�Z�K-����GL���Ϫ�*)���FH���!���=�-�s��S��a�M��ra��d�����\#�%�ȱ�������ۚ���@��M�#���K ,ʴ��Һ������;� �����#�[
$�����ife�;� �����#���lj�Q,X��,�,������GLj�l�����E��B&�)��f��s@���hϪ�<��恿�{�NI&I$�$�8�  $m��`6�  �$���IúL9� �v:�`�i1�,�.^pFR�-���4�S
��8��c����>V��)�˲hN�v�S��qY�u���r��v�r)�v�k�c�'�.6�N ��&��kH�7b�d�̱��{HsB;\^��;��v\�.�\�g�u�6f�$�v�����+$IБ��\�Y8��/�񨞷:�*�v�^n������3G\ئ�E��
L������z�h[w4��:�N�E2`���;�K`{z:`zH��]-�*��_�%uw�/%�� �`oOΘ�:`{WE�w>���tO��2&$�Q��7dt������]10=�06�jYA�&��6�73@���h���=빠w��h�n�%"q��IF�q�n��04-��8���8�s�F{\��֧p5Ѹ�x�HѓrE�w;c�<����#��t��p](�,Fa�|�fkY�'<�훠�ر
�
��Qid��KR�"H�P������}�U�Wn�fx`w.���t���vU\P$"m☈�h^��<��Z��z����r�QH�%"�yW��ں[E����Ӳ��:�N�E2`���-}c�>I(��zp�+K�Oq��>�F��&\�]s3�l�k�vϘ��vͻn�і�^��<u#s����T�b9bӶl��7�~��`{WK`H�b`v�D�T�(%ME$4/Jhz��2{�6>�az�%��V�Q5Iԕe����������T�J">HB�]��p�<Q���	�4�8� �V,H14R@��y��JLb咙���h��$��� a��a <��Z@�&(����6(x�A}s�F�'�����> xh�0 <��(��g��nIϽ��`�0�x�HѓrE�Z�Ǡ{{ ���ں[y@�Q,X��,�,��Lod��`{WK`H�Ǡ�4���	D�@��~���jp�:૶9G�����$غ��1=2��E�6�LD��<�)�y��_X�=�M �.u�bQB&)�Hhz�[E����Ӳ�iK���QH��@���@�޻���Z���@��F�%b��$�)#�=��`z.������~�W�}_"dx��tOH�x�I5��<���>��z_��}�G�y�Jh���%"q
M�6���u�^�^�e���tr�=�B�:ı���Lv��V�Mv���Q���_��͉LLod���
�B�^e+��b���S�3;YN��&ϻ�����|�=}V��:n8����$Z��E�����tx0=}R)$�2$�$4+�=}V�o]���)��΢q�j(F�LnK`{WK`I#�����Il�z����B�(BP%bB}����� 	 �-� �	 �bY@ .��-��ή�iZZ�ν��t%�[�\�9�D���N�Y��y{a��_�݇��l@"��S�������s�g;��-��#k�������D�gF��'U>``u�5��.C�H���p����ֽ������]�D祧Y[�h��2r��<���N���4��zq��t@lv�w{���{����L�a.�w&uɊ�F��kv��ǃ�u��.Ύg�3�ʜ���p7�،ˀ{�~x0=�0=��������F�%b��$�Fh{�s@�V�篪�:۬�;��
�䘖]ڼ�YLE%�=���:H������=Y�T\#ɑ��m'$Z���@�#C�����l!r�*�V!%����#C�����z���D���	���%1LdBn�]�^ ^ݠ�V��r��s�qT��u�ݗ�`v9�8���D�4=�M��Z������3wnK�n�UR*A��5SrN}�}w�I"A!�F !ZJ"#�"���X��̹,}ܵz�bAs�
G1F�#�1���;��:H����t��R[��R��J�Ř���v�����͵`s'1�z���X��)I��=�0=�������#C �:�1�.��)�G\/9��<6�v�tW9�:k�������3��vf��H���K`{WK`t���}�������uk5*�IP�[��v>��I6f�ܖ�͵`s'1ިJ�4z���U�&f�����rX��jʈHHJ!%��!DDU<��`}��;���%�ԓT�sM�Ia�(P����V�;�����v�By������[�UT����ʱfE%�=���:H������6!nm�&f��.i˥H�R�Z��\�zn���KZ��s�v�(lR;����H�(�xLrC�=�~Z[u���-lq��;����hs�]MR���vs2�Q�6}��V۵��ϧ����mbn�c�A������=&A��]-��F�mvZ�Ե�*҉�$s4-��<��Z[+Z�� �dBBD$�	�@XI �	 !��3߼7$��"�L���i7!�y���V�=빠yl���u58�P�(���]slus���'v�p��uE{r'�y�·����헤�1L�$����"�:�Z�=�0=&A��]-���Z"��E�V��1[����d���$�h,������nf�岚�t�Iގ�J�bYW��X��Y�0=���:H����t��$�nޖGT�MΦ�U)j�4��D�ގ�� ��������-�0 �8h `��M� m�8Od�W��{m:��!�	"u�,k%��=�re�u5�a,<�F��d���K��۱�L��r���Y�Z�^k:���]q��l:m���ڪ�����٭�"v!��j����Y����PQn�2�����6�ɹ��ju7R��@"%�A�;p!�Ӝn�3Tu%��մݱ�V�>�����`���{Z�kf��\�J�t��U�cv�M�ˢ#���ʜG4Z�d�/�?:`zL�ں[��&{��q�IDҒ9���hz�[��&����mK%�+�bJ�����$h`{z:`zL��g�����Hے-�Jց������t��(���/2ϭe��loGLN�0=���:t�h��T6�Pi���,�F&sOsùP㋝՚�]�2[Hͱ�g�f�n*��т���nf���M�_U�u�Z������=���w�~i��(�xLrCd��=���Ia 6��>�k�oGLN�0;�.��%y���X%�����=�3��W�{�gၱO��sލ�J�<PƟ�8ց�u��<���<��hzV��:6	��%J8�hW�hs���z��s@��MN&�fH��b� a&����Ә�6�I�v���v=�%$t<����i���iɑ��NH�9�Z^�������Xw�� e�}�C� dcnH���x��Lr����.��ޥc��
�qI�<��Zw�?�(������'�W�uU7�Y-�5H��].�^*1��bi��<���<��hzV�>���~�4���N71F���cr-�WK`t]`{�:`z.����]�WC�	9�YW�GF#v��Hs��T�;sӰ]rM����2{q{l錕7%��E�&�����lj�l	[ؕ�VF�����Hց�w4+�=}V�ץk@�s�`�R9�Q���+�=�`s��;5$�nV˰>��V,�*.��Ɉm�$Z����O��I�}�f�;$�R�X��U���v �a���%UP*�fj��;"������lr�l	w�E�M�ls�ؔ�,��]V�r��MI��\��i���ű��k�a�[����t��t�ް��~V�՗侉@��a14�hW�hs��+Z��s@=�թ��Pqᔖe�=˥�:vElwGLE����ƝcR8�O �Z^����-X��;��ef�Wr�Zoe����#Z��s@�@�U�{���.��
g�$��� A�X�;#G6�!CF2@�$$��	$d�Ri����+���"�b���+b�����h��p*���i���"RƐ$���b#�! �D��!���+��+�$����h{D�
UB�I# � ���˚R�T��jͮe�l�@     ��  H        m�        �[@         $   �m     ��             j��2�ۤj��V�ۃ�:¨v���mɗ�g�ӭ҈�L��NlY�/Y(�ʧdq����<u�*��	�� ���ݐW���ٝ\*�ؗmr���ά>,gV��%p�݂��x��ui5`��6ĺ*�S��^7YZf���K��c�ewK�
R^Jp���U�A��&�e�i̮�I����qs�^�{��n�< �-�(���=ttJ��hl���8��V-»�,�v�Z�nݑqkM��[��(��bt�Sj�76w+�:뛎ͧ!���\�D�.��̱]��nv6��5�Äݔ<n�,x��݇����'���ˊy=#	촁�iM<J�l�vK4�c_'�p�-�e@��eش�;صp�C���L�md��a�a�&~.�o��h;�*z�d�&xvt����m�Gh�J�ۘ���z�;���n7j������[���y�&�i4�ΌL�Ä�g���Z��(%���qS��i�m� ��R������C��/�*�l����hw�u�
=�F.n,ljڭ1��1Aɩ-��-�Gk+u=<� ����v��չ�nNn �:���\<�d���NL�ո]n0�D�K������]�����͛�4jƁ��I����UH�\�&f��+v��s�ثn�`�c$x�]����ܜX��۰R��Jt9��[��]��ݒ\�j��[\Z��6v�L�rD�����nr��i�*=�tl�:E�ZجK5�Ax�#����vH�Ӵ�.��D�X�(ڶ�{]�5 �*7Ku= �Z�v����*�������}M6��Hv��w����gW�G�%�M�t=b���z�ꮹ��jK�f���$ @�m��l m�]\&��wM�ݎ�w:��W��1�m��.ۑwZl^��m=��n� l����1�� �4�b�r\9#A���L��9�n�9�����eòn�wϝ?9��v�;lrK��ub/v����I��Ù,`D˭�inɚ�ڋc$�ڞ.Za��^y�6h�TM�L`j�����{��w�{��̏��������٥��L��ї�Y��/��`��g,�`���>Jbo'#�am(��]�hs��+Z����9g�Qp�$����̶�t�Nȭ�����^�g��wC�2~�m��ץk@��t��]-��]-��J�#3̫*�Z�V���t��]-��]-�ӥk@�gT�DdC	�nf��}V�篪�:��h{�s@뎥SQF�u��g�r�v����I�<�r)�����!L�3E̔�
Y-�Z>m�?���$�loGLE��[J]	K�Ey"�-�b���bG����<��v>��DD&�]ʙi��R��D���`oOΘ���=���$�l�:<x�N9�Q���f�yz��g���k%�lB�����1���*rb�ێI4=}V�ץk@�޻���4�D��8��N`�MO�ͺ��l󖃐���Od(Mx�n%뇭�	����-ć�d�ے-�Jց�w4��hz����A2�H)1�NF�oGLӦ0=���:vEo��U]��g�/��df9�nf�{��hz��8��0�t`�"�P�BXh1)dD +��9���I����nujF�&����������=�0=s�`um)t�D5$�$�
E�u�Z�<����^�篪�<��
��c���� �YL�Ƴg�� �����ѳ�R7<<<�B��F(���I�<����^�篪�:��h{��<v8�	FҒ,��tLj�l��[����=άXG���ڒG�y���+�����tL���U劳+>�$�2�D�ގ���0�u}�W��Ƅ|�G����w$��=���&�&#�Hށ�w4��������@����}���_&���D�Q(�<]:�LfC�']�����	���`�����1��9IH���b�����@���h_V�=빠��T��M�5by���]-��tI�������ubN��$Q'�R-��ށ�w4�1/W��{�����mbTD�+ϭf$���t��Ή��]-��tO@;�����0J6����<W��=���:.�0=�0Wt1]լ��� � v��m�,�m�6� $�J씼��n�sRM�{1���V���1^��`�g��x�"�4R�p�i�]x3�%;����L�v��f]Q�d��ox��+���ۻ]1������7��9"�L+��pa��;�^J9��2눊3z{d���iPvA���.v]�ݘ� a2�2�t%��2v���1��ͮⷎ�k��策?��wÕ�]ht��=k�nݳ1jn�2F,#ɊDcmI#����u}fl}ܵ�"q��sf�V:�2UUg؄�f[�������&��Z�� L��"��I#z���`z�D�����ؤI��]���W��R2�,���Lj�l�D�jJ"����Ǯ����tK����`{WK`lR$���t�������g#	u���Ʀ�v�ω��4>���hry�p�H�\ܩ�n�N��I�̶�"Ll����07WK`J���M�AR�]CST�}�j�(QȺ��Ͼ�������]-�����&�%O,�H��$s4]k�=��Z}��(o��u�wvՁ�]]�*U'T�2�/107WK`l�%�=�:`u�g��wC�2~�i����j�>Ȉ���\ń���vٔ�LӖ�!"ฺ��m@%��;@̻��cg���\�nv���ż�^��r�/�Ol��}"`n����JK`{�K��G�L��L�h�נ{��n;V���h�*�H�&��1'ut��R[6�>�>u��W�Ij�ց��^���:�n�rF�O�R-�K��=�:`u쉁��[T�J��VL$q��cqh{n��}���;��h�}V�{�U�8���&Y":�|Z�f�[,�����1��4��M7I�P,q�y$r@Dm)#��r�נ{���Oq�Qa�wmX5�6F��I�2�W������6R�ll��{+��8��y&Oэ9"�=����#�^Ș���=:���Db�r�j�UM;IDBO���X��6�>�B���>y%Z�򤬍�Fc2�,�^Ș���6R�ll�����������+%����Y�{����BE�����f�q�4����t�)��qm�P�iA�q�s�-ۏ��<��������ucn��"����E�{it��GL��07WK`J��]]�FQ��^}t�[�#�^Ș���=��� ��7��I�#iI��dL���)t��GL]utb�<��F&Ȥz���@���l��{"`z�Uw<�%�U�����,0�-���`��%� �8o�_;|��z��j�e�\s�����z%�нI�۫���r{9���;4�-Ց��ql��fӃ��j��ֹ�t]l$呪v�v����7C��b��+p��v��f�7X�ӫpV���w:�@��ۗ���+��k�=M0Ae�\u��=�g6nv���y��Kn�U@�-75����n��n�X�!:1���#����p���X�<�v�Uy1=�/Uv�U��W^��G�m����������ײ&��lN���Q�-Q�Y��e�;z:`u쉁�[eOqߔBM�5��Ne�)$�ۚV_~�����6R�lގ�ʗ-d�J@���@�@��������^��\ucn�RG��R-e.�����ײ&��l�����2��jѳ{�F%s���e����ۍ���kE�:���sJ닊d�r�����6�ܘ���=Է��v�7�,R8!6,�L�9{k՛�3?�����K`v�t�}vmԩ�F,���&Ȥz����=����빠r�נ�zu�i<�F5$�@�R�lގ�{"`z�D��ҁt�#Ȟa"���;޻�/mz��z�U�Zêq�4�jaF׎k�8ʝ&k�hj��z��k��np�n&��e"o2c1$�h���+���}V�����nU\o""�P'�L\�)t�oGL��06�:��q�8ؿG�{q�Z{�sO���!�]/�1b�XX1���RJ��q�&�`X�Xq@�X�>�	��H�	1!"B� E��r��)+b�@��!�#�D���^1(D�eZ	u���6H$H�Hf���y0�p0�,d7*C��A2��jh����y�g���! �P40�$Y		14\"X�%!1V�F�)�,LA6B!��b	! ��s7�1b�X)D� 1b "a�	��0b��H��X�a@#��u11]`�Ņ���#�$�h8D!��&���E�C�M�>���C��~_ i�!臀qT��n
� fv��z�
�W�\�@�∑I��X0;z:`u쉁�[e.��/��
゘1F,�L�9^�@�@돪�;޻�u��Q�$X�p���[k�N��9��v����Ƿ��d$v�r�r9���b��$q�W�h)t�oGL��0
�i�Wj�@�Ɯ�hq�Z{�s@�mz��Z����qǑ@�,R{���H����:R���P.e���ɉ'3@�mz��Z\v���_�H)���pyϧ��y�r���"(%~NG�y_U�w�;�w-Xy�6��t���F
 ���.���7cN�/#��*�'c<P9�'��uIG=tr3���? �S���ܵ`u�d���s]���@��Q(9����;޻�+k�<���:�h��`�p�(ř����&��l���oGLw��b��$��W�hqڴ������<�N��'�L�k3-�Ҕ������$LE���n��{�?��~�n �m @	  �l m��I�����wFmnI3���)�u��O�qM���ˮ���#�ӎx�4v���W���m�s�6x�2ki�;l��["Gf���$v�f���*�b.��Du�h�޳Q���/;�=����\b?��/�[��U�6�vN��v��{'.�6�I��ڙ�[�^������E�M���lJ4��u�I�p�MM��n��Af�a�%���P!��#��-�nh��@����Qa��u�d���P�I)6��H����:R���0�Z�yH��15$�<���-�j�;޻�m�@�.<�u����Y���������I&0=K`u{Ѵ��#JE?�Z{�s@-�hW�h�h֨өČ�52r���i��k�6�n�G���J�&I흖�?�s�`�m�RL�(ŒI� }��M̞�3�?D(��m���U9�3Z,���kZܓ�g�]ǚ�Q1~��*S�����I&0
�i�Wo$��9"�-�j�;޻�}�?$}��Mߝ�h�#X�ȞEH�8��0	$���l	)Ilr�
��
@c&$�� �٠y_U�[�ՠw�w4.>J���D�ME ���z7/Wg��^I�q��/"�nݮn+�AvL�3E�G$Ȱ�j��@�@��@�z�h��ܸ�i�'&�Y���������I&0=K`u{�4�)G?�Z{�s@-�3~�U_}�S{�`v��lo$�n�,PQ�$�4�f��}V�n<�a��(O;��`|�a�J*��2efff0=K`IJK`v�t�$�����߿1���'7�f����`w �Og��;�h��e��3��]y� �]��k3-�%)-���� �L`z.�����1<�0�dqh�]���A��}4W��[�ՠy�(+x)���s4�f��^�n;V�����n\�"�A�RM�ź��1���j���IG$���"9˝ڰ8�J�R�d&�������������I&0=s�`{���e�%� ��Ň8H�Ņ���R2�G���m�;\�\\.�B��N�7�,�`v�t�$�\�R�l�Ͱ��b�$� ���<W��-��h�]�՝�cȤ�Ɉm�$���z����}V�[�h�u��nUT�IuUSa�BOuVk`NS��	:c�:&�R�)YV�(�E�E�w���z��z��}V��g�ߗ���I�I$�$�m �	 �cv�   �M3v�U��5���A�x�;���ݎ�q�w]���в�nQ���:�>�Sx��s^\�l{�0h7B[
��x����ۤ����ȍ���\�N,��*�
TT�T���ٙ�*�y���=��q״�͔9�cxN&7e�*ۮ��Gk�Kf�gm�tՄ��:t~{�{�|��!jH��7';���u��\:r���{v�Z+���n��(s�@�V�dģ���女�^�n>�@�_U�\:�&E��P&(����z��[�t�'L`mJP�IJT�7~$�@�U�w���z��z��މ�L��	��9���߿+�����@�^�@�U��m�1��((őH�޳@�^�@�U�w���<첉H�Cj9��f)n���;,�=��x��_W:��,�6>�E���Ӟ��NLCnI$�W��[�)�w���z� �?r�ZO$d��Ԓ=�u���P"��@7�ﹿ���z��z�ێ�n���C9��t�'L`z�D��� ��%��:��JM�Ӱ򈄛�ͫ�����]��}V�yp��@���Rt�������(�Y�\;9�@-�4ԕ��q52b��5�����F�/u��w&�C���S�D棷9nc�q�$z�n��Қm�@�[^���F�X1BF��L�;� �$��"`IR:`z�f�kb�4�f�ⶽ<��� ���U����nh�JhW�����N<CnI$�8�2lřj��{XXjQ��ݫ �r�>y&!������;�S@-�h+k�-�n&�$J&��n�9���!���1Zc�pdA�l��v�;vo#���72bpP!�����Қm�@�[^�nYM�yAX��Hd�) �٠x��@�,���Қ�ë�dXH8𘢒h+"`IS ��� �L`uJP�I\x�n�I�nYM��4�f�ߋ�S��F&IW#�X4�R8#�� @
*V#PB# ��b��h4`HF@�sW���8}�-���P�9��p�;�S@-�h+k�-�)��UD�N!��F�&d�����������m��̝�ƹ&��3 Xv�t�#X��8��4����;�S@�Q���ƌm�$�fM�f��������33*�C`��_g�'�2bjI������;�S@-�h+k�=����D88�ĝQa���e�`��`q�d�j�Q4����%h=���(��Q`��`^�����[:P}�t�<� EW�� �����"��ʀ"�� ����"��� ���� ���(����# �"� *�"����"*�"����@@�"����"�@�"��",R(��"",��$`��V(�",�,Q",P ��B(�  ��T_��_�U(*�@U� ����"�� ���*�� ����"��*�*������)���ȁ����8(���0�?��(� T��Q@m�	T��  �E U  (�  �
      ��RQ��UAJ� �DUAT�PR�U JJ(I)JQ@� ��,   ��"�  @e� w�d��NCݜF�@/�@0	u��<��d}�Ft�[�9���  f�eu���e� �R�T�g��y�����@z�tU3w-c�����u�e�  �x� P �  �R�m����ܷ�G#y :&3�q�t�-ʹu��{ͳ|< ;��ns}������ ������oU��P}�[s���q�v����m� o{4�g�e<�F!���.�Q  P@@2� <�LO ��8�U��<8 g_mq��K���9זU�r�WÁA�E�����w��|��NC�� Oz1�,�=���G%� =}����ɮ����r� >8�     ,���=Ɯ�Lr�$�6
SM��9Ҕ�AJQ��
ce)JX��)� ܥ1��)L@�)c4���)Cq
:R���)JX�(�1���Ll�)N� �JR�h�)����ҔR�iJP΢ {4 ( 
 ��d �JS)JR�i��1R�ǁ��@����:�_3�� 0	|�d< ��L�^B���O]G�NM���w�@��N�1�i��g��pOHI�R��  ����i�  D��Rdԣ� ��T��D�  O�%M�R��   DPLRU=SH���t�����������$��sޏpo���"���o�DQ\��
��!EW�DQ_�QDU`� ���'�
���LVBHH0n2DD���S	����
8�*b�Qr����8��@�,i"7%kQN����8���f�c�hT��Q/V&	�r%�d�Lb�	@��L�J)L8p8"c��Cr�Ą�f�\�7�}�eq�D�ό�!���(e�āB��B%%��L.�M�J�Cl`��"`&�nP�$)��&u���2k8%� οg���J�Zi�V�<h۹6���Yqæ�u�A��Br�g������u�t&��c���@�&��q�A��Q�S���_�ĦL�ټ�@��W�$a"Q�!޺�x8i�I���pcl���Bg��!ɠ�I\g,3�+Ä�J���k�j�b͔)�
L�a����w':c��a�ı�BD��"�w
a���:S{����ʴ���\!�݌�R8��$��#V5e0B��g�(P�KX��\9��V�{�)�*��x�~$�P �L0���+� ��"�W2ky6��L\iٗ�ڄJ�Ν�]��F�:3�i�H�É2��`p9�ظ �f �:(�0���W)�40F���SOJ�t.E�`��1� ��Y.�a{��l XYR$(��(P8�Ԍ&��q`1��O�w��rlЋ! �!?),ptЄn���pȹ�tm� ���,0'3����ٽ�9������;d�q�t�0o��
��1��!!�|�4b�t8'���
0l����@�B�p��*@h����`2-�p$Dy/,]��D�آ�"BQ���Ȟ�Q�S8ɇ&D�`U8��L�ٓ*B�+��I���$���! )�2,)�����(�rf�hNnӲ|:�4$3�>X�d��E�H�Q	JR��ž�	J�_���h�My��>��M��׳H^�Ud6N�2���,*t�[��Rp���1I�b��K�;W-ɭ�b�����! �q�"��@�#�4�>
f�h0`�>��!ʖ.�#�MnnOD�����U/r�V<�O� 	&�@�!,,�d�*pFD�$J0�	X�
�R5�|����=����"�û��6\���#$�"C E�X�p�$�\1��.Mn��)��L1!���m�nt�FF��C&qI���+q�`�H�-z��L=8"�J0c$dv9\L����Ь�AO�%��ʳ5���zRn=Z5��R�͵)��3C�2�]L9�+3@���Zѐ��p�i�����٘P�k�"�*W��ZH�a��i��hd��&�8B�bX�c�R�kXS8ƸCP˳��0�ѽ������ȍ1�A��$�
r��l�`C������P�����$i��o&���[v)�ɠ��K�w�)�I�E�0)�cP�Y�T� �Ӕ@�1.R	L�cTd26�R��)[�!!$�(�,)R U!�f
��
�H!
�
	LHƸ#p`��f�Y��
�Kc��$ Q�+�WɆ�iZʄaJa\eZ�#R���������S*���#c p3�hшHS��!H�-����)���6c�w�89��{ڸW\���$i�� �ɤ�v��Z�M;xB�2h��Ӆ�� H|��������H)K�;0ё婨�����	�G�:Xf̤;T�'ʮ���B��-D���u!�����H��z���j�=^�H�!�xW�\e�E�E$��2_� ��׊U��o��ka4"��YY�~z�P��x<(�-N�h��0!F��bB�!XR4�*o��UjdP᩵wU<			ʡ�"�B+�`�"�`�xl��댘o�.4�ѿ�)��P�	�
�P�V��z�Q>ؕ���Ӫ������Ʈ��.1n1& XF�<'��ˁ	�1���')�bg\у{>��k�vl����X���J�+J��,bC������e�l�`@�!B"� p�2���̌�;
�&�Y2�b�T�	�4\ao.��H��A�]���M�5�� �"�1²A�Ij�C$!��"b�GM:$�3��>�Đ+�1�Xв��PE��R`�woL|1a��,��h`3�t���4����Q��� �|&�H�B��;�H 4rO��ʙ�ű ��I$�t �"h���u�`Ɔ��4S���M1
B�Bơ�P6e�Ӌ�滎��q��Ο$
c.���0K�P���|��&5���a�����h+��m�Ld����H0]ߐ��#Q�\��@M�9��q����\��&ο(dL1�8��S��Mk�Y-��'�V,2A�:��HA�@�rCN��C$i1�9bkg�J���@�r�)���3/TJ!#�[QǳU�V��B���}F��xMD��7�r��XyĨ�l�Ք�ìs�gL��2�N�!$E�{��H���zr��Ww�"j�M��#��
��=�n+���S���n��Y�Ą҉U���qԡ�<�y
/���0�.rl!q�5�8��.�5YKR�8��W�}���-&A�h��+n_��)T���*{�^#}P�0.�0�!��K��1�xo�$��Kn��9`sC
�˪��E �!	�]W�K�ٍ�v�c� #��/
)-���li��BP����D��%�W!�ԙ%�CL�68�q�[>8o#
�r4l��ǋ�)�.�a��H�e�;t|�>�1�F��8�:/�	�|�E��)�%H��������d��ܑ�#��>�0�!aL2����G��Rc&��ٲ1�!���N�t�8��Ai�F�G�N|I�dt�1���sP]�?3��MD��)NMmiLc�u�oYaXˌ��s��i y��L�ۗQ{wQg��+!D�>[�dHlHccB5�a_�$aB��O��t�v|m���!C]l>C�Ņ04l����b\];>>���&�l>2\4��1@�AQ�p# �d�Bi!(�)	�5�!��F�1�0��1�$aJ鋀�����F����$$����jE�	"F@���в+$J����0(aɌ���Ðd�p�JZ(T�X\��$"�X֚i�5ͅ22)�9	Z|��	�`AH�w�_��!��ʱ�rN/ <K���ńX�#p0٧ d#ާĒ2!8s4m �p�R	 �U���%~N��;���ˡ�#�>U}V��9Z�ߤCP�
a��jqyF�3�K�^���o�H�|}P�.c����6Ή$\p#S�C�c!M�i��0��-�a���k�W���|8��ݕQ�\����7�5{�e�W��P���2H�!!1�q��;��(�>���  m                           m�����                                  	��m� 6i�M�b�/�O���6� $Y���$/Ke �ų�H[��(:�5��m�)��&�MM��	$v@-+mi�����A�l$�f۳m�Re���2�o[�`�m������m�       [@ � E���m�hڶ�����f�j\�&#Wn���*��f�U@k�� �ͩʵUUJ�\3 � � �ہ[V� �����> l� H2l�mm�  8�i'L7[�ڱ�p[�6�`   d��j� �6�r�UJ�怨      �m�l�nkH [@� tݛl�m�   *�Z]���UIiIj��]. ͮ K(���v 4P                             �Jٲ�           ��  �rD�                                                         �|                                         �                                                           |8 �m�-��  ��                                                     ��    l�j�M� �+m�n�� R����-ҵM��i�l�ۀ$ lv�V�m�I,��h�o�I��(�R�l�wm�zvjR@iT
���  �8sm��H�`�5�M��h �m�n@v�d��� � p$۶� K(��z-� -���6Ŵ	$Y"�b��9��� 6�2���:�`�[j�a�a�ʩb�YYV�Rʀ]a\ ���l�K���[�T���Ԇ����e��  �6�l�\`�B��8ٺ�|���s�$�g��v���l 2  �-�L�-�x����z�oP	%��[j��VU`��HM�I��I�z�F�L��e�� M�      � $�H�f�v�6�&�Э<����r�ʫ�ͬ
WjjB@���;` �R�   	H�޵n�6��i����+�(�!H
f�!��mp��6��m�t�`   3�7@(R��]*�3t��j��MPgp�X��q���v�id�/6G�U��Vny�t�UkS�k��P����H6�9p�m8�vV���қ��;YyM&�6�[N�	�6�X��I�l[Dۮ7mۀ��� m��xm�l  m�:@$ ���M����:U�Id�屎����T허
ص�ܐ�v�l /ZG [l][z9m��9m���i��nh(6��6ض��8Hm[-� �;`[d	�k]���-�6�� m:l�;i6I���l�Y-^�� 	 6]�t�n��� &�"��d��sGl�5+�$�J��UUTk�8!�$򥱮m�l�#m�%�\�e�$sU)���PrC��n�M��.�]����@�/�o� �.�KJ��u[mUqz�6�;q%�v���c�AK*�r��Z��ƭ����� p�oQ����ڶ��R�b�x�G�l	�Z�JڔVW�;K�wE�r��ؙBU٪���+m��1sV���3�U�[ec^�j�g�N�2����
�����xjZ㴅�����bU���a.Lٶ� q��څp`���d��j�%C�v����+���>m�6�!l�Uh���J/l�	�'I(������e�T�ց  m��nƥ����l�����rt�젚VR�6�	5����fj�]���B*�Ț��s6B#�%�[eU�]�UQ�SiV��{=�evxgs T�쫧�j�'6���v%�mm��m��]�.�=˭aj��SN۪j��v���R��ba�0��U
%��٥̂����ԁR�U*�h�iJ�u�vĀ)�易	� � m��m���k@��V�
��U@@6N���:k���J���tlۀ��,��f���#��	 m��,��k5yV�[5<�`=�t��T�6�VP���� �*���W��YV0�n��K<�Γ��dW���UmV��ҩI�l#�	{)Y�WUk��죜����7S&�s�vl�@�v9q�p�'If��+�q{il��ev��,�-�#�V�k�[Ę�l�-�H ���ճj�W*g�5��p	[@l 6�ڪ�e1�P�U�.�VÀl �mJ-�i4�Ƌ�u0 �]�oa���6� h��p @p�a�6���E$��m�r���ו`��^m��pHW�����&7]5U�l�J�UUJ��46�m������	�U�m�۵���m:l89�m�%�M�6�A���6� ��β����i0�N�"I  �[��#],� m��Nٶ��Mi&�ڳU�Vک]��T�A���@1��eeV�W �` �l^Ku��0M�c��j��I�j���ٹ�]s+[J���Ix�y:ųk�S��N(�:t햪�� ���x��ӈ�M��$�Y#�Z*ʡe���`���ukg�����@�9���<���� }u�^y@:8���d�⫠����&����8�\�������e��[�c����|����]dѡU�T������Uee[�;s����b�1΃;M�������ݔ;�žuK���q����E�;d
;򲼺�dhl������4�גE���  6��n۷�kslHIdl5�ԍ�Lp��m��8-�E
�x�®�����;��  �B@6U��
���1�U�l�� V��v�lkX �  l����Ӝ�n�m+f�=��j퍫g�ݰ� �WgVݮ����a�[i��-��X`���$ H�g  �7Z�[�� $�Ml�pR���m�߷�I@�� I��     ��I�b�d���@������y����=���  �����b�۲4�Wh*�m�� Ku���%-���)�ll 
�Z�U��]��ƤvһH�v�۬��-��m���Io-ۭ��m �cT�t��]���t��@)�@-A���m�A� ����ľ&�ٞy]��U�6a�f���vx�rfx�zV������y��ݩU�ץ�M� t�9m���9v{m���K/J�UJg�ݥv�d��Y��m�����7�:�HZ�F|=Ut9���Uʜ� �Ž^�Z[R�?���>8����ն�m&g�|���9?��[��Z�y��)[
� T�U��]�ٶ�F�RmZI0�C�9/I),�����U�ehjI��p5W$�J�\��t�'\��������>t�=$���gd��m�F��-�6����m[m��c ��[��h����H:�RZ�5!�U,p6�V��Z#�մ�� �h��� ��/i�����UUUJ�*��h��h��` ���pF�,����l�    f��5� ���� ��j��Ͳ: `��`I6��m��lH �zMk 8-�J��[{�M�a�� �-�   ��� ̉6��)�m�p8�M���(5p�T���Ԫ�1Ur�(C��媪�����Ԭ�ĥ�W��U^kx���	Y�'gEs�u�6�e.fmm�u���T[�m�lI'a�F�$ m��wY5����v����Zm�v� ��cm�7l�kn[@6��[I 8hq��2W��m�n�   �  ��m�h �@i�Y������-��ڶH�맶-NkmmQ��-WF�5�U �l�(	e��4hIj�h�l��k*j����`R�Q�U\��J��4����i�j�˶ٍGYҚ6[xA���Ʃ0�&�<��-�'����@��   z�   � $H��۶�q�@�5�l���ٺ*�%�6��*�v�]���T�V�r�m[@I&NX`��������?� M�?�2�h"�
?����������~0���~@��Q�����(E?E�p���P�Qvh$� �$H�,I!	(�d�~Eڜ ����:��PM�@�����AB	2�l\'ʄ��Q`EN�N"���\������T�
�h
D��N�P� �T������ ��(/��QD�4h \�R�JL/��� x�c�HHI$X��!2�"@dr'M��B$\����!!DT�Q�R��	Z`�!	S`)�x9P��	 �$X�HO� ���R=H�F@ �T{""�2F��@"	^(pS"��P���R��	>ހ ���S��E�Њ�������G@���D6����* @D��a��T��`�����W:\��Ux(�@ z�WA���Q^��E~B(��N�{���ϻ������|'     k      �\����2��9�+ik������6V�s ��iwXC�CN��#+P�.�����nj�Z��QVY�U*��Q2�e��1m��v�     ^( m��I�       ��  �`  �           �    ^��`          �U�ʆ�Ԏ;)��ir��m<�y)��]��N1n���2d6�흍u�[W5�嗴�����=��z䶭vwm��Y6y"ޠ���-IfM�I����+��i�A�����Of�q@�9l�u�r<��,�%�Of{E�cR�l��Z�3���h��
���Y����p魺�U6j��D[�G$cs����7\61֦ۙ�+�Uݩ���
�t>��e穭&;q۵��YM�k��i��؁�����yk��<C�Am)�d5eu��/3�[utv.^�yA�km���W:6m�h֎<�
�گ�;��vڊ�k��';���!��v��fSb�=�j�=v���]+n�t[�:C�����B���H���u�&�5����35�g��@�A��(�<��d�lG��Iչ���:�s����q�t�� ws�R��沆�z�t�s�zQ�k�����#������6���w�Y��M�u��X2ʶ�[l�CtP9��+��"ZB�0o�1�II��2��9��'�&8Ή�=i�r��5(��A�ct�8���ۡj��ƢnS��++ƚ�V��]��Ɗݻ>�L�V��Xh�:��FX�	�89�v괥ʭP8�`�UuTv���I���[3�q��A�h/J�pq�cu�ܨH�2]N�p����೑�ZE���Q��ӳ^K`'v$�Ս6aw���n�m���2f�
;� ��ҝU]��TJ(`|�_�+���{���w����~���� �� �Z��=#�jq���mT2  �f� $ �� �cz+�]{b]A�=�g:�^!���p�B�hw��͋�<4r%V볒�.��z���ܒ�ɺ����S9S��epsF�:آ^��/�֩�ɂ�z6��л�q�۞,�[���i��l��=!r۴���l2� 7L?����w����z���ϗ� �]��v������x�/v6��.y B�" �oD�K��J���Rﳍ�Jhe�֓LRN)�3@�۹�[Қ��-뛚�����s� �#��[Қ�S@��nh۹�r�|xX�&�6�4l��o\��-�s@��4y�a�x�	&<	$4z��m���)�[e4}�6ҹ@f&�y:�Iokf��N�4iݐ�U���m�]Q�@�>�cQ��"��NC&1)�4m��-�M�)�[�74?^vA��7���	�dԓ��{5�_� @`��9�i`n�Vfe� ��<��335x���=�S@��nh��h��@?S���"M�޹���s-X��v�O����b�ݗ#i�	8�jd������h�)�[�74�����7q)m�z��W�θ��ŕ����`AQ3��l�`�y��ۘ%��ޔ�-���ss@��������0pq5���[e4z��m���)�{�K+�LxHh����w4�J��ԟ���zjx�/�x�/{�)B��\��)�J�b��������e4z��g���2(�X�����)�[e4z��m�����]Ձ�� �!n��!j�i�v������\p5����y�8+<G�*�/5!���|h����w4zS@?S���"Hn�ss@���ޔ�-���|���� 	ɪ�J����j���ag�7�;�������e��m��FA�G3@��4]�@�����f+]��9[���0j%X�N�ՠ[�C@���ޔ�=�m*����$Q���9�����ۮ'^,�墻��j8�&H3]�Xݭ<s��dr-޺��h���k�h���E4�2c�4m��-�M�j�-론���8�M�x'3@��4]�@����m��ެV����M�hjC@�ڴz�h۹�[Қ�Vդ)�������-론[n�oJh�V�Vz��RI$�I�{SI�<��\2+�6��	� -�8@    �j[��n�۠�n���:���w�U�8}��ɬlV��v��kF۞z�����J�Y���uf'���F;���P�&:�8N�\p��ێ.۞��Hl6��ݮ���XWgTe�[�7��𻣈t��e�Ƅp \�Wn�S�<9�q�$�p6ˡ��}�ܱ&�/ ��J9_iǹ��� ��6E�sǧU��=��:��n8�o@�q� z��s@��4]�@�������q6�B# �#��[Қ�ՠ[�C@�����<,S�B�&ӆ�k�h���-�s@��4y�XeX�3	'���Z�t4m��-�M�j�?u��<�i�d�% h۹�[Қ�ՠ[�C@����`'� ��%vNz"N-vꮫ�c�N$����w��SR�/"nH2(�7����ޔ�.Nc�3;�JGn�ڰ�Ots-��M�hjC@�ڶ��N�X���0���!U`�)�^M�ʠ�/��P�<P��oCc�0�&��@����z��ޔ�/;V�v_-m<c�㍩@�n�oJh��@�������q6�Ĕd�9��)�^���t4��hz�I���5NH�m��gs�J�=��nM��s��;�㦁�8���)�Q$��i�@�e4z�h���-�M��XeX�3	'��$4z�h���-�M��߳<�<H���{�"�r1�H��4zRʄ��F�	U<���߳l,s;9T2)"�&'�s4��-����w4�X�i��M�h��z�h��h���/�S@=�r���,�������'F�8�m��Bvp�8� 70v�CIp��,�r���̵`g�Xj��0����;>���1Hq�ԁ�[n�}���S@��C@�Y|��s	�����e4l��{���m��^dJ0�N]6�A2������`n��X��V��
'2�윖���a$��$��o]޻��)�[Қ��O5�C�8�X�$�v�7u�{)ړ$u�#Ɯ��n788���t�9�̮cȠƜ�LbR�o]�ޔ�-�M޺��;#Y�F�����)�Z��޺�w4�H�m������Ԇ�k�z�h۹�[Қ�Vդ)��'2�4�5DC���X�����	���[�.T�4�f��]PX۹�[Қ�ՠ[�C@��癞^���@�`�~��,��n!6�r��
��HQr� �`8@ �J �`��M&j�I{:M`˦Cl�8�x*7nӇ6Z1�CsΝ���i�$�M�]4ⶇ�l:0��$nhǑ�N�K���W�2e��fg�5�y�6.ۄ���y�ظn.�Ȍ;!rX嘸�o\t�Pgq�a�vB�YV���C]s��gb(�ѫL���t�ۨ�U��z�Sni�3ծM�ӹ�h�s܎n��Z��i���z�[�)d�s?��|h�V�o]�w4V�𤘚�%<N�տ�癘���a`n�ڰ3;XXv{-�R"I��9�o]�w4zS@�ڴ�k{�$xƤ�&1)C�33ۻ�`n�i`fNc�3;� �������7�1���[Қ�ՠ[�C@�����m��MĤm����9�n���\�:z��g3i�����^�W���@�m�7�6��h�V�{�����kb#�>ݭ,��,�lt��e��K�7w�*����w]*��-v� �;�[lb�Cq�ԁ�[n���M�j�;��h�2�q6�6��#��~�S@�ڴ���h���I15�፸h�V���C@�m��?[)�w_�<|��J�O<v�飔�f^�ۇt���Ge^|�r��9���zr�v���t��}�J����ݍ�@^o7��G�jH�c�4������s�����g�{�H�H�8�@g�O��΍]�if�Z�Q�XT�H0`�`�cE�2	oR�Hk�Y���qL�"\$*8�Q�`@� �ǒ����`��48u��H&P��5p'ԃ��5��R79a�IRQp�tB�*P� ����R Fƈ@�	��%V�#cd���50�HM5��c�L�-�L�PnR03�
9�cs�y(\�J �1c!(l�F��pbZE�
���jΜ��J�k#a����B��%1��`H|5j&�$�	�L`�.s+���&Fg @̐*Ɛ(��`dRr��H@� �V,+M�).Ip�#�!�2��Ƴ�K�: �"�x�8bA0a�E�7�TDJ�<z��>~]��D�(b��{�=�jMI9�{F���[;Ѷ��x���hϪ�;��h����e4
��:��"i���7w�(��T�O�o:�o ��:�2�A*���
��I��y��˭��C�Gz�[d��ש��[��)2��*����7��^^������ϼ�na#j�4��h��Zw]�u��:��
���'�(��t��{�J��馁�:�V9��I��9���CBo��I7��Rd��hl��]�~Z����ƱILbR����T/����,�����Ȉp�d�Z�%S����֖v:����+��� ��5X�lw���?"8�^G&sK�;�W����;���J8������|6��oX9����7w�(��T�O<�MtCc�0��CK�7w�(��T�O�uZ�vZ��� �#��@��Jh̬,}=�a����XlNƩ��ES�Ca3E������D%价���hh��4|�3��d���I"�Qx6����V�V���ꊰ� 6� ��������V������^���O\<N�^�7F{U��b�`�(xM�nFrz�.�i{;�;�d�k����Q��e3�*��D�^�U�����;��y�l���O]�.�6�����V�^hN�c��|7σ�<a�H��JT�t�uT7�����{Ǿ{��?�`�U��s�ս�l�����f�y��3��ضw\㜵�g�59�ǉ�p�=�������M�����XeX�3	$LUU{ܰ��Dzd��x�;�W��t���${~_n<��7"ɌJ@�>̭,fVj��ٕ����a`���DJH�ƘФ4>���oƁ��@�롡���w�@/$}��Hn	��h����{XXQ�	{��������e4޵)�fH$�r$�m[g�y;sKk]u�ʎ�i�sۓ���{V\V�{���P��\��2؝*�NfY3G�n�,w������ax@�D}!ݝ�[��2)�5SN]PX�kBQ��@A0�y�0TH�@YP��JJl�z�X��;��X_�@����a  �9��q��S34��.��f�?~�Ł��q٩%I�B�����XXݯrr&N�d��fXc�ԟʠ�� �����`{��a`s��,5D$�ݽ,��-jiH���MS�;�允�"/B�DF{�~:~�_����3�3-��kgp�D�u����ٸW�\4�K�.#���v����!�k�����|��%��ss!`gt�P�<P���^Vû���?5�-�S)��������ݭ/��d�s6���{X^��L��g�6��o@�4�����t4�瘑X��X�^8�0Ƅ�!R\FAX8
�K�^��IW9ͮ�kK�)��lU%K�3,sN��(Q�_�������`g�_�>����B����V{���W���G2�����.�,w�������^�s��w���^론~^����7q)Uv����;��Gc^L��p%v�����)�78k��B^!BI��q��f��I��L���W�&��v�I�s���	�*������x�7���NjSeA$�9�v��@����P�~���4{���3�/�^Q	/� ����}?��~jiH���MS�?{߬,w����Iz!$DD%3��x�;��v3Z�U*jf����&�,5DB�$D$��w�,g�Ł��q�l%�(���w��gg��"%$m�LhR��hf(�DB������}a`}�k��q:˺�=- =l���I�c���#�|�>:;p4�<r�u���������̨e��e��ܟy��允�ݬ6~"#�g�Ł�6S^�lU%K�3,sN���,/T(l�r��7�ZX�s�%�I)�������MQ2ꜹuA`fmx�3�,�B��Jg�>�=�������f��I�ܷ4XjQ	�v��>��;ܰ��IG�$�3y���O�CΨ��RʂI�,}9��؅�BI!@�G�}�|f׋>�����_fr��m ЋIj&k/�K���ʫz.v@� m� H   ��H���;Fn �Y݆q��X�q��]Xe0�[�2�;�56�u�������9ZD.u��lp�7��yH8��g����7g�����]x���71���[�n����8��m�%�����A[sV;@/k�a����T԰VQR都��}�wp��|�Q*��}nKn-���u�Im�gi7+��R�f�13)������Z�%�q��"*hS5O@��ް�>����;�s��E`H�	`	"BI	/�;��;����UR��j��U���ݬ/|BI" I!"L��W��>�3����D(@�BBBS ����%7US2��#uE���x�9��;?����BU_�����`��0��ɚʙa5E���$(Q=������XX}���a/��=���>Ua���##����@��B���^�{���ϧ1�>}�,_GpME�}�Σ���_l��nx�u]la��a�m��~��������R�Jۀw�ZX�V>�ǰ�/!G������)=N\�*��m�sE��ea|�C"��� �"��q���f���������"!%
d�O�CΨ�i�P9nh�;��;;��̈́��$����s6�X�W�;9-��LBg���3��<��	�@
I	D�w�,ͯ}����Q@�a!)�c����RN~�h�N�����A3E��ݬ,�P�" �"^�s��w'�vw�����N{�+��@�]�Rl4�-v�X�Ìgj��N0MI����̹��1p_�!1��K��#�7�1�Hz���Ɓ��j�/ua�
8ý���3�[�̶L��T�	�,}9��$��$�G�z���_l���y�r�>�idc���By��{�Ϧ��}��job�E�@|/��M�|h�~Z�_-cl� ڑ4��a�!(������`s��v��Q
}��}'�ɩrR�S5-�sE��ea`~IzB�_��۵�����������wκl@5�]�ٵ�D͕�c��9��gc8�.x�]cWc�{��W�;|�NI�ṕ`f��:�g�3g�����a�c�0�29�{�7���d���`{=�V>��z��B�;��n<����2x7ߧ�_m�f�H�=�������`��r��9�u*\�7TXlB����|�����;�g�ReP� K)B(,,U-�*�</� ��}�jI;�O~�3,��̩�4�}9���J=
��������ϳ-X�y2N7�����r��9��E���8��፧�N�o �{���ql�	�$X!-�a�4�1��m�8����{�Jh�tx@�0��Y��s����/G�$���&]S�.h�>����BS�B$A���  +1'�޵`w'�vw���$�=$�HX�Eb� H�Eq��؟��1pL��$�N�����?z�Z��=��4��©����4������"���A � ���Q=�������`}�k�IB �� ����߾5$��~�B�SQ!SD���vw����B��IG�!"IB��ߎ��~�`s��v�ҙ-�ٮ�I���!e��v��.pˍ�!��&��kX`�@�8\�,2J��A���BI2!'�΍�~�9$���۸V1���!
ߦa����F�R$cf�!e��("H�B�D-_ 5���B2���HH�ā$efI�p��p�a��@���#[u����S?��� ��_xb�>޷��[��I�K���2�&cD��$ ��
J���	�
�� �#2	��9�a
$�B��R�-�g
�"'�2P �	0|A���P�m``VS$.\}=����\   ?� �      8)$[+i��_nm�2G	�'&k��Œ��U@uY��[���s�Ĩ@�A�	q=,�	˫�Z�9\�1��T

��	��cZ��A��[     �  �Mm        �          �     �     H�m�      |q�    ^�}��ɋ�k�d#�vJ�c�m��tPt�ه.���ճ���'�sM0��:;]ujz��/\ۏB��` �i�U�j���I]N�1\+,�M�n��>�VtU4���.��$��B��pƽ�j����.�Y��Un��V�!�M�٣�n��ޓ�Y�.k���'�ڮ�ڲ�;���w%����C63�q��\=�q�{*vܳ[���Wvbr�۪�ӊ��J��#�����ٴMѥݛD�*u�0v�I<�+s`��kg��t�NMκ| �]�s�A�:����x�bv�ۣsՉ��([h�rLܪ9'8�ėy�l�����qs]�n6�{E�WNcF�b���ݞVy�8Y@M���~S���D&�g��_/e�&�Ok��!����JA�ղ���c�����v`��)/V�ml�sN���Q��!��D۳n{�Q��8��N���&�u"�\k�y���}�}�7����@�d{h�['���/ml�N��'nٵ��(Q�Sc5���nZ�v�e��J4�k��n\`�LѠB4��]�v����u����\��ST66���F��Y�wh�ku*�M۞	�tFژj�e���sۧkE��
-�ј����r`tm���̕zj��+8N�ni�`ڶB�ݺۂGH	k�{a��[U`�u!q�A�:6nB�M�� ���E�V�Ҫ�e���i܅�MT��,Z�Ì�o�ʟ{s�\��Ɗ�́v�3Z��3�93��=��@�(:W�\�]
 �� �2 U��|�~@N�P��Y�m���&4l�]  ='F�1���g.�����m��	  �����65/#��X�g�tsv���l�\�shb���^��V��������Z������m��s�w�}��m�P�b#X�ƩUNД��\p�]�JJ�:�m�ϛ=V����܆Ŏ}[Llõ�����˂�UA����H9�]��)ג9�O"�^�l�nW��ۘ��mY��[vS�;$u㗶��3��nrv����Z���w��ow�������E�i�ײ��?{�~,�2Ձϧ1�J#�72�����F�m1	Hh�w7���
!L��������`}�k ��Y��Z�o@����ՠ^�M>�31.�>4��4�0�F�F8�hN���	=̽,�+K>̵a�BO�ϾZ���|�3c���4}�MT(���p�;������9���+��T��z�Sn�Epn��ɼ���<���]u��7���+|��9u9������4�hޔ�/u��=���Q2�UPܷT��s�¤(BD@P9ʭ�(E��.�	�C�0����1��!�LV�UòR���@�d��@�H�J�Dn��k���o�X�r��B�$�dܝ��榢B�T�4Xͯ}�j�IxJϳ}j���x�9�idS�jf�j�Q.h��Q�$�}�����mx�3��,6"<���}�� ���MSr6��nf�}�s@�Қ��/��hum��Ȇ&�R6��C�Qu�u��Ջ���f�L����U�6;������"�ƹ�s2ƪ��2�j����x�3��f�����������������M@7����-��iԓ2��w���Dz"���BS'���`{=^,���_-`��1�F�N�w4��f�M��"�|"`Q�U��� "AUX"0Q�0A@�)A���k�g�ԓ����RN^��q.%ɜK�nnq�R
'��`V
�����'����MI;�3٩:y �@(���T{��~�U3)��n[�,�=(� @ �b�{�ߧ�O߽���_zS@�ۉ��Q�����ܶ�G������9:M˻ip��<y����e}�;dX��Da4�Jh���/��� ���
�ؓ��g�ԓ���z)��sU5B��4X��W�Q��"!(�=�^,{kŁ�v��QВD(@�S!�{�ST�&�\�ff�����`fv���I7�����͵`|5�3325T���TXlDyD/С!DJ~���U��}_�32Շc}�pG�� �������O݄?~�mT�N���U4������G�$�(��I/߿~������33-X}�7*Un��PJ�yö��띙�g�=��P�K�q�I��c�u�I��z���iL�����j�ϻXXfe�I%�"!}!���`fɱ��r:U#��:�V}���D/"S&{޵`{6�X�e�؈P����26�I�M'�����Қu����4}|�V9��<�uJ�b'������j�ϲ��Ԕ'���>�)lSU4�j*�fh�;��V�%ܽ8��>�a`|�D%����U���%��"HG���ȵ����M�[K��_��m�  8�UU*���Y�t���36��ɆC7���^.�îom�7f%���<�rXW>+g�kf�}(ۅ��l�ii�q�\K��5��z�B��9����n��;v����;0�Q����b(�B�&�֐m�=n��Vv��s��V��,s��Hu��e�,�g��?{�|�*!�.��S_�)�@Bn���*sl�v���X�N+�:���M�lq]4j]Y�p�w�m������̵`gӘ�BP��3+i�m��F�fffGE)�2�j�q���؄�f[����m�VӶ�y���m��0idc�Lm�f����W��$���[���D~������q��~�-���dfK�u$�U2�T��ߒIyB���z�������o�̹-������q���|��2cQ�4�Z�J�m?~I+��5$��Z�~I%zX�$��r�d�	�)Umq�;�X7l��܋q�C��L����b�nN9�X���{�|>5�6m��o�m���e��ϫ1���"92���Ӝm�٩hZ��J*US5RX�y��;�$��^Kد�J��M��6��6�v���G�%�Qwm��ֿE5SNj���%�>q���W�v�o����?��	~DB��ޯ��m��ߟ8�b}Y�J�d�&��3.�m�mqv�}���m��=�����"*���;m���^�����2�Z&��o;Yl��z�G�"�=�޶���E�$�����$�eJ`ْ	8�
�\��o&��GW]v���5sۃg��eu�YqZu�u!�sb�Vc| ??�ߧ����=�ն߹�vxG�,9��z�>� }����x^%9���� ���7_�?�_�R# �֭�����ݶ�z�[-��;Y��m��;��,�I���\g7V�~�5ٽ�oy���[ �A�V# �v���P�Bs�����6��W��m�,�.rj�̲c0�b�3{��Qʰ ����c)���?����l��m�����m�K�.j%22�Y�e6۽��v�$��(
13����������7�m��[-���	Dow�32��eә�T���1�[�\݅��ѧy�����v�:i���;���� ���q3�nis�\���LGT�m��~�m���oq����ɖ�����~~ n>���u.��8�����9�P��K�Jwo�����m����6���S��B^I/���m�{�����2�Z&��o�����m����y����n�m�<���L
$��"ji��Ԓ�"���y����v�o��]�ݷ�61�� �~P�����w� �{���JsK�G����}�6������g���n�{��m����>�2�������us���v�@xr�����G.'B����~����{�S]pHhq2���W��m�oT�n�{��K2K��-I%�>��|�m�1!�ߓo��\��DBP�e��wg�m�ܭ�m�����	(^�UO�}2�檓%JA6��������y������m���Ԓ_����X�jy&E�$�Ħ{����f^��m�Oqն������ޞq�����J�d�%Ԓ6�QV�o�����F��6۸��m�6x�m�>�wu������[@	�����l���{E�u�I3�  �@�  �� ���-�=m��\�\��;�C���!��f���R�8�a7cDR�x1V�qz�����{9�1v�IW֧��f�\c��m��"�nc3�ۭ�n�.��l����@��{����?�]�&~yl9���`�Z-�	T����v�^���0@�2��b�o{��\YwV��@��Q���m�p�.f������p��F;�������*�ꓙNZ&��m������|��O8�fl�4�o7k���os�L
�"SU6�o����~J�fmx�m������g��u~P�^Q�HWv�����\�!TI5S(uS�6��W�v�o����l��SRI~}k��$�e��ch�0Q�K��m�У�?$%w���m�>���m�{�<�o�$�@�������I���"l�]�ّ��m�ot]�����RI{ݴ��$��6��NN$��U�8z�ˎ�&�m:7fZ�9����=�8��s�s]�؄�$���ઓ%JB�T���}����m��k)�m������Kl�溶�^��}�X�jy&D��$����_���B	P�ʪu@;�@��3�����m�;�V�o����j���������~��s.��0G�m����l�{����"���wg�m�ܿc� ~1�ߪ��2�5�? �;�	~HP�r�έ��g�����e;m���OߒH^�UD��ǒ`أ�jI>NfO8�z��Jf���m����m���K� ~�'ӎbV���ӟsO��#���6gc�ի��\=��1��CqǙ�&H&f�]��͞�M��v��m���:�J<���g����'���*Y2`�xۑjI.��~���y��s�)�$�}���$��,Z�K�-<VH�8&Ḓ퍼��m�q��v�b^J�R�C+��i)�K�(Y"+&��!R�#�&,H9*�0%a$a+Y�T��60R6F��BT��1� �6�3F��5��Hc&E�	DզscK��9$Et�lb�q�dF A�@��d$+$d���0�$�U���N2$�`	�0@�F
��$@�aV$H�# ��p��`�'XHsI�	V�b DWJ�88)x
�8�@ 8���/\�E2#��TH"����g�[m��zs���92��U&J*��������J�ջ��6�ܭ*�m���9�ߡ%3ڿG�$����y)��I�)��${Ӊ��{�\]���ޘ��w�m�����ܲ�!�=v�N76w�s,�p Sض8��ӷ��k��ｾ<G��]Y�M�TWm�e��6��{�6�o������wD�~��ԒK�����lR!�mL�m��7�)���wE�m����m������AkѱRd��T���m��G�}m�f�M��v��m���1M���|���	I�8�~I|�]������7�m�c��5m�]�V$@!Kh@����Bj&�%ʦQ2`��4$*[�F@�HA�Q``�p�M�+�λ���ov�d{����(s�"I��y�\]�ߔOk6�����ݞq�ϻXU���{�1�o��R@5�^�fK/(�8���n.��s���Z�[�Wg��s����gٷ8�1���}1M��7�.�l͞&�m����䒭��ʲLC�LxD��RI~����f��M6�����m���1M$�S�/�b��I�q���G�)5&�n�o��D=��b�m�w�E�m��]T�9X�RRI{ݴ�?z����^��������@=���m�)�6��h�����^�~�٠{�;5$��D�T����wu�_w�w��d�o����1��ĩ	�]I�4���H-�m�    #���m������.x��D�%��7m��i�n$ొ��$�՘C�i��n$�����ug���SZ;<��7`�B:m��,b�Q4Am��ηSպn���JN�kvոӡ�D�e�@z|�t�R�lm�#���X�]\��7nnG����{�"#���wx\�],��ۮs�����c��<ra�}�]Ǘ;0NI{a����v1I�j7�U��z�޳@��X~���>�̀ulnˑ�*�*�Z&&(�zk�yy6ot�P�����E��鱩�27QIӕ35Vs+K�oEo{��/7����OGL�60�r��a�	?���`|�vl�w*���S@��xeY&!�&<H��{����7��{�‷��@vo'	��f�z��Vn���=q���\!��8�c:�t�b��5C�+7���3vx�-��}l1��E�@�k�U*f���m���>�k��ZHJc! V(A"!,Q"$E(�HUB��b0��0��Q`�@h��
-"���^�˺� ��Y�y��H�F�r8$���4W_���u�O�=���:��z����9�5�C�T%
<�7�(����OJ�>����W��#k$�cR- ��Y�{�~,{�Ey΀;5�\��m��BPJ�we�3b��V�g���ˆ��p���Ɨ�Bݍ76O&&6%<��xۓ@��Jh��f����~�0>�mX�z��T����J�oEy΀/7�����M���(Z�Rd��H"��������zh~K�����1�<P��(�e_"D�BO$��C����@��|h��^��ՠuf.�d���KJUX}�����%��O�fO���w*Ϳ���cFp�R�Ŵ�<�]v:��+;v9��1��/b��lp�5J+=A
!8�(y�dw: �ޟ�~%�ao��4
�g��2#	&)n=2;� ^oM���o7���^�����nBYU.���sN�37�`}�V��@��j�K���i)�����У�9���=�>�k
��_<�<�޻4�W0�F���i8hw&��y$Fn�����X�V����>��4��]�z�[̊naE��9,����só�pދ���+ۣ����vD����� ^oM{���[{�E�ř��"D�&B`䆀~���?vV�ɰ>�{���L���:UR�i9m�ۙ�{�
�oE�΀/޳@/	ci���NCC������;2w��9�eX�+��,x6)b&e9��K�3#y��t��<h����[vInI$����Z��g�gv[�(��`���J� m�  rP�]��ƸevpU�uB����Ts�{+v�/<D%F�5C��m�֎���k�2|�������i�'Xnu�d��d0�̓F�N����q�$�pi���udƎ�:�wi�W4��|V��u�T�e�	�˞�/xY��/��l���9�'\7M�[��i���t�eR�U����^.ٍRmO��:�������[`��ש�$$R%"��}��?{e4}}W�;��v�f��\��):r��U����̎�@fF���;�DƐ��i8h��Z���@=�٠w�w4�[�*�1	��@�Oq��fU�߻��?�DD>��]��Y�y$Jd&ȴ�m�{�s@��j�?W�hlm�+����ɫbS����kMr�:2k��OR�+FzIz!�e���)/'R)�<nb�,HRO�^�nh��Z��� ��f�^:��mB1�1%�MI>����(U`iD��W�Q}N�7;���ޥ_�{ɳ^���^DD��࣋@��~Z��>�3į_�4���@?gyզ&��1̺ ��sz��΀���@N�	��SɊ'��4����ՠ~���}�h�O)!��mĤU[\q��,)�x��⩲�=�GFy9ݸ�ͱ�s���G���� y�nf�{�4��Z}�h�]����ʲLC�F`�p�?W�h�٠w�w4�)�\��yR$Q��	�r- ��4����  A�	��{�g�RO��v�C�.�d��X���w]��Jh��h�٠�#�m6�#6	��/t����V�_m�w]��?������@���8�f�y75::������S�pg�ec!v1Zu�E��S#�)�v� ��4����ukl��H��@/�����{�4�ڴ�:�&�IO&(�&��;��h�S@�]�@-�X�8���Kc	T7U3J��OwoK��`��`�B�/�\BQ]��+��L�cUI���4��9���/�B��W�߿W@���Ձ�����e9�o(�Y8X�y:�[�\݅��ѧy���[�Om��Rzi��8kp��5�u���Ͷ�m�w]��)�~�ՠr��uS%Jt��i�����{������z�X�����[l���6�j�6	Ұ32��9���ԛ7wj��͵`upg*ȢD��Hh��h�����m����ui��BE"PsN�33*��J!,��.����̞��I�ʉ�+db�B ��5����)�p#��!@`g@�#��FfI@�H�	�p.�T"EB��@� �Y*0 ��Aհ��TbI�2N��s��9�r    5�      m���h��,����-�v�ghn��Y/l ۵yX 2�.�I�¤����<�:إ/r[J���Uj�U�)	Pnĵa�v�e�kX     ���  nۦ�        l     �          	     rA��      8    ]7I�m�v6�U��ƞ�j�X{9���^�R�:�,����3�g U�uT��^
8��٧b��嶭ú��S��]d2c5U[Td�4b����qY�6J��%�����z���,\�ZΎNnz�m�L���N,b��ɔ�Fn���r��0�r;�gdoc�j��S�q��tlP�sc��ɳ�O ��y��j�]@��)�dں����6�lm8��nw^Olh��;v.mykv��R��181�m��9:8���#��,����kP܎���b�,��pm���*���'H���R�2ڊ�VЧB&qO'���ۃ�{p'Qͼz���s�$[7R���]�=��܂J�$.���5���j�(7�J�Wl�����ɳC�G��K;S��s���T콶s��ʰ�^N-�(����x�ԸY��-�z�G��oF8�f�92\�����q��N���.ݞ�p� y!wIil<�l����{*v�í%�',놛$�[�@	�����49d�X�[�S�3S�}gu�ηa�+a�R�E.��Ul@������7X��]�64�TŲC��W<��+;����=���j�����Y�>1�B���U�8��������6�-�f�v��ݥx�cHMM�i7&�$��e�ζ7K�tJv��(��p��&яO1UOl�e����Y{m%r��av�T�X��^P�)�Ғ�T�+���%:�h��T��q�������<���AC�+���� |�r*t@�����9�s�a����W�E�n������,�a�� @ 2 
�Rq�W8�еT��ce��\���x8^W�:s�dnvʃ%I�Z�nMx�O�Ĵ$���q��G/n�u�a�ka2R�U<@�n�tnnDn����ɩ�M�:�����j덶^:箹���Ľ<�]nKs�Z�F)v��6[�͉�L���s�� |9�L��i�mn��u���A�q����m�����E7V0p�<ڼ�^�����o����s@��h��h���;�둤 y�nf�m��?W�h���w-^�M�d���T�(��Nh�=�ߖ�[l�;޻��S@����M2�UI��;��	��ڰ3���l����V��;�t�#�2D�$I&���s@��h��h������˺�=-
��%/Y\%\��m����􃔌\q�7mv�6x�f�j-/&������Ɓ��V�[l�;��h�9P^E$����?Wj��0b���I�jD��1E�0/J�5'w��@�z�h�M ���V���G	�qh�����m��?Wj��$�m)⌄ĦI�wu��-����Zm�4��c�F�������S@�]�@-�f���sC~}���gC �J�v'[��v�ލ�k�b�wW>{<�2']u�63]�f^�\g�;����V�[r����m��.z�"a'�b�Šܳ��16ffڰ7v��9�����}�J�R�"K$�4�SK�g���S��d� L��]���&��h��h�Ӭn9"�r��LҰ؈{�zXl� �ŕ`wu��9pr����I��%!�~�ՠܳ@�빠[e4�3�3ܫ���AJ9]�>�-\��;�6@ٝ�:"�ۅNM��Co#!����b�PXb���g�@�빠[e4�ڴ������IE&�UX�r��(M��>4~|�ۖh9��\�X������S@�]�@-�f���s@�άyVI�y���@�]�@31eX�rՄDB���P�Nfs<�T�1LRy&(�Zm�4fV2s���-���ri2f�j�� ��f�nl9��v�z�@��;`��Y�®x�]OP��6�~�����S@�]�@-�f�\/*�jJ�5-� 敁�����l�gu�w]��*ɑ�qG�����V�[r����m��9{�:�d��UT����;I&�umX���l����V�wu�&�IO�	�L�@�빠[e4�ڴۖh��=�~{�ߠ�h�%%�����i#v;Y$ڴ�  �     6�:;]��^��t4�F�˝;��l���ub�6s;7"mŸ8�aM&�ӽ��w[r�.�v�wZxy�'g��6��:�q�u;�{ol�;�����y� �/fۅŲ�t�[]�:�9�[��j.8�	��ō��]mp��=6�#\=�K���5,�*]1�����w�绿�wwz~~c5i`�W�e�L��J'`3lvx�k����<��Q�M]�o$���h�Ĥne����h��h�,�;��h�Տ*�1"S�D�`s'1��Q�36Ձ���`\��yR�'��Š�Y�wu�E�����w:��=�CD( &T�l%��qX��v2s��IBI}~Ϧ�}�|�Q���X�'3@�9���%mn� njڰ;���/��}�B*���@�5ӷ<!�L1�������X�c��[�yh��>m�>�V�^�f���s@��Z/qgS����USt9�`�YV�(�BIG�h���s�hԓ�ǽu$�q�� ����m�O�	�L�@�빠^�c�T7����[Vvr$ʩ�UJ&1)��^v���Zz��ucʲLC�b�R-��V����k�nfڰ3���%	f������mZ��[p;��{Z�i�l�M��;b`nz��2n^}77��X� }~Ϧ�{��yڴ�h��9�d��X�&I�^빿g�y���y�����gqeXQ�<n���&`j J�;c������	�%����-�V�F(P��B 4�!V0CY"�Q�� �HX��`�Tr9H?,(a�B A#�$!�R2h"J2I	��e�U���q����:�s�����)��dx�QDŠ_]�@/\�@��s@��Z/qgQ*��U6��; ��ʰ6�o ܝנ_]�@;ڒxe�I��R%o.�ٛO]�J����W(�9�liz�-��qB��%<jd&%2M�]��h�q�"�sVՁ�;mT�*���n�f�����z�^��Od���=�^�;�s@�άyVH�xLS��E�_]�@30ʳa7��j�ܝ�`b�Wc&�LRy&F�Zm,�/u��/;V���""�A�{�n�I��1ܗ9iҪc&��;ܵ`yG��߼���- ��h�[i�b"��Hڜ[He�Q��# Mb�np%��;�B�����Q(��b��9��j�/�ՠ�ey$�8�s6Ձ���1I�5Qqh�j�if�{��yڴ^�Φ'��H�D�'�[K4�w4�ՠ_]�@=�&��)�Q@�T�y���X�����;�nW�w;�,��#D�%�9�s��DD,��|�ul���V��-��VM�Ʋ�ׅ�M�e��h m�  mp 1����itt�ѻ\����u+�,��r��]C�8�:�d�h�ם���J��D�:�4�;^upq��ua:m��/���2  e�Cr�3�pRt��u��ۦ�w8;^L�X8���x���X�2������\��nd�Nv����pG5��W��̛���w����q�>�4��]�w[�y�M� �l��v3��q�Ga������������s��퐣�m�����nW�u�s@�v����*C���L���U�^�����ڴ�ՠz�3����"Kjdz[w4�j�:�V��+��Ӫ��Ci����l��_��-�nW�u�s@����1BI�#�@��Z�ܯ@�n���Z��Թ5 ��W�#�5��^e(��x�V���섘�!��G[��U=A�qh�r����s�h]�@3w�� ����RH8S�u*ԗ�~B�W ^+��c�ԓ��;u$�ە����#c��ĲG3@�v���h�r��������� �Ꝇ��[����[6s2ց��Zey�T�21I�qh�r����s�h]�@����;�5���t&��iEܱ�ѧ��]������j\�7ct���{���o���oV�o@����s@�v���h� �=9W!�8�m$�h�ՠuv��uW�u�s~ď�����1H�"h*i�����8�l�ER�!(K�Pك)��@��h	sIq��B�C"T uL�0��,� ��%ΰ҅ �Q«� � md�#�,%H���aك�1@��,vQ�+�H��𱘇�F*@MhM��♸0���il ��i�L�@c�9 I�U�("$> ?4�@����`��)�|@�x�A����|
�h�B,@8(��)�ڣ���p �
����YJ�ݎ�@c���'
f\�)dR-�nW�u빠w;V�ي�/�@:߼M<x��s!<�@��s@�v���h�r�����O&	ưR��o:��=ؑ7Jիi��[�rv��f����^8�d���LbY#��w;V��ڴU�^������
d'�)�[�vrs���׺�l��Zs�h��yR��'�dmŠz�����h�ՠuv�����2G��$�F�G�u�s@�v����I�f"�<�rw�N���g$nx�I����w;V���Z�ܯ@��s@����74��ȓI��\�ݛ��%���t@&�Ѝ���{)�B�b��h��1�H4�G�k�U�^�o]��ڴUŝLlO$�%"�=V�z�w4�j�-}V�{�|M<x���=޻�s�i�M��k�:�V́�)ȓ*�It�)USJ�TC̬�`n�k�8�M��ܼ�?z���"<s	����-}V�����j��g���AB!^��6���}��YZ��닉�b���mb��.����X+j l � ���-�����shWn��ͳ��j�']��Jv:;:�\mZr�)����=pt�a�Z\q�6�Z�u�uQ��JbN^�3m���PQ�{6{nA�l�c'$��qQ���&凜�����gr��r�7+�ۇX�u�D�"�n�Бi
��I�͘~U�<���-�q&d%�nsg���8�c�����v:5�6��Z�۸9%�ҠGc�O'�!̌Ry&(�^��ܯ@�����q��������eT���Kjdz�w4��h��@������*�#s�M�����Z���?+r�޻�ɍ�A��H�_U�~V�z�w4��h��:�؞II��h��^�o]���Z�����cIU�.&
U^g=�Z�_]p/nD�#�[q��m�=�0�"��`��U�x/jֶ����V{=�`fOqꄸ�纶lꝉ6�d�Mґ�U4��{��!%��]K!D]��v���ٰ3;��}=�XC!3�x18�_U�~V�z�w4��h��yR��'�b�E�~V�z�w4��h��@�����2,hq%�52=޻�s�]�@������(���܉0Un�(�z�6sp����w�7������leku�j�ń�E�8�m&�~�~Z���y�'и�w6Ձ���1Jj�Q.XUS�3'��T%�>{�f��͵�w>�@��,�cƞGI�qh��^�o]�=��y�7��Z�ՠ��������G�[n�����j�?+r�����#cQ)�K"�4��h�V��[��۹�o��߿����t0D��bm̛�t�{sd[tk�g�풵��e�c��.s�r;����q���-�+�-�s@��^��^_*C���LQȴ�ܯ@����uz�ՠ~��bt�48�(���m��9wW�Z�Z�nW�9u����Ʊ6�s4>�3��͛vw]�ǘ�l2#��%���@8s�o]5$��͞�Ó� �DR=�j�?+r��w4]���U ���JF�hP~d�2��0vɶg$�&�����s;m�m�w4u�q[��AH��ܯ@����uy��}������o5<$!<�@����uz�ՠ~V�{|�#�W2����*���rl��Ѫ!BP�bɰ7wmX�{��B���EA-�M��ڴ�ܯ@����uzb��#�I�7��[�����9wW`fOq�b�ͤ�"!B(6 ��H �0`� ��$ R21wp�ã��~���RK�7'f�l�U����  ڶ 6� �  ��rQ�Ō��P�h��q-�㞗y��c����/9���������uk:�G�N�SŻh���л���Hn��7ѣǱ��Kyo3�r��'c��3���ƌ%�V6g���\�ݭv��3lL;�+Xz�l�۱��l��R�v^����ݛ�|n2�@� �m�1�vkn�����1On.��;��u��,J�'n]��bK��=�w4]����@�������mF�3i73@��^�k�<œ`fw-^�I6wL��T�TKi�)������ܯ@���˺�|��MJ�)ʒfa�*��$�y�f��͵`u��6fe� ��șr�7PUP9U6	���X�6l̻��nW�_z�I��$#q$�5z�Y4�+���Lj���:����S�Z8�ë���2H�%1�dRf�˺��w4�ܯ@������L!���a<NcRN��Ѭ���h��O�vw��ܵ`u��7�DCf-�B�ʢ�u<��f������۹�r�@�����0��2,hqQ���۹�r�@����[��WXڎC$f&�Nf�˺��w4�ܯ@���ֹ���"i7���a��:�{c��9�d�q:�]�a�6N�I{f��i�v^Dԑ��"��۹�ۖh۹�U�^�긳��x�BH����,��ٻ�j�י�`ffZ�Q
Az���x��I��}��Ws���42Q�A�Q�I%7�{j�7z��꜉2�T�M�1,���*�@��� �ܳ@�����ܘC!3�x4�z�w4�r�޻�]�����-��N<�]�Z�u�x9�9؋�n��e4bü񂁸�28��<2$HF)<��f�_nY�[�s@���޻��z1c�dX�4�6U*�3�j�f�͛w6Հ_nY�9u���!�����U�^�o]� �ܳ@����2�/#jF�MH�z�h���tjN��T ��9�jI���uL��.J*�]T�>ŕ`lF�o י�`[�s@;�I�,i'mH�m���M�UU�t���z.�D�r�/m�1��η'M�+z���E�'�h���/>�@���_nY�_q�dx��ĲG3@�Қ�w4��f�o]����L!���a<�4z�h���w4�)�v^�eH��Ԟ9�G3@/�,�-빠^�M޻��z1c�dX���&I�[�s@�Қ���N�ӹԐ2� G��[�� ��BL�e�!�H$H�HIKX���bB�K5�J79�!IB�"D$$!�H��HE#		�	�2�PȐ")dY��H"��b@��0c�С@6BUa���Jd�P"�]����R1H��JH��k+#�Za���H�ŐU2�dB ��L�ԀA���dE�
@3_c��@���B�l(�s�!	6���� ���!LC-c���'5>\�H�$�� $R�F�)/�e>��Q��o}�     m�      �:,$I�E���6���c��5��s������U�땵��P.[��r��*��m��hت�������].�jL�Ԃ�M��L-XԵP    5�` �oM-        �                 $     �M�      8    [�ۙ����q��������g�m.d�6��^B�^[R�B���+Q�uV��࠹��۱����v���c�'rc5US�2�[�Ͷ�U���HFq�f uSt��1v8����g�U����Cn��_S�;km���&Qآ����<���P`��$:���/Rkm+4�d��.���G����W<\;�ٓ<a'4�2[r4�ܘ<Ol�����{�ax{a��v�-`�^[�J� ���YN�4���oa�m`תN�T=���'Wcm�:e�:��/12v��u����hQ�Bi�9v�I���<�q��3�A��N6���:��S=jKn֢�21�0�7j���J�����I\�q�gl�jȾ�:Umڀ�!�3m�vU�CԤ�J�:Ӹu�c�˲�d2�2��lr7Q��=3�Qq�a9�l��D�n�v3g�2q'NI)C]��=/)Q��{q��z6�=Y��u�����gl��\��a��{ml���I4�l�Э�UU�N�y�dt�6��c����9�e5�d��Oc@�f�]��ŭ �nB�� nM3�9��gUn�`��C���=�����ƻ��M��ۓ�K�#�-�<�:�� �t�ɳ����GY��$��
���Ѩ�����s�äZ�V8
% �"��(wT�c��W-���A`#IHlXiU�Uf�6���.����2�f��9�L��Ae�zi�UU�nP��sA�2�c�<P�D�"6�p2 q�C�WY�x�9�KnsUM2��C&\r�I�YRD �� -�8@   m�`����v�R�3�n.wc�nۤh��h}���]����N��xG�8-�
��v�����Ķ�jӥ�=���v���ӕ����[5�4�X�=E�b-��yl�[m��2P�j)�Ms�����G���ūF��E�S�����nGHO+��c���{w����ھ*!�3���N-�1��u-t���-��op�[���^Ӛ_a�òT�ִ�UV��Қu��}�@�۹�{�L��ڑ��@�4�w4�r��n�}�M�a��ɒ1LD��I3@/��h�w4�Jh��h���H�<JxID�I�{m��/�)�w[����4�;�,�"Jx�I3@�Қu��}�f��s@��������o׬`�4�]�wu[�;�x�d�]�<n�{<�]'1�����ַ]�H�$���fnڰ�U��fZ�I(�̭,��MkeQJ]R��U4�$��;�@v�i��33��F��ޔ�;���?{Ѭu�,x�b$�4m����;�����4�.�����m����Jh��h}�*�RID>����2��qS.���@�4�w4�r��n�{�4��Lh�H$�r$�m����rt�a(v�x^8�'������)��GY�QLD��I3@/�,�=��h�S@�s@;޾BI��E�'�h�w4�)�w[��ۖh�w�Y�)��aUJ�ϻXX�e�5BJa%
d�qmX��V>��R(���
�2�P�I�n�Xۋj��3-Xjw��h��|�!1�1�	� �{,�=��h�Jh��h�cm�q]���t%=��d�F����^u�{v�R�e�sX�d�k��0E���bX����I��%�bw�צ�q,K��}�Mı,K��Γq.��oq�����֡9U[�{�7�ı,N���n�Qc���b{߿l�n%�bX���~Γq,K��x�L��L��2ֈqS55-˖M�f�q,K��}�Mı,K��=�&�X��"b'}���&�X�%��m��\!2!2���찙c�ʪ������	���%$)�z�L�ı;�߶i7ı,N���n%�`q �"�N(��Mw���K�2�uiM�!7PUST9UW�&BbX�ｳI��%�a�#�����%�bw߿l�n%�bX��t�t���{��7����G�s{a���U���i�Ӝ@�
��f�p�a3�Nɉΐ�8kz|�T�L��uJ�p��L��Yܽ.�X�%����4��bX�%��=�&�X�%����4��bX�'��|��2̙n1q���Kı9�{f�q,KĿ{����Kı9�{f�q,K��;�M&�X�%�Ӿ�4�U*��"�i\.�	��	����7ı,Nw�٤�Kı;���I��%�bs���&�X�%��{�RviSR�Ԍn�*���!3�%$,���Mı,K���M&�X�%����4��bX�'1�c��n%�bX���O���Z��Qn�����{��7����n%�bX�ｳI��%�bs�=�&�X�%����4��bX�B�%b�!8J�o�UU33UUURT�Ѵj�q���e�X1�tu�m@m��	  �lm��2p�Wa�Y2ˑ=m*�ݩ;l]���km��Y���rd��9���:/����̼�N��vo�������NL���+L��#L�ӓ��x��=v��Yִ���� ��S����n�p��p��WcE���t�<�dI�"7'^Utm��ѭp����{��>|�ql���*��-ٽd:kc�g7&v��Y6\��vSN5��j����d2V�{���oq���}���Mı,K����7ı,Nw�٤�Kı;���I��%�b}=Mn���:L���*�\.�	������7ı,Nw�٤�Kı;���I��%�bs���&�
�*I	��o��n�	����)��\.��bw߿l�n%�bX��u��Kı9�{f�q,K��=�{:MĲ!2���5K�d�T��uJ�p�ı,Ow���n%�bX�ｳI��%�bw�=�&�X��Bb'�{�Ɠq,K��s��I��!�ɖ��Mı,K��i7ı,Nc�ǳ��Kı;��f�q,K��;�M=�����ow����P�kc �D���v�C����I�ݻ��O��&��75M:UJ��E"�i\.�	���ݝΓq,K���Mı,K��4��bX�'}�l�n%�bX�w=��f�jT�H�3S5W�&Bd&B��٤�;�#�*�� ���E	D��
!�A`2l��`: 04��:S�2�22B~:�'"X��5��n%�bX���l�n%�bX��=�gJ���I	�����T����%���ZMı,K���M&�X�%��w�4��c��"b'q����&�X�%����+��!2!wL��T�UH���\�i7ı,N��٤�Kı9�{Γq,K���Mı,JB���p�Bd&Bd.�&�e���&Vs��g94��bX�'1�c��n%�bX��}�I��%�bw�צ�q,K���Mı,K���LY�8�%�*�3���<6��^݇g��[q�䭝��NJ���h7+ւ�p^ӭ�k��{��ı;��f�q,K��;�M&�X�%��w�4��bX�'1�c��n%��	���lI�]47LN��W�&%�bw���&�X�%��w�4��bX�'����7ı,N��٤�Kı>�{�$�i��d�q��&�q,K���Mı,K�w��t��c2$8
�S@R!��7Q;�sf�q,K�ｯM&�X�%���OR��L�7.I��&�q,K?9����Mı,K߽�f�q,K�ﻯM&�X�%��w�4���	��2�E;5CR��H曚�\ı,N��٤�Kı;���I��%�bw���&�X�%��}}�&���{����~����əhUn�+/=h5n+(Zv�^/���|��xGD��0���mq�����UT�-L����/�L��L�����n%�bX��}�I��%�b}�_oA���&"X�'�{��&�X�#!g���*f��r�j���!2��w�4���#�G`�'=���j	 ����4��H����j'�%��8�͖Jt�USTUR�\!2!8�篷��Kı;��f�q,�1�Ͽ]&�X�%�����I��)��	�5h(M�*)�uW�&AbX�w�٤�Kı;���I��%�bs���&�X����Buݝ���!2!ohؓT�&hn�.3s�I��%�bw�ﮓq,K��{�Mı,K����7ı���\!2!2ٚ�e�IU.��D��Ģۛ<8�rmvٳ�z����ylI�+خ�8o]�빶�*��w���d�9��f�q,K��9�{:Mı,K���4��bX�'y���7ı,N��z�9�3sr��2i7ı,Nc�ǳ��Kı>ｳI��%�bw�ﮓq,K��{�Mı	��̹jvj��SL����U��	�X�'���i7ı,N�=��n%�bX��}�I��%�bs�=�&�Y	��	��U.����jfP���	ı,N��4��bX�';�l�n%�bX��=�gI��%�b}�{f�q	���e��j�'.YU57�+ı9��f�q,K��9�{:Mı,K���4��bX�'y���7��g��t�w������Cm�0��uL
�vv՝#أm�T���m��'�}� � m�Y�kU�\̶.�6^����U�y�3���x��Ń��:ڍ��hM;�6예�+U�p=���/V��ѻp�V��+v�n&�vB;0��lbld.�ck�n�i�L�v���pv��ME�W������ �Tu���w��CrX�X���j.^���ﹾ?n�,���s�szHxlm��s�I�s���&,�!q����s�%:L���*�vHL��L�����&�X�%��}�Mı,K��}t��bX�';�l�n%�bX����K�Ժ�Ң��j�L��L��n��n%�bX��;�i7ı,Nw�٤�Kı9�{Γq?��LDd/e�<��3Ct��R�\!2!X��}�Mı,K��i7ı,Nc�ǳ��Kı>ｳI��%�b}���I��!�ɖ��Ɠq,K��{�Mı,K��q��7ı,O��l�n%�bX��;�i7ıe�kN��N�E"�i\.�	��Nc�ǳ��Kı>ｳI��%�b{ﱤ�Kı9��f�q,K7������ߍ�Yh�m�mu�����`)��pQ��8'd��ε�%s&E9��fJ	˩��\!2!2ٻ�p�Bd%��s�Ɠq,K��{�MıL��]��ڸ\!2!2�36�]L�KS2�4�L��L���ٸ\�)���� �Y ���D!��B�%hi����K���i7ı,O�����n%�bX�w�٤�O�8���'q����j�'.YU57�&Bd&B��q\-ı,K��q��7ı,O��l�n%�bX��;�i7ı,Oc�;�Q$�I�U5EU+��!2!vw'kI��%�b}�{f�q,K��3�]&�X�%���^�Mı,K�<)r��P:TS&f��p��L��_f�&�X�%��X����>�bX�'}�~�Mı,K��q��7ı,����������籿�c�Q*���Y]'&��lqxK���Ǔ�s�GxuvU�u��ݭŅ�nrm>�bX�'��߮�q,K��s�]&�X�%��{��t��bX�'���i7ı,O��y�3�d1�2�c��n%�bX��{��Kı9�wΓq,K�����&�X�%��g��M����"X�=��KTR�U"�T�;��!2!d�g�p�ı,O��l�n%�B��)>�I�ci�0J��]G_�Aq� ��`b|�Q��^mHe��")"��n^���,7�Lc��	��Y�#A0�`�tmޙ�^+�UP"�(�bt�� /�t��Pz+� �v$ � �Ƣ}�νt��bX�'���p�Bd&Bd/��[�e��PH�nq��7ı,O��l�n%�bX��{��Kı9���I��%�brw'j�p��L��O@��t�jI%��%�M&�X�%��g��Mı,K��}t��bX�'1����n%�bX��w��p��L��Y��fZ�U2G3L�U����uv�Ǯ�ݹ�F�q:�]�a�!;Fi���	�c��p�������7�����}t��bX�'1����n%�bX�w�٤�Kı=���I��%�d-�Mf���� ���S�\!2��=�{:Mı,K���4��bX�'����7ı,Nw=��n%�HL����R�5.��TS*f��p��V%��}�Mı,K��}t��bX�';���7ı,Nc�ǳ��K�L���R�2fh,Ni�+�� �,Os=��n%�bX��{��Kı9�{Γq,K�y, SC�(u3����Ɠq,K���9�C�-�1��&�X�%��羺Mı,K����7ı,O��l�n%�b�;Y��p��L��[���s���`��(ݼ�z���a�cl;�l�ph8�1IGkM�ӕӗ�	NGF/����Y�,Nc�ǳ��Kı>ｳI��%�bw�ﮓq,K��s�]&�X���>�Pw�F����_=ߛ�D�,O��l�n�c���b{����Kı;����n%�bX��=�gP�Bd&Bd'�fm:u5$��̡�+Mı,K��}t��bX�';���7ı,Nc�ǳ��Kı>ｲ�p��L��]�y+A�L�:N\�ji�7ı,Nw=��n%�bX��=�gI��%�b}�{f�q,K��3�;��!2!l�k4�2] ���U�n%�bX��=�gI��%�b}�{f�q,K��3�]&�X�%��羺Mı,K*}�%�Hؕ���
�!Ȱ�8wy�s����cV(9^Gg��̝]$�t� �� m� �>� ���ݷ=u�s�mx�;��i۰���1t�8H'a� m z����s�)���m�a��gt�;4�Nmi;��)��^c�����X�K�e���i6�ä�ڳlr���C��Œ�k�m5���{�ěiѝk�c2�X�=r��ig<:����EJ��{�}���`��^0ʥ��vS�j�����y�r9m\�a��84�l�vt�R]nW��ɉ��Ȗ%�b}�߶i7ı,N�=��n%�bX��{��Kı9�{���	��	���jZ��]%��:���Kı;���I��%�bs�ﮓq,K��9�{:Mı,K���W�&Bd&B������$�T9��v��bX�';���7ı,Nc�ǳ��Kı>ｳI��%�bw����	��	��fZ�ꊡ�*)5WI��%�bs�=�&�X�%��}�Mı,K��4��bX�';��\!2!2�L�6YH�f���I��%�b}�{f�q,K��;�M&�X�%��羺Mı,K������	��	���ٙr��)9nf��R�!�w��]�:6r�s���`�U�ڗ�lp횈��G/e���{��7��;���I��%�bs�ﮓq,K��9�{:�I�LD�,N{��Mı	��|�W��L�T�r�uE��	��K��}t��T���`!4
P˸��bc�>Γq,K�����&�X�%��w^�M��0�!zu5�%�@��j�T��,K���~Γq,K�����&�X�%��w^�Mı,K��}t�!2!2�j�L�ԺM�T6:���q,K?
9�߾4��bX�'��~�Mı,K��}t��bX�+�ݝ���!2!oUjZ�.]���794��bX�'y�zi7ı,Nw=��n%�bX��=�gI��%�H_f���	��	����ڤl���)x
�û���{pi�<�s.<�<=���������j:�7
6�����{��9���I��%�bs�=�&�X�%��}�ʄ�&"X�'��~�M�d&Bd-[���*�&��H��w�%�bs�=�&��#���bs߿l�n%�bX���i7ı,Nw=��.�	B�p���]�f��U r\c8�s��Kı9�߶i7ı,N���n%�EA<��31;��wI��%�b}�{Γq,Kľ���t�jI%��C�W�&Bg�I@�"{����Kı;����n%�bX��=�gI��%��Vb'=��Ɠq)	��'�ׁ��R�D�,�T\.�K��s�]&�X�%��s��t��bX�'���i7ı,N���n!�����?����.MG@2� ��rz�n��J-��
�����ñ;@����Vmۖ$IN�UT����&Bd&B��O��n%�bX�w�٤�Kı;���I��%�bs�ﮓq,Kļ�I�n�u%����p��L��_f���� �&"X���i7ı,N�>�t��bX�'1�c��n%�bR�V��R��I,Ni�+��!2��w^�Mı,K��}t��bX�'1�c��n%�bX�w�٤�K�d/�Y�H�j�Jt��\�p�Bd&Bq9���I��%�bs�=�&�X�%��}�Mı,�A 	B($�B(�b�A� ���� &5��ޚMı,��][���:UTMU
�ST�L��X��=�gI��%�b}�{f�q,K��;�M&�X�%��羺Mı�7�����+�ލ�������tg��d�	�v6�]�;���NvݴjK5)l�8#N�d'!AC����B���L��]�{��pKı;���I��%�bs�ﮓq,K��9�{:Mı,K�I��6�MI$�3(sJ�p��L��Yܽ."X�%��羺Mı,K����7ı,O��l�n%�bX�ǧg�q34U"S�K�.L��L�ܬ�p�ı,Nc�ǳ��Kı>ｳI��%�bw�צ�q,K��Hw�t�)�)����;��!2!v{��i��%�b}�{f�q,K��;�M&�X���D���I��%�b�o��s)7RP��j�L��LO��l�n%�bX��u��Kı9���I��%�bs�=�&�X�%�����������E��u1��y:��\����dj�ꠠm�  &�  k#O��0j��7�k���V�9��v�V���OnzƠ6��v��ߓ�"�86}lq��Ƌ��������ږ\6솹S������3�g���v��3��:P�<��a3��+z�\聧�b�Y�e�K�Ɗm�ڹ���G�9��+�әw��Q�{a���U��j��� x��Zv-�te���]�p�<��]��ɸk��'"X�%��ߵ�4��bX�';���7ı,Nc�ǳ��Kı>��+��!2!}�͊ESUMԉ��fi7ı,Nw=��n%�bX��=�gI��%�b}�{f�q,K��r��\!2!2ك�-jUL�UB�3���7ı,Nc�ǳ��Kı>ｳI��%�bw�צ�q,K�w+5�.�	���)d�MNB���3�g:Mı,K���4��bX�'y�zi7ı,Nw=��n%�bRg�;W�&Bd&BkLͤ��ԒK1��&�q,K��;�M&�X�%��羺Mı,K��q��7ıL��n�\.�	��;Y��L��ne�AU�qn���:k`�.nL�ϫ�:��a��甄���՝��]]�%o����7�ı9���I��%�bs�=�&�X�%��}��R},K�}��I�!2!{P��t�)�)����;���%�bs�=�&�جE΀�GN�j%�����n%�bX��u��Kı9���I��%�b^t��0:C�(l�����!2!}���[�bX�'��zi7��1;����n%�bX���c�t��bX�'��R�)r�$%9�Up�Bd&Bd-�_��q,K��s�]&�X�%��{��t��bX�'�����Kı>�}�H�j�i��9�4\.�	���Y�I��%�bs�=�&�X�%��}��7ı,Os���n%�bX�wڪ���̫Q<�[�jƟ<k�ѯ)��vhn���'�̩���..����u�l�&�X�%��{��t��bX�'�����Kı=���A�?"��Ef��(]�ix���
˩��I�7��)���X�'��zi7ı,Nw=��n%�bX�ǻ�gI��Bd&BkLͤ�i�KS2�5p�B�,K��4��bX�';���7��A�H0��Ш` (d�M��5�{:Mı,K�w�4��d&Bd.�@�nT��T�NXMQp�%�bX��{��Kı;�wΓq,K�����&�X�䘉����p�Bd&Bd/j����N�MTԎ��7ı,N��ǳ��Kı>ｳI��%�b{�ﮓq,K��s�;��!2!?��Im�R:N�����]8���n�a{v9vW`ۮf�N8W���u�oa�ܼ��>�����w���oq�����4��bX�'}���7ı,Nw=��n%�bX�1��Mı,K{F��MˠS �ӪW�&Bd&B��]&�X�%��羺Mı,K�=�cI��%�b}�{f�q,K�}�����&����;��!2!s�ﮓq,K��w��n%���"b'=���&�X�%������K�2ك�-jUL�UB�T�;��!1,N��}�&�X�%��}�Mı,K��}t��bX�Da ��X1,JH�Qj�S;���{��p��L��Y�m
|�NUK�9Ɠq,K�����&�X�%��w^�Mı,K��}t��bX���w6nL��L����M�a,���AU�d���ZAՇWb4�f���Fœq���;O>����G��������,N����n%�bX��{��Kı:c��4��D�K��~٤�FBd&B���r�f����ꋅ�ı9���I��%�bpǻ�i7ı,O��l�n%�bX��}�܄�L��[�Y�t��t
j��uN�pKı8c��4��bX�'���i7ı,N�>��n%�bX��{��	��	��qj���$�m57q,K�����&�X�%��g޺Mı,K��}t��bX�&"tϷ�p�Bd&Bd/eK�MˠS ���M&�X�%��g޺Mı,K��}t��bX�'{�Ɠq,K�����&�X�%��P�?!<��$ct �e�R$�{RQBXa�2��0���L��&3�u�$ eRe$pJ��'D`�m"��k���A�2or�U��	$$L�@	\crS B��0JZF����� �P�4�
�b��������ל     6�      U�Y���%s �;f#k+�6�5זt��D� �Uڴ(�T�xZL��<�(-�s����Y�+Ur��Q���T(VUKh��n���     ^�M�  rY@        �`     H           	      �l      �    t�'�$��h`����n��bJ@뗝جjh�z�8�`�9���H�t!5I�K��������T��;FyM��`������ntd%�6Y�R�N�J<쳝-U���zI-v�PJn'�oej�y ND��C�vwkl��.7"pn�X���N�����vj��f@��&Ό$c�힚�\.�ri=m�^�E�u.����vi�EY�m��q��el�s��s�<�5p���#��B����%��HZ�N��&��"��נ����iq�Dp�u�ܝ� �h�m���t�J9�.�7q+�F��ե��u���/�rs�6ݶH�vxݥ�T�Bn�.�㎸�@�D�BPM�5�n�L��2ؓ�+nն�����//Ta��Il��[un�U���j������mJ]��xv�{{Yy�m�nM۷mî6,�ő�Sa�5��6�KՒ�;G^0�ʃcv�n��ϗ�|��F�P�b����X7K/crت��-��\�Ne��a��u��m��OUӍ�].Ȫ�pp��om��5b9�:�󍛣�Uj����Yi�OHsj막�R�[�t��ΰ�1r��s�Rm��s� �s�sy�Aƽ�������n�=��_gTr�x�8�x�Tʁ�c|���*�u���s����7d�׾����GN�Y���	WY���V�vr��s�D���UL�]r����W+s���c[9L�3j�S��:��L��:!Qz	DB=E�	Dڮ�&Wb� �/�B���'Q��;��8�1��9�q��d�"7k�&�j�tu`E����� H ��l��e��J�r\Spi��8�Ƙ;���Î.��L��<����[ny�hH.s�����zؽ���MX7#)I��s픭�ֶ��\��$|��<:wnn���pb˒6���6^��ղq��Q��vgm���|����t��^���=��F}���{��9P>tD�D��b;t�s�G�]�;��;�8��.���8��8o]����U����{��7���g���q,K��w��n%�bX�w�٤�Kı;���I��%��_fе�U2MU
�ST�L��,N�}�&�X�%��}�Mı,K�Ͻt��bX�';���7Ĳ!}�Z몁L�9R��p��N%��}�Mı,K�Ͻt��bX�';���7ı,N�}�&�X���Mi��ʦ�ҩmK�9�p�Bd%��g޺Mı,K��}t��bX�'{�Ɠq,K�����&�Y	��g�n��fh�	NY54�N%�bs�ﮓq,K��w��n%�bX�w�٤�Kı;���I����oq���s��[8X)G+ �n�,����6ə��&2��ؓ\y��Ԓ�:A5SR:�p�Bd&Bd.��ٸ[�bX�'���i7ı,N�>��>���%��g߮�q,KĽ���nS"��m����p��L��_g��I�mF8���'y�z�7ı,N�>��n%�bX�1��M���*���^�<���3@�A9�T�L�ı=���t��bX�';���7ı,N罍&�X�%��}�MĲ!2�Y�H�j���"s34�L��� 1�׿]&�X�%����Mı,K���4��bX�f"�/�w�&Bd&B����J��j�Y&q��&�X�%������Kı>ｳI��%�bs����q,K�����L��L���NW&�&��m�l�7���+���9�����rp۴1��
6y�ۘmۗ[Xy������{�K���4��bX�'9�z�7ı,Nw=��n%�bX�1�{MıL��Mi���T�t�[R�i\.��%��g޺Mı,K��4��bX�'s�Ɠq,K�����&�~����w����������p���q,K�ｯ�I��%�bp�=�i7�z@�#���J�0�X�	���@`�AѨ���{�4��bX�';���7ı,M�,�T��:USTT�p�Bd&Bd.罍&�X�%��}�Mı,K�Ͻt��bX�';�zi7ı,S�-Zdc��n����p��L��}��f�q,K��3�]&�X�%��w^�Mı,K�9�cI��%�ow�����7�X���z�Sf-U������\�]Yw<y\��[d��W]�cm�$.&3�I��%�bs����q,K��;�M&�X�%������>���%�����I��%�bs�}��3�TU2�Nff���	��	���z\.�K��9�{:Mı,K�w�4��bX�'y���7ı,Ns�臩�S$��R*����!2!fVl����bX�{�٤�Kı9���I��%�bw�צ�q,K����!�\�d����UU��	��	����+�Ȗ%�bs�ﮓq,K��;�M&�X���aBR ��XE�0P"EXA	 5΢w:߱�&�X�%�ON��.s���8���q��Mı,K��}t��bX�������O�X�%��g߱�&�X�%����w-��U��c�鎌�`�U����ut�^���n�u��F;쐝�*�ٵطjV����������4�ս�빠{zS@���ZƦ��G��o@�z�hޔ�;ޔ�{.Pm�(%�q��빠{zS@�zS@�}[�/���&�ca��L�=�)�w�)�w>���]����0�d�DFbm8P�<P��@_oR�3�x�}��TUTE"�dq������jo���|� m[ l ��  �`�j��V�-gJ��4�HB�rμgT�����+����6��b���"�]+r��۝�Z�{tH���\`(�m��v)d�4[��jX|Rk���������sKlj�9q��zm�R�;Eܔ�	����4��ѣ�hn8Ww����l��S�u��G��a݆#F�w�s���n6{v�۩������Oz�U�6�~�ĺ��Z�>���K�3����%���d!��?^����4��4�ս �ˬC�524�������4��4�kz��s@�����ۑLOCR{Қs�f��w-XlB�	<ܽ,�-۩%��	#��s�ށ����=�)�w���z��Rɂq�ԉF����j���.����E+��v9��z���鸤뭹T�AA�#z��s@�Қz����ɠ_Ys.M�����ol�U�%>^�/z�M��t<ޙ�.���/��&,�H��M��}V���eU�
nm�7+K燐e<��Ʉr-��ɠ~�w4�)�w���?w)�R`Qbm�&���Z�6%��� ��k�>}̪�8~�!�]p�,�[t<n���ݜ�D�]"��n��h�zW�lq�j5n�ƞ&�hzS@�_U�z��4׮��SSi�"��&��4��Z���@�z�hzS@��c�1�fbds.�ǽ�4��*'ּ+I$���:�M�v� ����lp$�&�����:���޾�@�[d�/���&�ca��L�-�M�}V��ɠ~�w4��~�#�M�0R�]��z����s����a�:�`@.5��9k/��v��0�~m��_���<̪�9��[�8�w+K��&P�d��I<�G"�=V�4׮�oJh����b�S�Di�4׮�oJh��U�M �wZN�Y4����sTXlD(I=ܽ,�;�'׽�s�8��
����b�Hǂ����5$��޸��1�OCR{Қ��&�����k���3��~j`� ��ȓI�z�z���תk��d˔�Ӥ�p=�v����2Vmۖ�k$�L��G�r���?^��-}V�����{�r�m�9����4ץ4_U�w�)�z��h�\˂p1����Z����M�m�@�zS@�]�L$P1ģ16�Z{Қ��&�����k�}|��*Ǌ
8d�I�m�@�zS@��Z{Қ�3
vI1%$��T�)dǂ�+ʷa`َ� �H �    m�tv8�ChՊTg��Ψ�[4��c]p���5���<{tF���MɌ�.޼<Z�z�a�[�`�:���m�� ���uZ���ù�r?��=w���.l��+�Y0gӓ6� �tX�&����	�r��s���ٽ�vB�c$����.m��X�ݤ��l�%��w��������?�|�N��]okg�3�������';۴jK4\���LX�q�� �NI��~��-}V������ɠyu��hs"Kx���Z����M�m�@�z�o�$z���&�N9x�G�zύ�m�@�z�h��@��c� ��ԙ�z��hz�h��@��s@=�V�ls	���$�@��s@��Z^����&��ji��V
UWk�-^\�B�G;ۅ�v�0��bwl�	br��0Bn6����Z� m��@[݈�6�iP���D���[����@vl�\��k��{�X��N��@����-}V���Gs<�#�?$��9}��h޻����/�)�~�^���8�&Ӓh}�/���@}�w΀������4 �t�ĉ�ƞ&�h��@�����ɠ_z�h��`ْ	8܉4�O[8�f�Y��jRr;sָF�m���қ]�V���&�MIx�qhޔ�=V�4z�h��@/a�Zr��7�m�@���k�zS@=�V�lS	�DҒI�[�s@��[9�z P�3�U��	��E(�FY!�aH�� !�� I�����A�ă\J����D�S�H�"c�WJ��K�0�&����@�FH�(� �`�1 �0p�!��G�!�-,>�c��(e�t�#o�1��q��;�U�<,��)H�'������A	�HK���Ds�#qH���\ؐ�k�f���D�HG(��ͣ
K�Yp�/�b% ���G�#��0���JƌhG���U��N+z^�*�8�@6��j�N�v"�C[@z)�i]�����{�U��‷��4��!���bcp�-}V�}�M�m�@������(5�J3mŠ_zS@�[d�/�)�Z���lM����ٕj%^�%�u�1��<h�����1Mv�Nq>�ex�5��v���i�>��0z��hޔ�-}W�~A�Y�{~��,�Ȑӌ�m9&�}�M��hޔ�=V�4?�"D�IcO��-�M�Қ��&�}�M��Si���<MHhޔ�=V�9ԓ�s=���N!H$�A�%\*S��+�O����RI�sآNC�6��z��hޔ�-�M�Қ�y��������(��H��}��Xс{ldطz�l/*'ivv��`7.?#i�)�
DҒI��ύޔ�/�)�z��h�.e�	��6��4zS@�����ɠ_z�h���b�XD��6�4�Jh�l����oJh�İ⼙#�?$��=V�4�]�ޔ�/�)�~�^���8���rM��s@��4�Jh�l��<�2�v�"JIU"�Fɫ��+v[�tS^� H+j l H  ]�`mTcWgF:������+N�p���)Ӹ��pv��7/ný�o7[���7\�e��7b�H�7	��k�,s&�-$�kV����*��dc���Lu�Ѹ^5�n��٬��87k��9�[��r�y�ێ�:�탊���j:=ng]�^kSʩ��6N���+˦6L�@��v�]��kk]6k�c�o��˜t.�,&�����y�k�������?��}�����eW�IB��m� μ_|�M5$i�hjC@�����ɠg��Vgk�l7P�e���M"�X�4_}�����k��Jhe�ѦئD)JI&�}빠Z���Қ��&����\���a��L�-}V�}�M�m�@����o���Ӂ���5�]�pQӹ4�v;=�ܛ��r`w:�Y��n8��#y�E����n-�Қ��&�}��y��;��;������1�$��극Η �� 4k3s�5$���n�_zS@�ֽŒ9q�M�$�/��Vd��
!7������ګ \�[1<�$k��&�h��@�����ɠ_z�hz�Z�M5$i�hqŠ_zS@�[d�/�w4_U�o���\��A`��h�v�Q6:2q�g�6$�1�BgbLq���Cv;s&�ݥCp�=V�4�]���hޔ���M�L�R&��M��s@��Z��4U�M�e����LcQ��fU�΀���I*�������ɠ~+|xX��D�<M���v��>y�U`g��V�({����<�#�?$��=V�4�]������4��'��1ĜI��=v�f�m�{B	p焌��/d���t�0��nb�"M8�$'	�_z�h���/�)�֓@3��ى�y#Lj\�3J��ea{ٽ���37J�/�w4�X�jH���C@����wZM��s@��4�2ք��9�m�@-�����oJl�R�A �^� َk�RIþu�Ȅ�dr@����/�S@����^����%�͊N6�D�ײ�1j��<����)ug÷����u�vM]�d̘�n�$��_l��}�M �i4�V_(5��Ln��֓@�۹�_l����%�����z�h�w4�/���}l��?{k�Y#�!�Cc�*�b!�wx��֖w���^����;2<P��,i�Nf�}���g� ��&���@	$��{�J�UQ"�/ch�1Ɏ�IV��Yd�� )v� 6� 	 tZ��Z�:�ŧ2�gX������t]�;ms��Yj:M�Z&Y;�t}�v;����,P��
�ۀ!a8�[��:��\όbh�0�vy�8����9x��E��b���.7j6�pezv���[Wn� @���
�1���nK��j���D�G�W�T��A`�P����uv���qk��՛9n^.����p�{��*G�٭�^�z�h�w4��pέ	'<s���^������e4�)���ѦئD'#������e4�)��&�������2YD�5J��=�ޖ�O� �i4�]��/�#��D�&7�Қz�h޻���|�}�}�����$���]v���M�|���q;a�@�� ��>���6�e{8;Zz�4��$��֓@����/�S@��������D���d��/�w5D��T �֧���jI�;�MI%�h~���EBƞ&�h���}�M �r���s@;�Rjf]K�NXMQa�
"�/K �յ`_z�h���[�ZВs�0m��XwU��"�7��nmi`gݬ,����~�����2�A*��m56�a#��C��z���b;��:�$�n�Y�`L�d����z�hޔ��,�?V_.$ۀ��5�4�S@�Қz�����;ǅ�����Ne�w���ffgb�N!�~M"gY�ѩ'���jI�؉a�y24G$��[i4�]�3����DD=�^��n�ڕM9s3�!4�]�ޔ�/�)��M�ʹ�tS�7����(x�iK��%B&�u�6�����2{�9������cOs4zS@����[i4�]� �RD�ڍG�������MٽJ����Iy$��-�cn�����9�`��X�e�oJh�U���F�b�I8����3�w4zS@���y��5��:�l"�  0*� �"É�d0 ��T�T"4�o� ���ǽ3�'������&�5�4zS@��� ��h�w4��YM������q��[�l��>�h�ys�:s�����s�r�k>p�@pQ5���^}V�[i4��)�~��a�x����Zo\������h�U��g���>��Ǒbi��s&��}��k�Ϫ�z���y���6���74�5BI��k�7'5���j�RI%{��`��trL˩u)�&������a&�RQ���_����~�Ԓ�*��DU�DQ_���*�EU��EW��Q_���*��"���������"����EU�uEW�(��DUv��*�좈��"���(�����*�𢈪��(���(����(+$�k*��� &��B ��������	��>�R���        
0�"A��f��w  ��L.6���JP� e:	A�X�WN�"R�kc4ҕ� �(S	��62�(1�� 0B  ]�9�q �     A7��� ��" ɐ�i� O�j�R�  @   �L`�a4� d�@�S��R*h ��  hi� jjT�h�b`�F�0`�&�"	���$ڙ�=L���5;�O/3����DGdH{��?�*ڀ�	�����A(O�����i������F����`���Dru��� �E��"��E�5k2o�J�D8���4�Bj���                   �<��>B(��Q"*�q�q�]s��32����i���O��Zz�+u�����Eđ��))�C!�#Jb1�I&�&��h!^3�yl4\���82k&���A�$��� SUIJ�B�h�V�̵K5B���v(W+Q�Y-�`+­�YLl�aP�C��!
X咉Uu�W�i�D҉�M�C&�K�
'/�v/0�D��
.�+u@�ѱk���Ć48D? ���i �4�1L(��)�Č�$�BJ#R6�kt��W��6�=��BET�G���-@$X��Y! �X�HX°K��K�7Sy-�k�k�V�JR5pp�� 	@Ec$h�ĉ�DD�#L*$a#!B ��$H��IIA+i"Q��(�1P��@#F�SA�*誔��jƘP�HƱ
�������i�`�q����*�E@]s�M�P�.�\���kjҤ\nCʷz̲qhD��ds2�1mmOr2��Z�����Keo��kOCTyq3W1K��^�/��][�g&�j;{f6��7o�?҅�8����k�����6Q�8���^0�ڏ3�,�<<ky����                                                             �xz                                           ������餵a�l ڳm������
6�m��H���jH- -�mv�x�m�m��m��G[;Ci�9E��s�                                 ��                                                                             =�       ~���߿cm�h�k�bMhm�[Kx� ��ڶ۶�l��m��l�.�(����ڳI*�������m[IճVܐHknI��ɥ�.�k"I���j�Sv�@%�n��?�� ��$��   ��m���qm�m��m��`�4PZ�%H8�Kh�h��i�/]hd@$���M�[�<�e����^�%��6m�m��"��amp�.�L l�m�[rZ` K(�e����<mη�G���u;�IM�k��ٳnΒ����L���-��uH�]��\6�[�C�ӣm��h�۳[�{H��jYȆ.�4� .�[H�:mN����ܳ����l�sa�=]�<+պ��T�$����xЂ�n}��U_Z|�4���u�=g&P�@!�t�P�E<�-}$C�K�c1G�@ʜ��6��S`�B
�q�9� �p�2��(NT\��C���4�
r�Tr�2$��9O��|�A�!I���
؄J'�p
�� Vq߶{]xqZ������݀          l        :2[[^�Z-I���Zu      l              ���\M���N���s���n��;Uin���v��ֳ�$פ�v�v�����[-�v����t�Y׫� ˭,��*���ڢ��n> !�
��(z��<����w������ � :ݶΛ�� �S�Mĭ�M5����Ļ��Y���KI������#?~����2���_�վ�[�6���V��ӂd�l�3,�=��;�^~�"�����'+��A>�daV{����I#Mռ�W6㻮��G��2,�\��7��[��k�d &�&F�[')w<�k��.�d��:�^վ��L[ӎ	�l��̌W6�]r�ou�+v��~z�����{���[�����   :6��M�   ٤�׋��ĉ��+Lt����HK�����gW*��y]�-���jn{�r�0�}`L�`ĴD�+wﾏ���N8�<_n���5�ʋk7�&��'��ec�N	�l�6�\ݝ�k���G�g�8�'�y[��ޛ[x�}`�%�
B\���un���;oDmr��9�Ҽy�OYKq������	�d��A+vn��n��z]Ջ�޸���v��    t��l    9q�]I�	$��M����	 �p�L�Y�>~�X���Y8�]r�ou�,��w��%����r����=K��-�w�.�9�WfS���U7Y\>�R�	i�8 O��X����}[��P�ưx����
;���d@�x�j	h�`R��� �T�aE�E�� �:�|�ΪUWmg{�x!�h�G�v�E���C`��}�R�������+��{���L�mh<7��u�g��Ųf���kg3~�d~�����/��wd^�Y��%�ܴCr�+Ӷ�׽9���{�1�UO��X�?z���b�7�     �z����    ����ܶ�k;;$�sl����d	��}���vަ� 8D.q�@:�}�[�"���]^�,�l����K����yo�޿�6QRZm+�.�ou4�����I�� �+1P
��o:D񓮱�� ����A�{-f~��_}�w�����j!N��tTּ�|O�U�x�=�Dy����O�|��)=q�7��$>�M&5s����-�����H7/b#>�wZ��:�� 0s۷n78�W � 盵ǿ~��g��`���}�Fv�|g�'/돱~��ܺ�aG�[5����d &&U(�cCV^G_���������I�"'�}��Wh�~��q��~���Z�'y���~���   9��t    	�:���\�m�n�\��-3�`��DCtR�z����{���.#�x8����,w�|d����o荹��T�/y�ȵ�=>�� )	r�"j����D��߽�������ܵX���{�n(��#H��f\�_�M��v�&A�bY*w�:���L�zr�7o%���wg�ѝ9��{�{�7��ݿw]�.�&A�����l֛�~�Y���}��k�8�d׼g�wo��=:V笶w�HK �[i��oskf��kv�����l^����6��p�����?Rxm-�T����'(��B2�UCb8��HQ(e俿��~�����~                     sf�mY%��[6�җU�u�P                       )�r��u�Yt��T��$9��M��j�is8��w]yz��k����O%���K��&��^�$�e���٧n���g2N�VU��\�v�ΐ�@�ҝ�O N�v��� �= %�ɰ    �wb&�ފ��[��&��`[1��8����������U��7�u�Sؿ~���l���[Y��j���  KLkv�ǽ���}�~�K�{���-滫�YJq�Uw�n�_�HK�Cnɼ��:�z���mtם��~Ȉ����72O{c��u]��P�L��	�l ��L� Y����yjq�Uw�����͚���""���>�ͪ]W�&A�&RbA �U�S���i�m�^�Ŵ�kԽ�[{[~���S�mU*�[�    ���  ���  �v�f[;i��5�u$;���<����)p�j��0^~���N�S���{���i�ffc��˺�j|��
BX-8@3�[w^���>���u���R��n���#�ݵ5ޜ+2�w��2���� {��J��j��~��w[��}������Yt��=�{6��[���g���j!L��<��N��[�s�]=l���Y��׼�w6׾�"2q�Z�W�^��
BX ���v�k���X���{�kv�R���1�ٵj=��Z������    ��wK�   ۥD�j�Kg+�П��yݷ�B�`^۝T'���ֻ�wsk��F���������O�~YY��W�d��e�d����?�od}}}�V��b�+���xW���¯=��gWx��HK����;=�����ͨ���m�MG�my!�!�I*%0���A�����0) $�  "��CE^��O�QW�O��>��j�ISkW��i[I-I$��U����n�wѴ�%����&A�bY*`�W�Uk�zwkv���b��+��3�tB���P�/�"=��"#o�غ��ߨCm Va�{)f<;��K1�w��K��V���,
�4T6��eW�U@  [k,�`   6$��[n��[�]�c���D�����bcQ��|�ޛX�o/ΣW�s�W�(��P?`�V?I��Z���x���Ӗ�1b�}�*���	�l �Lj`��ؼ:�e�V|K�kM$?�M#
��~�^��C���>��i(v�F��Q������ɍ_
=��	  
a66�_^�Z�R�}��ۍ_b^�Ͼ���E����*ϷK^�ǅb��^����X�������c&�Tj��E�n׆����sE����yb��^���@�<x���y���«k�ׇ��Ewݑ5U�ə@
~�}j�we��_1h��O�T<f�������J�T��Z���/��{@    ��Y6    ��v
껭�n�����Zl�L�cz����X�ݴEc�cɯo�Ф�xr.��!#!H�T>��-w�Ǟ�=W�R���Y���>N�<�;��7���0r�Z=>I�}R9�V=�+�}6��z/�
s���x*���)p/^:@��|��I�'��}�r�x)
��ۅ��Mn��x��T�-\>��~�('ӜZl�s����'z�|��W�ϻ�h�Zp�������qݜZ�т�{�4Q�>��SE{;j������L�""��Z9���o�x|�0~�~ص��h�Q�}R%����Ǖ��h�=��un�=�!ڨ*������~���W��篟-�����                    ں���:�]�m��$�Y�                       �<��k��[XT���6[�ݥ�U�,�l��i�ڂ\�r��M4ʛ,�u�]��vB흶]g[g;9�]�Mg�q��s�j�YW
�w�C8�4�D���wv   :IN���   R[k�KfE��]2���~w�����)p%.�qwv�c�P�{8���h�]іC�H�l+8GV�h�r-���^���ާ��׿�����:�������ДzΩ��N��"��M�D-
;���V+0V8��-xT`�v;�d�r���?Z�������ׇSR��P�V�/EB�[F�����شt(�:�x+`�u��"�&������*��֏��Gt��l��q���kE���U�e��UP�^��_��^��qk�"�Ђ:��������Q5*��^
����/�֎ţ�t�R<�=�)�gM�Ee�7߿y�z�{��n���߿    u���   F�����X-���4�wtP��'m�c'��<�;O��}��R<��-h��%B�|C�^C�P�o�-F�
ţ�{:檩@�.��f�{��y�ry_?>�]�[I��`��X�{h
ǂ���qkG�:�.��!�¡�~��UDUL�UT(��UQkG"�и��^
�Ec��dM��kF7葶�$5�T��EC��t��@d-���t  �cl�֢���蘥���ʣS�h讏�&�x)dC��ikÑh���E���%�i%p�V2���QR�`ۆ2m8���OR��ֵ`�V8��M�GF�ݴEc�QJqʣ���q��Q�&m�    �M�Y6    hv$�v�cM���FK߮�:����l	|�:G��-���ր��ñq9d��T<�f������T�Y�#�X�Tx�~��ZldΆ7��<�;��;��ݴIm>�P���E
c�ŭ�/+�F�#�P����֎E������)p�j���{��{�{�ӿ#/�֎ţ�G���\h�Z�$�)R �T*+HNyQ"@�$�������=1;z��Xۆ��cJ�i����|+u�ͯ�܌wz��j̟�E/���AHK &a$0W�áwFY$�`�}��-xrA��x��^qc�g&�~�_E�����}�Ŧ���:�y�w�����6�\h�X�ɾ��������8�}�r/�te��R<�ھ����   �nh�    빤mm��fm�;\����6vԈ���V�E�мM�/C�Qb��赞����QvOL<�C��t��߻�'��}���R�J]t	4�s�G����8��ojt�*�vG�����K}ۅ��t-����[p�VI�����`^۝T_]�~N�;�y�u�'��M=�/��mh���U��>��*<(�P�}�Z��tx�n�&A�����?b������Z,(Z;��'���=�#�8���h��ƔЯ����e�c��ߢR�J��޻�y�w��u���'��=��=�KGb�軣,�����2���SQ�-R�_Z�]�     ��%�@   ��ҺI��t�Vr�\��ηׯE���r��M�����P��8���h��4��'釢��q^��ɴ�E�C�D�8����±�_��  
�*������)]ӔC�I�J(z+>m�������9�B��M�į$��R8��֏��xzw�O�Rᔻn�k�ާ��'���6�x-
;���W�|ں�9�g���;�e��R<!�Tv�E6�^	�v�|�����Iߓ{�3�P�[p�׸Z���ñD�=1g����&��[.���ׇ��^���"�	t���'{�g��$�_}����GGFY"�����{^��p�c=L:��P����V�E�*��� A�b0�I#��{o_����}��|�                     �,��'m�k'6t��ͬ��                       w\t��T���#4�l6���G��� �Zh�[Isk�kwl�]��-�J\�[uY˝��iWW5���O"��ݑ,�ӑ7���<��<��<���>   ֭�t    �;��m��4H�l�����)p��k1?;�𽣱G���z+
���6�x-
;����X�t���h�_�޿��D��bBT�?j����b���n*�_~y��M<]�P:���^
������-i�X�п	)�'釾��݅�����d &a2�F��F/���X�֢ǂ��{8���h�ػ�l����{ݸZ�ȴt+���*��h��Q1TK�J���o��&+�b��~�x+
���m}�y��4��6�b�Ղ_b�_Z�J��HK �2J��֏��wFY#�J4]�xZ�9��z&�����V{׼Z�����z������   [��M�   6-�3�.���L�iq�>y�O[ע�`^۝U3_>N�<�;�����6�xY���?}����X�ϋZ<��b���!计x�`곳ꨊ��D���q�Y?
5r�Q�]'���(M���5v9"�N�oGG�xv(�'鄴V+0Y��=�M�O����)p%.��{��y}���0U^�-xx/��d/*߹��h�op�;���x��x*X���Zl�G^Rz���y�~N�;oS}�𿒜��X8�w�h�xrk�����h�ǂ!|�OgŭGC�WUDUL�U
f�&"f�\h�z�c���֎L4vY⧉z*��YŭGB����b����AA��     $��&�   ���]]"��4�cmݳ	K�)u�7�}'�v Qה0p*>i7p��A���_}d5���}��-h�������{�Zl�,���|��{�����Z[J�P�Z<{I釂�q{S��^L:�u�@�_,����zĀ ��}��Q��G�9d<�G��ۅ�����ݴ$�)	!	���{��+U���'�;I|�n�:M���@�\Na/EC�mO��e��_1��Q\p
BX���MS
M�f
o��k��xt(�����B��{x���P���T�HM��T��=�C��mTET�UUB��!UU�r-����X�V@��4���h�Q�'�
ǂ��o�m|�{���y�u���   [��    i�%��kn�qRn�>�==z)�` ���ؗآ��3S񛜫Q�	o��_FY"�Ec���֎E��x��|-�E��'�j����`۔�Tb�?}=j��s&�3�.�-���uV,��o9�X)	`��@
��]�J���V��D�q���NR�yV�c6�&A�ba��]U��\�����uo������wԻ��ͷ�pL�`5��e��ou�+}��]N�0��w��^��r��=�}��    �j��6    f���^�ۢ[&����wl�Ui�`����s�s�q7�wI[��|��Y��2��H���D�{����yI��][[����w]+�w���2��6B���'=�~Xݝ�����ԺG;��$��xU�g��%�
B\� �����uo�����Ϯ���}h�w����	�l ����$��ak�򭧽�wV�mr���f��][�Ǘm�'�q���c=s�v�&0yqo׿v�                     [�~d��_[_6�,0v��1&                       e3i�]���w��%�&�m9o�u�"m���f�۶�3vMj�\Յ�����Y���m櫮"�YM�E�<v�9Z�����:�y׼���}����   ��K6    K&��m�t�&�Zv��L�`
d��b��}�]+���y���v��d ��fW�HK �[h]յ�\�GYY"ܮVU�����}�c���>��m��쉙��L�`ĲT� ���u��ز��w]G�.kR|\���k�WV��}b@ �i�����}^�����J���Ud��Łj�s����t���j�z�]�K�R�!���w�w��w�'��}�xc]��u����P{qK�!���A�A�u��(;�:��(�����9�eqQq⺂u�\ne����10�T�N������݀ 'S��p   c;K]z���MI;V��])p/\��O^wy�. ��;�7y������!qq�<޺�A�T��<D��S]c(;�:�;�������U���uwn ��ʫ�]���1X�U���7�A�A�����]L��-n�7j � ��[���"����z�A�SP[�;���#�9㩔 �1�A� �i>̋��"�f��j�D�T[I��wwn ��������3����Dt�n��1����u u7sk�w��Qq�X���]�wwEd�ws(;�8�;��B)�&��*Nݹ�e�����;�5x���eq�b3���]f�2Q��;�P{I�x��VPwu�&�bu�}��񋻻���(�jm4�6'�Imwڶ�O��W׃�W7�=�e������߀    Z�9�    "�ӛiF�L�n�l��%.vΖ�O����}{+v��u�>���[^�\][�}`�%�
Ih`���w]+>�����=�{θ���%��n�9��2��H��ư[�����FVD}��q\U�+��WX�,u1X"R�,k2�XГ=g&3.�u|u"��&��i�vB���6�{��1FN׎	�l��̌]�?G�^�x���u�n윭�ȫ��|�=k���;_X)	`��-"���~^ڼ����ͷ�Η^�wk�[��     �n],�    l]��In��^�VC�P�������7�ۻΛ�����X���������_ao-e~�6��L�`
%��-�&߽�6�ͭ�;��y{�9k�N鼼u��%�
Y-����ji�Ů�p��(����w]+�a�{)gC�Vx����	�d��Ac�']r�0A�7V�y���`v�EU�ڞ�  D��`�utwvZ�߽k���pAμ��n��`-�~�   ���M�   2KդI�-�lҥ��j	K��sn��r�sʷ���{#+������쵓o�z�d %�$�X�_uo����7~V��zn���w;�yu2�
Z�0���\��>�W϶��H��>����.���+�W��
BX�%7)�׍q��uv��>{k�{Y�{�����*W�#芇��̼�X)	`��@
�vwvR��Fk�Fw:��w���]V�&��=��|*�z�RI$�L)D����������r� }>z�\ ��Q��ԚD�}5�12e��(���B
"~Qf2	J�q@���R��$$P��)P 	b²	����>����KF�
�}��~H��
��C!�n��ξ���=���W�__�x������`�
�G�������򮡢�����4{K:��B_ ���4����������o�_���( �V����/����`y�����5�`�Ǒ���}�R�"?7��U����/��> �y�����8�����>�(������~��T_ f�ab�I�f��zTOӏ+�w(�p|}_�Q��@h�F+�� ��H�H Ȥ���� � � ��� Ȓ""H2,�H�HH�#"�Ȉ�	 ",�"�2��DGU=�M(�(���b�dq7�V5��nϤ��r||
���E(B"�$P�BE	#$P���}D7���8����A��s���y��;���9>�����?f}'!�}�QF��&���=���8�]�������������}����N��<����q�.5������D|��S^�������{c_jC�) ��
�#r�"?��~�bz&Q�T�����tGf����2��|�0`�Q��|f���? ��֎O,+�Ѡ�:9#�B���Q�@��M�b1F0��	y^!���AA��h�?�D�����������OW4���?>��6z���Җ/�r�=g�����{������`��O���zo� ���� ?��J�~����#��Xg�?���������|޽��i�Ԍr�>Oi
0@��'�����O���!��x+r���8�؈";�*U�|�؍����,>C����=��v���k\�R�J�S� �����a��C�~�/�Ȃ>����a��ho9�y��q��c�+�C�G���
W����]��BB��]�