BZh91AY&SYN�� V�߀py����������`0�=`  >=T)_ �`#� φ��UR�o@Aw�w7P�Q݇ ���{^z���sࣽkA���C����ښ��l�� (   
���1�UML�F	��i� ��A%I��@      �ER�z���h0�2�4�# h	4�)��� &�#  F#�D�0�SɣF��&�5O�jOԞF���y�	������44�hL�LFFMݶp:���0?��TD5� ThP9��� DB²��>������Q	\UPB5�~��-R��I!���t�d�+��|��ǣ��ǿ��ӆ\ֽu�SL��}2�j�ywq"$���K'���W||h�ˮ:n%Էr�_{����*ny*��\\��)�'���q��UT�Q*D�[u<��^�I*��N�i�jm�Ż<Ӊ'4�Ỗ��B�Y��'�t��w��\^)���;�u9cX�^�͵)l�fv1B���JWfUB%I�Cz�y8��:S��J��p�O�r�[:t���B�1�e��I�1�cC��9�fB8�3"�0WC� �1�1�c� c�1�6X�4c�p�Όd�>gF1�c8�4 ���9`����4�epc�c�@�1��1�b�2�1���1��Ψ��iьc
��Q�i�a�1(c$c��1���I��G�W+�UYp��a�z�o[��t���D�U�i�la�)�q�c�pc�9�j�c4�D1(dc8Θ_,��f�c1�q��[!��1�4��Q# ��c�c$���1�4���;��qC?��2�̏��?�91�x��~���=���?o��s9�	�t鸜Y3Xd6Sq��
�P�R���UR�U@Cҷ��4��e�Yd�I	1XQa�n�n{Uf�@��5a��<T�R�,Uxc��9ѳ�D�Y
�+W�6vG2B�k���Ã�o�&��D"j��7�e� �aV�,`��v�8�5�I�4�j�DN�&JL��t�ګ{k;���Y�ȱ�RL-+�+W3hS �Z$�Q@�V�-��*D{RsOx'��M�O.�TaD(�)�DT�!Q��iǛ���С
c"N���(T���y�\c9�a�F��� �.�Oʶ��f�
]��acw��>.é�k��х�T#lm�Q���gK�] ��ZFE�*���]�6�a)�1t5����4�v��sx�SetͼVb�X(t��+UT&t����dc�]J���4˦���ڳ2�����s\�Y�s<��t�rZ�o��1���X����Y�Lq�n�;��h��W��Dn.��.�ظ�SvA{K��o&*j��33"�^]����܎w���Ū&K��v!IW����BÑ���t�:Z��2|yÑ
J$�lزLGj��ǵ�,Մ��Z�+I��i�iK�I�Y,C����]����3X�mm�Mc4��v``Z�����q�ز���]+�ue��e�k�ck[I
i�i��-��.���uę�[)hW��-Vg�6�l��J��>�7�>�:�@����(�ͷv�Ո̢p�!+�(�3	��(��q��58;�m+qbj������YNьܝ���G� �u�t��:^ʕU /Rэ�����l���J�4t���X�Cq�JJ��a�K`�4�4� �c�&˳�����e�Ћ`�/�f�@�L��-�!��+akף	��m�:Q�K�� S�5J��j�jhn#l��J�\l$cŻ8�C�H��"a���!�b����(�]a��f�Z/M&\lkv�����m[iX�d˫s���Zpš5p@ ��+%4��6��K&�LJ�m�%p���T:��j!��^)M�	f&��RU΀ߞ͚�Y�g�P���V,ɼ2����9��.n<#K�'3��m:
�PB�B�PB���P�� <�$�&FP"D�����,IbJK)cIbJ���3&D!�)���x��>�1�Gf��l#����:ٖ�lZU�l�-iT�e�kJ�k-�T/("ybD�,H�*C�.�m�K�p�q�&p��l%�n��6�;M��Ѹu�F��7���6�;F�����Gf��m�v�a��m���l%^�kʿ��f��J��(��xЀ�БU9	�� q�
��&� #��rX����}?�z/�^u����ձ�<bNU(%R�$+D~�/em�(q�g�о�����Y t$G�À��0ʪ�9cl$QE�U��\�㏆��p�(��Q�k��b
�hŖ�9K�eX�ł��-(�X4ؚJ�%�1Yar��m[�M��Q�1	B3 �� ���#Zi�K��Zo�4�6��Bކh���r6��t�*�~� /�𞋅�gF�z ˤ�*�*��b�ǭ��aj ����7�'V�����9ΈgN�Ӣ�fg��%c������g���N���gS/4�CSHAQJ�wK.��0�^#��$2�$�QӤ.���ёF������ǜ6�,�2C�v:zC�y�a�|I(@�1!i�SJ���)��{��;��!hg.w��#�\ �h�ջ�,�\�q�� }��U8��t���{�B�!ͱ��	p�l�!�C��:3�[<�
ΘCH��cN���sm!%�|s�w�w���q�}�Q"�""D�|m��)�P�1��������Hp�X��# �DP��nzΪn~�˺�[���9�<�D_�DB\�����I�!׋��1,\9�e &$��q��Ѥ?NSO�#��E��|9��#���<���
#:t:0��餶J����z��5#��Tt��>��F1�� �jV�@ӓ�<� D2�'�d]}:2�e�v�G���%����υh��>B�x��G��T�� ��3䍍A�
:D�+�@�-G�7�E�9�}�8�{71�_�)�Z�2�0(eY��<?�*d�.�tf��x.����I��~ V����#��w{��K�G �#(�������v��a� Ϡ��E�$�=���$�82-����z�!�P֌��;4��yIv#�!�GVao�Ae�(�1��1o
�z�GY/�re@��cG���B8��0���9!C�\E������;���-kF��]��]�N���@W�� 8��$AAd��bt����vLkRٶI*��.�Ud|�sϷ�SUG^Cl��i�Ɛ�Ɔ�h%������i�����6�l�	k�Gpu��0���b�x�r�SIaX�e �	P�4yE�4�����L�ᅦ	����C��j*�*�*����������TUb��������������;HI���;����;����D%đ����h0c��?����o;$��]:J����"!U���
�7^�Z�u��2�H����4a����'�>�l�<����_��^�$��/ǋ ��ƅ:A��z��� [�?�˳�Va_:>���kx:�9;�B�g��ξ���6h�X�A�b,�	$�K��	}W|>���tiQ����J���G";ޒ���tf!}��_G����\$挵-=��׭y�6oЮ�;�$�?�|��͢�Ic�b���e��$��Kg�O��}W�p�8S3���RA�a\>�QC[æ�߲k<O�������:D3�� 22N�Jᆌ����z9ҭrv2i+� ZA�vq���EɄ�8A��O��^�����5�#���4��4AQ8|��1@1�*��s79� E
X���;���"�\Ƕ�-�|���Z�{~��A��Oh�����	NJLgGD�� ���'��{�)N>DaC>Q�Bdt��2����b^&@��%exb�\	�!�̔�X`ag��F� ׆��|��D�4�WE)�RB���#�]{�Y�jyRQ�'��!$��$$�i��r9����F��a�c<Z��3�]io�߀�*� �]��1�s9��@τ�#F3K����(���H��!��	��p����,ac.�a�R:�Y6lB=VrHs�2d����}�� �Ðw� �p��|�4�3��j���sh0߆�hC6��ɜ<k�Tr>Y�: �pk�bG}��_d_D>�a�(����A��I��:dۑpx�#%�t��""��"�5�m�b��{���sm"Ǟ��W���\X��eFʬPQja�r߫�_3�trh�����4c��i�%Db*�s��QJ:� [�:���b`qa	y�iV�-�馌��[y� ��1�+ńHiBj�$#�q����@@�`Py��J@H��d�B""	K�,\HBa�S�h*��Ӛ���m��A�`�!�A���	��o�9a�x���×���4Ha���HJ�u���-��pd�%��l��C��h�7À(b.��aD�����2�|)4	#��$��KH���M�F&C�@�|��Q�~�$�3��J'ṗ"\Zje,��v.����pF�Y�7�G�lLG��]��c��1��83�, w�z�	���h3OH�(�<fH��B��ԑv	�x>�S8x�Λ�cӝ��!�U3�icLrE�"MU��[�4�C�IĆ,J�2�g+0��z0����#�#5m������ů5��<t>�ΈA�obga�ƖO���I�Qbֵ�j(ӍfkZֲ�eU.�f4��u�;�z�[w�n3{c|���_*�F���� '��cC��[6`��w��M�� �!lƛ`�Zoע ��eQ6�T�01������f˃�3��l���s,�1��3Fp��F�ã���^yǉ"�!�I�D,�9��5ʆ���>E� Y�%��nI� 3���t����Y���ҺP���7�F)Y�'�8Uˬ�;��8�L �X3���9!�͝ ���<g��f&Np�GJK7�yw� ��� �nj�A(���:��Ӆ��:�~�-I������f�$��F3���	��Uwe�s̑��F^���
.w!��Ä�$%�f��m��tv/��%8O)U�E� <�[��#����H	�:����E�&
��8�T��1���7C>/�]}ڎ�y/��e߈bl͕��"�Pm(i�T�e)�Ԓ0���8�`�1�,�F$�
���Ckh�cY�f���v`@�]�	5���`%��I�g�R�d����w�熜 �c$�6I#d"�%��p��*�#����͂�#M�S���?G�	fä�>p�cgII;�$��ꍳ���P���B�"	�Q��ay�W$��iQ��LU��~=��;���L*�N���xh�0�uN�7���� ����Y�᭕��VjLf(=D����.����̊�1�$�S��$�W9���8i�\������Δ�1�g̚X4Gϐ�4fhU�9O���� ���2��kn��J$�%Q ��m0F""�BV���؁�m6����"�gןvn9��Љ�|���]H��G ]/a��O�_�(�#����9�
<{8��Y��0������`b�AD2�F�"�P���PYPۣث�O0t��� �S�����E��$�7�tB����{<���wFΌ��b�ث���������.��H��<0�Vo�,�*��JsL�쌲�S�Y]�5e�{Ҹ�#��"E���^Ά�æ�c8I��/LI$>�!a��ܥ�ux�~XS�ć��/��zx$ڲ���Y��fo�Mʹ���]%TZ�(���j�햚���F�@﯀x*ZLH�R@P�.;�t�0�$f�U�dӦ,�t�\�ջ���
c�yΆh��˖�,Ġ�m.f�#�q.J��j9���RR��I�X2P $H� �Rl@�@;v�i4�ȑ�P�;I 9�@#+֮ �2��P�"�a�k��=�>-�L4�s�ą.w���'���<o$����A}̠:1�t�|7b�c�a|��p$����\5T`�X1�W�di��	������Y�^�e� �{$��܊%@��lr(�,��3���$ZHՌ�.���
�E�p�:0�I�|��a�0$�A�z�f}��,��zvJ�{B{��+=%�\���"��x�g���KJ�)�{ьD4 ����#��V�bgJÓJ0Һ�dA�]��0<���7���(��ev�D6|I�DA̐� ���yE����_V��`��lo놛�/�mKq1�I�����>I����
�
��RJї�0VE��nTz�+����􎀛q�J7��ᇌ�����De)"�*�NAc�S��:Y����
�te�\��`���<Eki�m �BreY�e43J�!;�*��bA�C�v�h��0xϗ�N^0�Jh���^M�2����o��L�6Hv0a�L&��%_��G2K0���Y�N�=eo�8��Gyl�W��Wq0䐩 YFBTan!��A%@������4,��|t��F�,3����(e�S׬�b��oǈ؉(�I"*��f{�R�Q�/8<f����������r#�8wG&���+Q�� Y�s���z�DQ��J������J{�\?����J���E.�'�eA���sR���[G$���<�JP�4��˄i��P�La
0�H�(¤�P�E��0JȢ0X1%)`��d�d��R�]e$��$Hr���,�m�:d%IC��F�@$�pE�AD+�� �A��BATj�Y[��PG�
 �� ��o( � M�Bk���	�1��M	�j�
&%�p� �����T�V���Uq `�P�A�2����mO+�:������p��THȊH(

l���e&�{���2զ��"?h*0@O� �*�T?Ȁ� 'Jo�
u�G���VE������`T1T?�E���q�Ш~@�M��[��E�b\@M>:�n��P� ����m�d$��BI	$$��������*����*���ATUEQTUFH*�Bx��ǹ8��پ�T ��W?F������G���O��� ��E���:�7���������9 ��_��������G�S���E�<�>�JUA	��@���m=2��CӴ7�+�K�Q�@P��`'� ��?�u����)�=�ʨ!��!�Q��9����-����	㲆���﷎�K`ZlHd���D�Y=���wR��Ƴ~�Z�D_���x|�U��� ^4����昞��yb_%JVAm_, K�@�	 (E"
��@ �D"�QiTH�"ET�! XT� AH  ��i4�>�P���	���0��a�=���,�P, ,�2(ȣ"��2 ��bc��s15wk~��!������#3\@.�����G�����	����� B�b�:�^�K�-]��z�Gz�_��l�A��:����0��%�>��Hk=�!�� ��ܶ׆}ZjwB�k�'(��� �P��I���r{�*�w�xk�{!�;M��P�<`��];PC�=�}'�CS�Hxc���j)"��w�{,
"��5�HB&AhHQ��0bd]5��q��	݇����
4��? [S�D�h" �J�@��S!4[�J����.��i�N��Oi� �V�vx��f�3��q�t���w����9�EE���y��:������7w���ζ@�9�_?���=$�='��=>�N���!_}�6�n��'pq	ت���F(".&����3�ޛXu�0ܼ�P��[�)hh1Vx��Q|��!*V��9λo�ę�M~̹���e���hn�&ˋ�~}A��@ײt
�!�5�C�mh�C	��s�7A�s;L]۴l�@ٟDD� I�-�J�l	��1�)���ɶ	D_�{˝�mÝXl� ����C4�w�����V���ۆ���n9C4��J�!ޕJ�1Gų��v��rE8P�N��