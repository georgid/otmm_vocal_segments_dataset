BZh91AY&SY����R߀pp���g� ����av?DJB(�E*� HUEPU )@""�@�D	R)(Q.  =J�E*  
�AE!%"B
��B�@QB  ���(����$�P�� �**p   ! �	 *� X ;�2k��ƺr�r�� p����`��h�U�A�G��ER����AW3��=�������&�h9�t�hWm�@�R���fj�3��h���{j*�E(8�B  (�P .`�9�T��C槟uל��jvq�]n N��>�n
Y{�j9�w��o=ã��� ���Nw_-m\M{Ҕ.疇��@�����R�r�T�u�'vڷ;�U�>�_Z�����>ʹ����ͩr�}�Px>��P� �B��Q�� }*g������w�kͯ��v9�< ������ݩs�u�Ǎ�5\FU� �3�ӈ�zE���t��W8}��ϡ�>���Qg�w���;� �>'���|;.}�S�����P@   ( � ���> d3�ɪ��8��P7I3<�8渘�M� �bdX���Pr���� }�/w>y��N)�c� �b��r7ͧ!�k��>9P@  
�Gu� ��2ԆL�ˌ�x� �F3T���3�b���S�  �qw�^ F:��8��&�[�Ó�@}8=2iF�{��gĸzP     P�z�M��R� ɠ    �HIIJf�zL� 4d��'�UJ�z�       "{J��J% �    "���E6�R�@h�   
DJH���)�C���di���������������_����}����"����EUt�**��U�� AWI�����`�"���傂*�w�R��AUw���hEU���5��5���i�Lј%�T	��12�ԦBPhsO�SF�7�ۣ[�����d"��O-I��6Ì���Aw�:U��*�����FE��y˚qϺDi�ggtO���%ɧ�O$
GsJ2�y�
�VE�IC�g~�u[�-7
���Y������d�f�=H֯���p'�D��X7��F�@�.]K���\�z��m��н��99�%&&BP`�%	BPd�	�`�����\��2��%ޡoN���ô���V��3�y�b�E��#�g3�5s�=�T=8�8p�w<��ۧ�.2%F�8#���g������'q�P�R�8P�������K�J=9Ð��HOK���f�xy@�e�
6=��(JLK�h49'���XÐ��Qփ�;&�7
���i�o��9QpX��K=߾[;�ew;�=�o���rs�����j}�8�������/��[�s��>9��ui�ș3ٻü�/�r�|*�5rvLo1��:1><�Bd�Q�$��((r]�Bf�O!(O!7t�����d��O��y�,#3�5NG�D2j�}{�����.ç�Z�<��R㖢��pխtugGFu�n&��Td&�K���H�ɏCz��͝F�|��_{u����uo;��!�I5	�M�Wc�O��,�e�tJU8�������{��Y;O�c�;�/�9���k	�>\�{�>����i�um�uh�j@�Ib߯Ig�Nwv4/���p��}^|�;����~(����,�{ߙ��c%�T�i�#��8�M9���V��#g����ь:������>ぢ����=,:�Uu�����4�Z;��k����J�J3�=��(06jĨ�y}׻�!�v�Db5��>w�Ɗ��Ө05j�3�ؖ.�-th3f^`xe�`��ך�8Ld%9m��ѝ�#�{q>5	��P�%��u�BƱ��ߥ��k}�i^J4��-��#��ܗ"_d�9)���w�N�ϵ"�F$�P��{�G�"�D�7x}/��zo�i��:{��c�M��}�L�.�xwO����a&��!wpJ�g
F����[���l�̝}A����g3�:$����(��Q	�l�l2��CP��'Z�����0k�ԍN.tvBP�%�%��QF��kHԆBVL���:� �=>c��f�Ox�&��G��R9ޱ��^��(N��7	Bw	BP�%	���������d�E�y�z��Ϙʄ��q�:�A�Q!�a.���]�����$���Ρ��p���s��9�d�X�*�N�ӏ��¬�t��@��}<��\7�>��[e}C������V�>�0K�}!̓����
�v]��p5����{���;N�F��sn=Fh�ȳ^zh:�{��V1�[ӵ���e�g�� ����s0��Mו��7g�O�6�ӏ
��缻zs���t��7�!,�F��ƄPzz�r��J��5!�Hf@aL�JP�t�u'Ldl06���ܧ)r@�Ƭ����8=)�d�G4l�rK���!D7l���D1r:^q2q󎉊��:6��v��Щ%���V�:�W������Z�����9k�澊Щ%�29Jj�e�|�l�2ȇ�rrq��4l�V��Y�}	�N�7!(2�f�4;��'S��22]��z�0H�,�iMYx�����M7{*Uө�Ó�F	$a�b�<������u�W���PŇ����$N�;Hw���6%�縹�:���	!�7y��m�o7��H<J�W4�sV�r# j�w�.���b���yHϺŐu�MBj4�偤�'J{.��F��C]�{�+V�P�@����*�+��i:>��Ic�L_�r����§����8]���BxӇR�C�w�w��:�N*���_��ڽ�cH꙽�M�����{l�Va�OQ���2N��=�Ѽ��t��v/�5�z����>uaBn�5��:z>z:�5������F����EQD� s4ޓ�[�����q�Â�LӋ	���;�w3�e}�h<e�k����M8���to�;�,�iΌ��{��:���ʦS��;�Ŏ���u^��߽j&bF	 ��������� �q	c�y��l$"�S���D������v3���sz^���}�xԳ';�������8��97h�[�\GsI�-Xh��]8G�������V�|�zrNubʁ�ox��K�oM��,{�#*3}ӨO��7�,8����#�����FB}	�'z�:��(N�(J#���Js�;��W���_z��j��b��Ny^{�x�xNJ��	��gSB��O
��;Ǝø��6#��;�h0��:�	�y�Y
q����;���Y9���e��8�q�a�oK��Y�dnOL�0�g��g1}�4��3�3�8gS�u	�tGQ���z�N�FF��@ı�(��>k���ݜ�Z&;��"&ע{w7;�9������o�Lŋ$k��*�f�'{�L�,P᧺�=��������t�e\�u�R[�{���<�Of���/{ީ����p��͑B�s�7r�M4פ�ά��G^�wg����N>�v��P�Ç�{�Qެ8Av� � ����!����>@��Us{�ߺ�x��Vt����v����7RHS��m��� ���J\s2'0:;�v�#7㩒��)J��37�4��⫝7ͫ������>��d���z�K����3�!�	���>���{ҳSWO�˾�C�ȀcPtO�(����XB2�;���?���︖��N�Py.��p�GWe8XĦ�C�"�jϻ�.x":_s�Ϸ�A�s�1}����V�Ż��5��=�$Q������js����z�=�����rs���� �ȳ0K1ݴ���qѰ���rk�C�j0�+D᣼�����(JR��J��>��L����.l���f�V����\��w"AJlX�T�|"�8t�Y3�i8!jԃ��nr�N�q��	$�B��.wC��-��1�.9`A{�.���Oa(KI���پ���7�>�M	����8�&��D��4cq�@����`����K7�2ѹ3Y�[C!)�l���`���d�Y�RdYi5dĄDcHn��YI�� ��%.:��%i�)��a������t}�f��������~�hI��<!�N��u��'Jv�;��ܹ0g�9��\Y	�(X������uFw{yu9�t��{��������~�{*��Q�9v_o�y޳�W+/gN��*=�,������D+i�N��Y��y2^�k��{�{�m*���-��8!��T�B	C5�g�iï\�]~t_o��h��i�D��/*P�2��{x'~��22|F	]�\Pg�{�������>]g���;9�u�T��]_s�}��g:�!bD�Ա$'��vzk4�N���`񨞏)�RgD�Ͱ�k����5sy<��}������.}m:R.��iĘ����!+=�aB�!�r�k�L���=4gqU�&z��Yh��O����R�:#�d���'���n�BEC�y��U(y�S�Yha��f]~�L&��I�yLW�%����2
Q�{Ι�P�Q�qub�%�9�O_b9�m4��X'��̝dԸtV���9��v��Ώ,�'�y���mEM�����}b����bD��<i��`�`���Z�Db�lA��&}�~*���U�Ø���t����Q,;�BP�y�r6`2��'К��M�� �Pc����:�D�a�J��%	��%	B���1�=��'4�vf�
�"b_W���m�p����HUOs�P���w��%�ݝ|����.�:��$I�9�L�:�p���睊v:,�!�$�Ϧ�3���]���ӹ�ŉu��yo3�/'��U���<�|����w	�n0�H�Z�N�{�u`ϰ`G^z}9��&���#������φ��i�QVT�������x�o�6��$��~�u����=,ğ.�/#������)�BC6�f���L��f11`/����.>`��1��-�%4K����a0PFG]�ܻub��2q��]����,۴�=�y{����%��'W�K��S�7���MB}�bu��JC2�x�Y9>GR�bk ��Zt�J�N��w�>�����!���g}|������n!ɺ��w�nRw}{����8���ُvΏK^ua٩q��L�'j1�*�5�jĚ��b�Z������'w��A{��go��b@�x�[��4�)gJ}�L�#���Bs:(��c�7�Ø!�nq���"�אZ�79J���/�j0�a�e�y.}�$�{�^f!<����!<��p�}�P�&Bn��wtώ|�|z���Q�z���tB�a�с�e�.g�9:t�h��8�SCV��μ�s���qfd.�*�@[2�4�8$�t��Xq#:\��)t�e�knj��l��ܸ�2�����:O7��0�:�����I�&SD�Y�a�Ѭ�h�0J�`&BP�`��$�A�bD:"��u�M��@�U��C!�3 )��JrL�&�r7ր��c�3�yj��$w!��$!����X5�&6��ޖk8�J��!ќ�g	�ds������OD�(Q&K7WO�CM���}�}�&��d�����y<sN�!o,�g������]R��v#xɝ�{�r��:C!vnwy��[�����ro���z��gH��9;Fw��<sjI�|F�Ve�(�!(J�di��^�a�w�e���A,U��/G��7��x���������S"ԙ,�\�AB{+�q���%���'E��w�������]l�1#PR/.+��_J�',ٮ��]�޶w����@�<���D4Ѳ�A��]F�o3
s,��PhtS��a��34��`��l�g�������o�g�����ݶ�h�                	 p  -��         �  �  ��      8                   �$                    �8��˦ʹ�Im@R���n��n7$��$6ؐ����km�@�� l�M�V�-ɰ[[m������j��UW]6^�K9�Ζ�sL�l n2RT���l�R�c<�W@U ��UQ��ko`[PslH[4�:2@�R���Ơ9��*UU m��'�9����6�u����`  �  5�0-�� �@ ڳ-*�UR��i����P� n�^�@���dQ�.�i�����l۵ջUpR�J�Gp�TQ[P�1��^�׋�5�  � �n����FڻD����ٮR�Ie� S��vh
���VɎ7
ul�R�mWYF��Vy�����Mk :mqmm�۰  �I�     ( ��                     ��p   �h 	      ��                ���     �  p��a���e3E�H    A�     -�@ � �m�   �    l  	e��`�7� �u�$ �`.Ҭ�.��#e띶;se�)˻Vi�A3l�c��qC�(�+�Bb���n���F���jK[b������RtݛUYF���fLN���UQ�9j����(���q*ލ��UN� h��y�Ö]�d��2*�KUV��Om�k���̝/mu�Kz�Իmmm�5����۾ޜ���1ڊP���Ilv���N{�:�:�zC��z�'��Þ���=�C��ۦ�Hդ�	77$�iV���T�j�V4R�pR�媭�y M���p�5*�VQ���z����c���� ����[�|��۶�lT���ӗ
zt�`�C\��N�l0�0,��p؇n +9�n�U�CX�WA*�b��ڪT-�9��;U�Wl,6�:L� C��d��.��*��f�VY�[P*���E��Α;k��v ��p�l�6Zl��͵i9��4�/D�ݖ�4��  ���m@U\� <ڝ�h��Ӱ�ջA�U;s�;�j���n̪�O'@v���'�*nݕ]�%ݻV;�[��r���C#p�m[�2�T:6�0gx�B�.{Ӭpu��YU%�q�o[jKg�� �'D����6#[۠��t��d趁�l9z^�M��;&�۶6�;�WU×��`   [@Yצ�i"� �V"0�����\��нq��l� M�  
��ɑ
�@UV����Ky�A,�=�����[t�[H5�u�%��A�N�� ̸^l��Up�Bx.�e��3uW:�{EU+�[��5U@J�6Z8pbDr	�v���#�,�IsZ� �]z�_���zA�ě�,�t�e֢��v� :�-�8�K{&6�,r��bɽ6�`��+ڮ�tZ�?�G��ݶ{A#�$:%�֛+�N�ú�v�8���(�@VjU�:��f�s4��Q(��fU[b��ז�rI�[x-��t����^-t��[H{(�꽵u�	�� z��˱��]�^��S������J��jÀe�`�^@A!"ɓ��H ��J�ղJ�Nٵ�mmp��Z�����W`2EYd����ȝ��U/3U��[*�s�A���Ɨ��gU�q8Ii�M�����eٵl$���j�i����d�r�t�̑�l  �t��m[m�YC�ٷi;snٵ�m�"� f�����0�G^�k�@O�}�H8"�`L60ʄҎ��zP�m��t���Lkl�   / �e�ԐX�i-�� �
�SX��sggE\pLX�W(lUt�	d���j�J�UR�ʪ�/n�@�l��n�m��m���UT9�����yY���h	�� ��ѭ���Jt�UmH% =V��     ���H��r��v� �  X���HSe6YV(�M��6�c�Α5 �
^��`	zv�"^6[v�rK��mP K5U���A~_���-ϴa-�ԔU@UU[R m�v�����?N�.� ��:�RKh�l���9�M��j 7Wpm�` UKh����$�5��-�Rg$�]��
H7b�m'@*@M���s��M�79�0I���UC,0�Ar��Q�ȫu�)�����BD�5���j:�%4�<6�mqm��vYCg��|(�8���Z������q�0�*�Sg�n���Mv�R�K���J�V� � ��L�ۍ�����7:A�X��*m�I��X�N�6���ltI:*��e�^v9����Q�UnҒ{5j��wg.�����'��e�8#�mD�ziYTf��T:/RIms�ΐ8d-#UU*:�<�
�r�vQ��+�j�s��b��PY�m�ض�rT��A�l��� ��k��,\ �6���`'@m�E��m�m���@,k�m��h��6ͺI0m�`�  �]�˴�c]���fh��Y��F I#���q�2 � 8  Mmvε��-�l6�Ge�r�۶   ��:Fm&�,� � �%��-��X�Si�m�pm�  �ۈp�Z�x  ջs�K(�$�M��  �[d�,�� ��` M�[@   ڶ�a&�(p 6�۳m��kR�GY��"�m ^��[% m^�)���l �u��Z�luKu����^B*�HJ���� l�H2��k�oP�( d �Z���� �` ���vv%��j4+*�utH��68$$  	���H�mmm� ��Kz�
�ʵIST��R� ����d&�@��֪�<�m!� ���۴�t�:�(5�0I�&ճlm��m�� �l*ޠ      �%[I6� [�tn<�z�i�nr�mZ� 	;m6�k[l8 ,��[i1m$��UWj���\K .Sk��0 ��-6q��-� m� g]���[v ��mmM�  ���2V�l���^HI��I 6���ZM���m7k���	#N\ [@ v��`[@ � �[Yi� 5�&�UV쬭Uj��I  �zӃ�k-��E���G$��ɴ�Y&��I�`���V��T��#H�uiI��ﾯ�$�ێq�� Gi�aj�U�r�Bm�grĨ)���2nT
�,����-īugF��]2*@r��_���g�疠*�u(��C� *�(CG��:f�:j�.ɢ��r�x;5����dd���f�:�
�����zڏ����>�5
����m�ԯf�}����8�W4\�HH㝜I=T���msm�i08:��Ӱ��N�ˇ<�mi5����[hʵ=�vZ��T���SO%�Gd�vں���m$��7)�:ꭂ���BnvѤ�{�ݐ�E�P� 
|��VG�W��M��mk�7GY�i;�n �8ՠ�U� h�7SJܪ��Pp
��]WT��]m:C����xY*�l5U]t���g��Ce���d �!��j��,�Hy旙Z\5�Hm�6Z�mݤ�g �5�Kz��¬��ml�UR��"nY�#������I�t.U�+i���;EJvk5�]� �X�����y�DN���T��x������R�.�	���T�i���рv�m���^*�l�u�]��.�N�R��64�����^�Ǜ�6���ms�x��tHlc 		�-{d��GK(�m�MGh��ywj�E�f����g�;,`����V�����Q��q7S��[���R��ω�P    �����m�:.��Y$svmٴ�l����Ųk� ��   p��u�6��*�l��T�ĵM��6��e��^�m�m� � $��l��AN�M`���<D`�i��H���I� nۗ��[d4�t��H��J����+�`^x�ix����t�p�\=��W=r�D<�fOga���$�ۇvE�����tgv��m�˅�v��vv=;u��98vc!n�aw��V���k�u�읝vX����l��{b뫛���Hz��D������v�Ҷ [���u����[���    �m�9��l���;�)F�U7+a [:P  mB@ �����r�ڶ H	  �~�~��b^�b��#QX�m����Km �[n Pƅ��յ�ݻ �/0N���[t�E^�<hn�7h-�,�T�]*��@v�ڪ��骓"V��Ge[��j��n9F�:�c`�
d�C	�x]\�2L���ݺWo)�Py�׫�y�Ht,v:���Č���im���q4���N����x�u�9k�Z��77(
�ggKm[���Pl�m�    8[\ o{�������E�����?�US� ���~C���U��t�h��?���A�h�W�;\�E�G�:A;^�O존@��ҏ�)�C@)��C�AKQL�U10��DS�R�5TMA0LT��DL�LAD�&�>G�� P��L�)(�z � ���� ����!�j$�"H	*a�	��� ��	(X(&�d���(
H2dR�()FH��i
d�VIF%�dUv�>���OҀ�|"�B�"hD��Z X�|U =mN�]���S�~<A\@}DGH��C#$���Q<�

/��"� �U�P{0Dp::����EP6��
��h�A=t*�>��,@�S0Ȳ��D��E(�$�*D"D�@ Q�0�LT�Q�_@� �ЩHx�|�	�_�f�_Ed �@�'���$q@�6>����YN�Y)��B!W~��"= ����*&�v�� �}��EU���?��������tpO�
��QD� ��JP!P)REiUh(����Dz{��Ο��5m�  !���[@[A!�   �`  
��ha��9y�f�n;nWi���94gH�X�Ƕh�Y�G n���[Eu]H!A#i�:ẛ��ĖD�.����U�.]�m��"��� 8�b��hl   �mm�$�8� %+�� FN�N�hܖ�l��sZmg7��Y�@�����d�ڥ�7m�5�C;:ݹ���:�ma+�ݔ�Fw:�.�s�8�zprn�#v�A�mlkbwn��b�oh���an޶<v��p7jw�V���m�0�8�&�GIq�	:i[{mJ|hwbݦ�]�*W�]��1�B�l<�n:`ݫ]WmBbz�Л�z5����M��8D��U���j�:y��r��.R��2�m��q��̮��!�6���=���)w��M�I35$J�Gb�72�ɂ�:���lhW<�u�	���ݚ,/ ۤ����\�:B�)��;OS������a9b��^q���U����
C���m�5۸ڔ�iCo�<�HS�n�4R��ݦMLHn<ڠ���gl�����NpX�2�;s��qv��-���6c���=@U[ ��d�(ֶ�bq!<i���c��R�U��ݳ6��R�N��nv�6����m��3�v�!f�7ְݻ%�`֝�'n[1�UUŎٺ0�w�U��[@�4��m�ֆ�Y-u�*�T�b[�YZݩbF���lP�7Z����hE��Q�6�ω� �$�[��7gLV��֝�N0�㩺��K`� e�>ZS�<u��t=�l!��w�;�&�K�L����]��9���ZqN��m�:x�.'//.b��uv�4{,���ʤq�Yms<����	+���k��\�P��@��tm ���M��ns�N�긞w�<�Y�u�V��n��saii�e���9D-��xU	UM�L��w`��wa-p�gY�n�y��Oc���|��<eͯs�nt�tH��0~w������ht���=
�c���I�+�'j��J=s\�y�-�PpYc;H����ԝz{�\tlV^��Sn�".*ڷf	:!{rnx��؟�8�g=k��ۇ����Gc=�s%o��ݶv�ۜ69v|Vխ�t;��5÷N��,\ݤ�E�M �5�&X�����;;.�4�ۭ�K�e.:m��.�7]�v���m��+vN�aH�� ���C���]�lg���/_����ǽ�O��9�8rv{<dö]�
�/d8pe^y8�p�r1���e�^��`�y07�?�w< �(��ST;�Wn�I����x��� }�s�>���_{���C��i�m�{���� �˺�ﻞ�㹦�+aM	5Wm���� �˺���<�s� �����.ؗ��ջM�yw^ }��}�|`��x�#�~��p����j�y���8�Co\r�S���t�:�i[c��M�v�B�i� }��}�|`��x�]׀z����wbR*��K��|�� 1�$����� ��� <�����i�TM�ݫ�N�Y��� ��V�R0����!Z�t���N�x�]׀{��{���� wr�St;�E���� ��� ����������.�����K�mv�ՖB4��������4�+�����[=���M������۴�&��ό ��� �˺��w< ���M�V����� ��� �˺��w<�s� ����4��Ve��Yn�����RK��뫸|W��o� ��� �λ=�t��'��U	�ٚ#ڕX�H���Vޝ��:����j�*�jݦ��>�>0�w<�.�������Yj�Ҷ���5��]�wtǷ����QnM���u�s�\x�U��)�[@�L�֘S�� ��� �˺��w<�.��>�/st�j�ҫ�e;M�yw^ }��}�|`��x�
9_~n�t�`�n��wU����X��� ��V��}�&��hV�m�v�xܻ� =��{�ﳪ�Ђ�"ZTw�~��U���Rhbh�I�������yw^ }�� >��w"�~
�]ۻ`�� ��J��+��Wۮ�:�T�җM�J��V�&�+���ջM��� ��� >�����Y�g��;bꝷx�w< ��� {�� �y�z���Ŧ�@�իv�o 7������>0��< �{ԩX���豦��w<}�� }���s�6����WcAul��������J�}���ݫ|�Ƒ�QAa�D����};�N��,�i�p���`�+��+�lU�R "���p�׫R2��t��8u�&��6{>���<�M��8���d�ǭj�=[��fX��{v9�<�&7�3ۍ^�-G��:v6��JC���q���$lj�i)n�mN�\�4��8���;��C�so6}u!��X�,=�]�\;�҈��S�y-�r���7Y�V�{����n���Pw�v��ݴ�S҄ںEMӮ���ճ;���~����1vZ
V���2�RI��#�}�x�w<{ό�_z�6��Wn���i7���������wH��8`����Ԛڱڴ�j�x�w<{ό ��� {�s�>���M0WWt�j�ݦ��ό ��� w���s�>��g��;bꭦ`�����< ����y�}�8�J�[��Ć�r$Sn7az��F�z��VR,�\�:�䶵�{s�Xj]�Qa��lw���s�;�>0��x��R��>*�v��-Ԓ����#X�F&���k*��332I�b����
����be&Z�4�)�.�5�~� }�� ;�s�>�.���H�ҫ�e7�w�|`��x�{� {���\�w���`��`��x�{� {��w���_z�6�h�`���6���< ��� �s� >�s�7��Ppݫl@�%j���n�8�wQN7eun���yLL�9�]��Zu�3�D��+Bn�o =�s�;�����x��xߺ�M:WV]0l�v��;�����x��x��� ��]��:T��m3 >���{��+��QE*��3ޑ�}0U�~��m UjջI����}���>0ﻞ pwR�b��"��-�o >����|`�w< �w<߾�U�]�6�m�]Q&��lm{h��J!�Ǚk^r�����2�m#rFRu
�u%���-I.���{�����#�	�U?7@�[�f }�s��s���x{����_6�Z.�$�m� �w< ���w��}�����N���ݫClI� ���w��}��>�߁��}�ԗ��9eCeJ�:庑��� }�s��s���x�,��#����Z98Ҽq�#yU�����[��w\���r5�C���fu͋7u6�ﻞ w�� }�s�;���=W��SI���%m$���s���x{���� 8;�"�WSV��7�}���>0ﻞ w�����֑GR�B��K�f?�~��RKޑ�{��J�����x TJ���;�&	6� �����}���>0���5v�����m�c��ҥn����7q����h�������g��'QŻZ�znۙ�q��`���wlNc)ͨN݋�������c��ZӠ%��jt��nx.V��R�N;k��!��;Vq���:mԬ툆���A�r`J�)>}k�Wc���O�X�<)��� uFYK5#���u��8�-��:�G<��l�ש.t�I��	в/EKz9t�ۛpO{������;G}���8�Apd�vN�]rNVN�D��DnN:m�WmB�E���k���ڡ4$�M��7�x��x{���� <}��;-ڴ6ě���_3��@�R,۪�}�VG�u������V4���� }�s��s��s�>��W�v�2�`�Si���� N����x{�����i60T�$�m�����ozM��C�}����/�$�&'t���ݶ!9톫�$�f��VN�rmy��;%9gJpKslܩ�RǎT�r�����>������s�}��;����8:�Lu%e���|�L0������}s�w�=�G�e�c�T����~�۝��w�������9���]N	؜��[�߾��>����|����i��{�)+V�\q[c��>����|����nwﾹ��m��pm���6y�A�S�CnNV���8ڦ�GN���Me�]�ݣ���:�P��ݸ��9t���,�;�۝��s���:��|�%N���l�=����~�����O{���f#����������-���߮s������m��-xe7����R�aդ�vm;���ΐ�(�;�	��|J�`!�|,2�%w:4��D�8aSU@I�O��b|���gVYbfܐ�*�5��A Ćt����h�vmuـ�&��iְ޳e�MQ�F)$[K��f�h��Y�V:Y: �@%u-	��Fh,��Z�1f�{�� ϻs��]��rgutB�ge����1�ӦM�y�t=ۻ��0Rҭ��Tby��c�)���!��T4֚ùs
�L�"|�'B��$��f��.h��L��a���\�h��1�&b ��X�RT��<ͅŸ,`1��҄x�cbYm)AL�+1�Ia1=,ٰ����a	�'}�Oܲ� ��D�t��pȨ��^fީI2�d��[b�:޻z4o� ����wn�	&���9���Bǚ�;��;���"b)4NP��34:XS�3����h���G��C�Dئ��PW�P?�ȫ�4�>���;E�#��O����R�������{��$	4�Қ�&�
��w`w`v�zu@�)J}�7˥)JO����{��/$�����IU4�D��0CEWW�ܥ)���.��)>��s��R�<��w`w`v�zuC>��y �YE:��X�s�;]=뫍�۞�W�m�V���l�QjB��&������I��{�%)>��s��R���9���)<����Ѐ���9����)8{�_�A��I�[%�g`�`���빂Y�'��_s�JSﹾ])JR}��Fqf	f����)+R����-��,JO9��r���s|�R����y·�JR����R�������Fo-�7��}`�)J}�7˥)JO����{��/y�o�(Ip���ppP°qe$��#�r}����g`�a��~mRT�iJ۹�X��y�9��)@HO��6��=���_{�a����bC���N:�Vڊ��u��i�7a�89-�[\H;��5TI=p7e�j�Zֳz�o}%)K�s��JR��{���ܥ)���]�E�%)9�ߺ��w`wc���H�9��ɠ����ؔ����`�)J{�9�JR��y�9��)J^��o�)J�9�of���[��������R���s���)>��s��C�)}��})JRy�u�0{�K0_~K�����S�]������t=�R��s��JR��{���ܥ)���])JRy��e��0��ٽ�[�Cܥ){�9���(� ����s����������)>��s��R���L�O� ����w�[���p贻��ݖ]$f��%���r�ԣN�Iq�f8
L}������}Y�$v�g=e�ct�.��b�{ogpX���F�`�O�o�;��G�I��4�2�n�"\���G���^���n���znO<r�� �K���Dg;� v���'7m��WA���9;���7k�6�]!:���ɺM"tb5��ͧiZ	����?�33'6?X���`�[��������ԥ�un�2�3��cb�s��C�OW&�M�f�&�fj�݁݁�|��3������H�r����y·�JR��s})JRw�/ߜ��&:Ո���g`�a�_�s
R��=�:�)K߹���)I�=֨g�݁ݽhJ ��"H	����wjR��=�:�)K߹���)I�=����R���o�JR����p�[-�l��f�����)K߹���)I�=����R���o�JR��y�9��)J_W8kVh�x��e�o})JRy�u�0{��?����~�R���~���)J^��o�)J���9�Ǚ�6o���iڵg$f׍ZeF�s�`}�OdB)v+��"����I����RWn�8��~��t�)I���r������R�����`�)J_r�k\�[7�������)JO����{�Ƒ�$��,$�0̢����lƇ,�]��K�~�})JR}�����)O~��t��3�������͙�٭�[�Cܥ)�����JR��{���ܥ)�9�])JR}��Cݘ%�|�/�YIZ�����f�	fd���\��ܥ)����t�)I���r����9���);�.s5�l�Y��z��:�X=�R���Ҕ�'�{�t=�R�g��R�����`�)K�����=�w�t��[�vu{[�ؗe��y68��%�z�6e�]�QZ�n(5͇3�z�Ҕ�'�{�t=�R�g��R�����`�)J{�o�JR����
J:����g`�a����@� ������\��ܥ)����t�(����|���I�H���CAS�޺R�����`�)Jy�o�JS҂t/J����=�:�)O�߿M��ë�߿M,n��I]�`�)_��ߺ�t�)I�~����R��>���J�	d���\��ܥ)��rٯ�kf�z����{�R����y·�JS���k�)JO9��r�����t�)I���a�-Q�ov��cS�����ck
�v,��7��qz�+���hj��D�J���ܤ�[�qf	f?��R�����`�)Jy�o�JR������3�0K0��_~���)c�)U�޺R�����`�)Jy�o�JR��y+g�݁ݶ7Tۻ��$%3Z�[�6[�oy����R���.��)>��s��R��>���JR��{���ܥ)�}�f[5�5ekn��wJR��y�9��)J}�}�t�)I�=����R�e��JR���Ü-kfo3ff�j�o��R��>���JR��{���ܥ)�9�])JR}��CܢY���~M2�-j��8�����N�n.��r77b�[vC\u��z��!F�;tl\�y��ŭ���޺R�����`�)Jy�o�JR��y�9��)J}�}�t�)Xut���KT�ҍ����fqf	f����JR��=�:�)O�﹮��)<�9�4=��B�������f��z����{�R���߿~�{��>Ͼ�R�ȁ�{�~��r����o�ҕ�%���gߕcbtnRY-�8���﹮��)<�9�4=�R�s��Ҕ��������|��G�jJ	�*R9U����ý~��Ř%�w��˥)JO<���{��>Ͼ�R��v���ߟ������F���њK��A��cn�|8v��br�Ckv�rQ^��i5�BV�-�cr�Y|w��n��WB�����I�p���#sݵݭ��'�܆��.u��ŕG��\��z�lv�t�g��嫓�([j�4/\�غ����o��6́����qv�v���KxK�Ûk���]j�HX�N7nw��U�vz�o&۩6.�=������{������w�����D��^��V���l>��h8^�t����{+�Գv�]����]h~��9Ϸ��JR��=�:�)O�﹮��)<�=�4=�R�?��~mR�5.Ue[�%�%�{�ߴ{��>Ͼ�R��������)Jy����0K0K����+��(��=�R�g�s])JRy�{�h{��,d���o�Ҕ�'����Cܥ)}\᨜'ⷎT�v���ý~��ŘR�s��Ҕ�'�{�t=�R�g�s]8%�%�WO��4�5-(آWe�g%)�9�])JR{��Cܥ)}���JR��y����)O�p��kY����h�m�뙹	��.q��o�D�Χc^[)v�廤�Uo�����{��Cܥ)}���JR��y����)O9���JR�����[�2�6f�oz����)J_}�7�D�x�8`�
�K�b�f%�B8�`�+�oR���u��r������)JO|���{��>�_sz�T���G-r۹�Y�Xw�߿C8�
S�s|�R����y·�JR�ﹾ��������,��l�9
�n�8�)O9���JR��=�:�)K���R��������)Jy�Fs�5�fZۻz�Ҕ�'�{�t=�R��}���)I�Ϲ��R���.��);�ߓ$JL���mTX<�[l�ht�K���=y͝Y�;�oO�zѓ���{s���n�W*ڳ[�{��/����JR��3�sCܥ)�9�])JR{��Cܥ)}\�"p��^)Ru�w0K0K����3����)����t�)I��~���)Y���]��ë��~�[���Q-�����R���.��)=��s��C�Q_:���:�JR��}���,�,��侮~��P�ڝ�����y�9��)J_}�7Ҕ�'�g�懹JS�s|�R���½~�3,�f�oz����)J_}�7Ҕ��	����������o�Ҕ�'�{�t=�W���������gb�<��ܥQ�-���!��w�e�ug9&WaP�.Kn�4I�y��[w0K0K����g`�a�߯�Ҕ�'�{�t=�R�}���)JRbBS54�5TEKQsW,�;�;��R:R����y·�JS��3�)JNu���g`�a���ɔ��F�ʬ��)JO<��t=�R�}���)JRw�{�h{��<�7˥)JN�Ü,�ʷ�Z֭Y��=�R�}���)JRw�{�h{��<�7˥(IOz�2VFb��&Ib����#1H �1'	X &��������)J^W8kVh�x��n���)JRy�{�h{��<�7˥)JO<���{��>�_s:R���:x`�߭��T���cX�e5���<�I�h��E��[_0�4׭m��;���#�l��}o}h{��<�7˥)JO<��t=�R�}���)JRw�{�h{��ߒ���&��c�;m[�%�%�{�t=�R�}���)JRw�{�h{��;����0K0KtK��������K��)J}���t�)Iߙ�9��R��J�n���}�Vσ��l#TUII[c$�T�s�Ý~��Ř%��9�])JRy�s��R���}��If	a�ߗ��YE[kvl���S�s|�R���
A�s�C�)�5��Ҕ�'~g�懹JS����G��%��4g��(�t~0��ç�u=E�/�(1�!.5�{�ue'I���A�l���Yj;{`�H'Mk@'_0��B�w;�D�B9IE$+�N$�w�a�4u�O�z�J�N�Ka�4;yjޝ9�da������٢�͚p[8�1��s��%��-����ݴR� ��$c���`Usq$pbX!`��KL�y�O^Y�������K7�H�'����')ey�����j"�{��{�a���p8��5��3Ek��'w+��gn�n_:ăz����z�ח]xt��6�		62b(
gG�Y��gp���pF�Ś �Y0R9YE��7�ĮT��V�Ndfu�3Z���5�j�j3wf!�64�A�d�I!bOw�N#��!���{����M��M���Y��9w��ԝ+-�嘺�]z9��:u�j�����J>��';D�.2�9����⿆�{o�   Hm�p��	   ��   ��f�����XÎu%�2�p֙G^)e1��t��6�zȰ�]Uƶ���3�і�ٺ+�ɮQ��ս�洑O%Ћf�j�m� ��@ ���m�   �m��$!M�` 	.��m� �6�3���ۗ��A�i�XFyg$N�*��di������#�.���F��V�9I|�t�
{4t.D�Zɶ�睔�=t�5Y6�p-�K�ͮ��oc�t�\��ݧ{H�,v�%ͻv+@���L۵�+�q���j�mP
���*�^^��|,)[d�Y�rNv��=̹醫ZOVv�.��m�5vNSK��0f�t��[�5]ǵ`�xbv;g>E;IV�Z��<)v�r���s�\\�mFQ��|�CmX�,o]��b��ɢ��LvQ�Վ{>ݐ�Z��A��s���3��`��[�T�@���&�;\襗��ғ��Z���C�vζ�8��W�1���jv۳��B�E���Y�o>P���z��e�	=1Ʉ��Y�^b���):\�iu����F �8��T]͊uv�rUV�9t��n1��%��rX��.0��lq�-�U��ރ�\���m�^�n�ێ*���ݨ闑@��Y�׾�/[�I��.���n*���j1�f6f8G�H�N�iW��WH�����gU��MElUN�U��L��e}�]<�c.����dۍ�\�[�5s���Ns3Պ��g��x�sh�붻V��8�ވ9�Q���:E۫v���u��+I��G:�N��23�
����r���ۀw:�L��\��6��'kr��d�L��rt
�a�n:�KoZ>�x麞���4�=T��	�Xgds+�ED�����-�;ظ��=�9kkp��y۬�dD��8��'�PN^��i3u�kG[A6m����n��<@ \r�
���@uqm�g��/�����Yc��9g9�:P;� �D�����>S  ��&�TS��������ww�G�/�Щ)TQWkhJѱ�d�lev;ډ`����3V������]��L�\u�s[,�K��]H[	u�q1T u�g#�Սl��G]N�v����-��=���7k������$�����[�[�tb�_����Ѯ6��Jp�D���bѢ�����{m�g��z���y#bն����X�k-�z�Ln�Bԓ7!b�N���Z���w����$��8"��$�Ud��G�8��w(�s̳n.�uf�y��#]����6���4F�Z�mݽn�JR��>�~�{��>�_s:R��������R�s��҉f	a���?~�IZI"�ۦqf	)����Ҕ�'~g�懹JS�s|�R����~�Cܥ)}\�Y�\-�ku�[�t�)Iߙ�9��R���.��i<�߹��)J}���t�)I�������KJVF+��3�0H��_˥)JO<���{��>�_s:R�);��ߡ�Y�Y���}\�RP�JӶۥ)JO<���{��~�_s:R��������)Jy�o�JR���,3�9���8�:pr'Y����'v�ٛl�����g��P�v�w��M�}��^��u�l���)O���Δ�)<�9�4wW���&�p�m�t6�$��m�U����}wnbB��2�0�+)��Ŋ����0il'Vh�ZD�49�Qf��X�� f�	3@iQ:^�9͢��-Y�nΨ��;3��q�3SLTCCUDT�Us�{���=����7gU�|�E��B�Ң��O�f31６`��,���pv��X]R�J-��$�Z{�w)/ ��:-�8`��n�ߧ�U�c�I�9s]%�(�-��fv��7%�0�z��¥v^�%73�]$NE���U%z��g�N�����www��)������lt��db�.�$�����ď}w)/ ߔ�	;Q$ꬒ��jK��߹ė�Oߞ�ǰ�8 ր�܊J�%	I)�PRQ !���������pʸ�3���Q �MTT�V`~wv�fwd��,zyt�I��UW���f���wI����Q5�O�,fw�v���K0J��}+�W�X
�V�*$��v.qۜ9�Q�n�S��K�8��벻��5vz�SM�
�C����@�0}w)/+�~�7�:-��#.�"�i[�ƙ�{�j���7e(�3�Z� �T�vwWT���n��I!���K�7�5N�����Ł��ـ	4�,�*�
&j,9�ݜffh��˧ ������~�}ׇH�� �P�Y�^f��%����N�];��h�� ?UUW��L�;���o�tZ�����O�g�w-��k�`�'��z�z.�D��옜������-�+6�c�{V`�J,�V�ww|کy��eD�DE4L�T�V`�J-���ϥj�ک�����ݿ30��(�tSN�4Ֆ��vӼ�/���tp�=��n��R^�"m:�]1���y8������;���߳�`-]�0)J.�_��g���ߵ�^��a~7�̌��2����ｫ0vfngfۧ��������@�8`���Wwm��m�����|�s���g��p(�KW/- �k����eN8g':;x�h�۹q��ub�7�Y��sm,Y�z���Fh�m�ԻG%��Rp�jc)�5���X��������PMG�7Vۣp����V��nX���/��x7#�����	i!����뺃�5��y�obŵ�@]+��t�;��26�Z:���l�m7oIa-�s'5a��Zk
�v-�[[sg��5J��34T�3$�5��twt���)���B����)���~�w�W��Z�!��R�d�jK����qf��;����ـ(IM��|۱H*�j�b��j����T�ｫ0����;33�g����~��+����B��i����&**jh�gfg�����ـtwt���)��ۇvn�,�����"�-:j��\�`��@�8`}��K���g͐�-�V8TWqWlR$�ہ�sIm\�c��3��n8�����殮~�{�����'t�b�J����zE�I0���vw|BJlHJj���!�������T��w���ݙ�ڨ����-S`g��?3;��3���M����jh"�"����uw��$����������vfi����p߿W��M�	13C��B-=�%��/H�	#�������0���j���"d橆�h*�jl�|�����3��ÿw_���t	rE�o�]�V��j�[����y���v�q����#�C�ˋ۷%#��]�n��I��ltҧ�Ӽo�$p�>��s���s���{ZP�+�u��ӀrQq4�DM<�1QSSE���ՙ��C��hT	X_��?��~�?��wW$p�7�	ߔ�Q��Ztշ��"ʻ�^���xЩ�M��0�óY]�Ł����#TUMCU:3Z�n�kz꿈	�\Ph ��}��~������>�ڳ�;�OwM��q�5SPE�T��M\�	*E�~f���a��������6}>I�m�ӿov��`(��InW��n�ūdO&�p� ]��j�T��VZ���9� ���fٴ�YWlV�L�=�۠K�,>�%8J���w��n���q���ի7����~��]B
G��P�����p߿W����%����0����!�?~i�&O�AU3S`n���pJ��}�����X���s(ltҡ�0�Us�;��3Ͻ�Ł���0�\�Ui�g�"�IY"�	�,p+,"��)`���N�N�U?�" ��g��~ﺿ�~��&���y"b�*��>�Y�ljS`}{��=#��z���D���<q�q�0h������ֶ9��7a�����A�i��?�2i[|��$V܊�;w�/��t�G��X��[��s�����0.���bj�H����jl��j�����ouq`}���cR�wg�BSU5P�EL�\���}�x��`�t�z��tJwN����O�f��a٘f>��f �wM��}�U�33p����|X�z��j�b
����*� �Ԧ��>���<�"�ϼ�`��tH� 
2���eq�	̖h&�LB���Af0�e�$�"rȪE\��qpb`����6{�8o-�V�pY�0i�yљ։��s�2��F�v^�Y�,�5Q�Q��+����O��𜰇<�U��s��|QvW��m;=A	۠�n�Au3�-��m�F�z�V��t�8�n��ݧnb��ohދ�xW�M2��*�=����iT㳝Z��pK����ƞ�W��j�{�^:f�8������Uգ��qۆ�B�Se�����=,��cV��[�,C�t�v�i�u�=�M�W��mƆ��hx�X�߿v�T�	�pu�V9f���w��<�"�ϼ�`��2�V�-+�*��-�ė�~���f,��� ����`���G��X3;70��r��&���y"b�*���ov`��_���H�o�.�)HWj�D�V`~vghfg�;3�w��`lj�Հy*E��wgw�������_�f����U.�i�-+Li5�}{��=#��zM�:�E�{�.�*2��ݴ!�VT�����&z�ӵ�i���Nv�t�oS`�]��wf`����,�:�ʬ�v]�Iouq`g�K0�Jl���8ѻ&��Cc�ʤ�R\��~�?�3�	�W���(BRJ�$�1֦�XLV�u��-���0�hMZC)�f�4��CB���f�Z]@��33c��fae�h֣A�TM�9�C�d������B !������$�S۬��u�\������s|�� ��B��f/����W`�+�LR�q��6�O�N��ٙ�7���>��f	/����9��%h���H��Y������{���wW?~��3�K0?;����(�b*���(�6gZ�Z���_�0���ð����n�_�(��>�wT�h��A߅vZ���7n`T�3<�+��\\6��ojwn\�>�}���jݞo9I)� �w�0���};�Y��0�;����� ����n����!Q%5�����)0��
�{җN ���=� �F����*i���1�k �����8`��~6���;�l����x���)}��s�y�4u�1�H��u�܌������ӫԇ㡲������6I酕y��)Q���N�-b9��LN�u�F��a����J��p-12�c�Љ4���ef�����0^�2�1s���~����w����(瘃h�y�" vc����Hh�����CR8�=�ZA�b�5PG���~�J����r�g��mf���m��=<~������a���P㢌=����#�5�2u����n�xw��)�l,�k�0�Έ�tF���l��
����Q�~]�����"�����|��.)(�F8( ��������}��ԗ~��~����ٜ�v�/� ����Ł��v`	)�ggf>�wT�G�(���wWun��$�}�7@�,�tZH�}�K���*��bu���j����9���ӏFu��;Wh���d�:�����ˣ�un�i��@�,~��8�H�vff�fw��uv`.�$����t:i5�o˺-�p�7��\�g�ߪ���s�n��@�Uux�-�p�7��\�`��@�д�l�Sb�L��ߪ���w�_g9�uW~k﹮�_RDY%G�f`�� ,�w�ԗz%�쟈�hrKt;ot�"��U�~���� �{���_�-Ye	�4XZWV�����TqiՖל&Ml�nv�ϛ����e���{�[f[i��!%i��X��?���8`�t��H��H�ݍ�M~m~�o��8eUW�7��\�`��@�븹M:.����ę�o��t�"�����ߗtZH�t��j����Z{�u��.���ff.{�~�H���E$�X�����>��8�H�3�՘�Jl	vf~,C#3�
�IP�{����U��[���p��gv|8v�j+��+�lU�v�v��Dʻ��cZm�=g�x랒C].��9vwA��[t-��m�[�su�s�x�o6��:�G���l�e�'F@�Q�i5և��j[��l,@�;9�OFwu���b�\�ۚ�iޯS���|}s���s{6:�M������x�L�]56�:;���9:�C����������ƿ}�#/��{^2�&�t�.��� ��Bn	�n"��q�[�}��w��غ!�Y��sW:yW{ڳ �IM��O�Nӡi`�B��%v$��o��~����l$��ϧڧ ԩ����g�]P�vU�����:� ߗtZH�o��t�t�Ӱ��+n������ϧuN�R,��f���d����j�����:G ���'�ȄJH�����וs?~��������T��j��vӥV�7j���!�;��Zնe����E�6��zqOG\�ۗM�ݗC���3 �{��rE�o˺/ʯ� F�  @Cʹ���] �N�c��`�fb^bk0��ܻ;���D�" �Ԇ(K�;������4}�S�ym"��{Vg�Ɋ��	�PIP�wy�ߚd�?4S�3S`{g���	*E��ٙ�#��ـtwt�BݤU:�V�'���^?���0���`� �
� ���u{�~�w�}���^�-��രt�Sb�W�n����w�_�B?���
����߫���`z7��`	*E��8������ۭհp�y�s���w<���Zz�i�\��z����V��p�v���BJl��U`	*E���8���0��������:8]SRUЛ�i�o���	#���M�%�s](�XY% ��?~?~խ�-�s/SO�Uu�wuq`g��0�lgwq���R�E�{�H����r����:7�n�?��&y����u~���� ߗtZ�� ��+�6Յ6��N�[ﺹ�s���C0�Jyz�W�r����{V`	֔��������t�ݓq�7lQOE��n�u�F�[WL5f5�ة�I+I��t:v��6��j���.���~�b?��@iGʺt���M�DT��5L5��� �R,�ڳ Q�M����V���3㳻��;�A����)�&��&b&&h�=��0��jU�-T�<ƭq��[(ֳ6�7����I0���һ���<�� Z�L3���;�CS"H�� u�{�>��KR�Bm���n�M`I�����ffa�wg��Ł��� Q�M��������ߊM�ml2�g�;r$��7mѓ�^���Up-��i�]p�ۍ���S��]`U"����0��73���_�����K�����i�b�&�����jS`d|���R/�3��%��P�~�r��/���e�3y�KY�tw��`d|���R,{ڳH���H��X�J�R�f�0F�33��3;4}����7���=�j�a(��ӝJ��ؿ;��x�-�p�9���aݙ�wW_�(��3�IN~w}�ww�����B��UUl��p�;��=�T��kJ��E,Vy�['��Ҿ\�G:�����8��3ף[k:n��5�=�]v�F賛u�n�g=�<rځٗ�N:�oo3� R��Ϯu�dmۤ�M�/���ۊi7iӐ�4d��:[RP}LW9\W��ͱ�.��Γu6{b
w�ܻl�[Q
k��rٮ/k�/.n��.��C�v�մ5���s��gu�ƻp��-�x�$�'�l���m�y�ǆ쐭P0ݲ�mu�hr�34|۫� �Ԧ�ϥ%?��fq�ggv���������.�y�jx�)�*� �IM��J�8�H�=��fs�@b@��/����X����+�l�<�pJ�`{�j�a%6{P���*i�z�zɻ�xfq�gw]�Ł��ـl$���vwvv��\�pCj����� b����,}�Y�~q��a���OwM����N�R,�֖b��8f�V�:n���k�Spu{x�p�0�NͰ9��7U*�r�;U&�!^�߯���Jl�V��5*G>;8ó�4�Wf 2�ffy�*Bh)�f��ϥj�|4#$Ī'$ �p���U!��@������n��{��rE�}~��U��-�"j�h���R�X}�Y��wfo����'G�ߦ�����pZ�����hv�UbI��{��rE�o��-��gv�|X���疩�a�b�i���:� ߔ��� �����c�a�~5v:��Wc��e�b���� v&v糛��s$�8텪n����5��7WI�iӴց����ZH�{�t��H��B!�v7������ZIH�v�ݠ7ڻ0�6}+T�E{���*�O�f��t�"���)`�	�0���W3s����)�\L�1���,G3��ʰ�T<���[=ޜw��V�0ª�����fX���\�`���8`��7@+��f&S�SPST�M��J�88��˺��7ڻ0�����&&QMU�q��[��.���(��쀫��N=�`�<�����Z�u�hv��v�aK31h#����՘�Jyݱ�ٚ�N�N �qiV:alV�ē0��M�:� ϧ�N�R/��ggf��0�zF*jXh$�b�0�6}>JpJ�`}��n�C�jR�I�ݴ��k�~����S�%{����k��?��]U��������� S�w���;�%�[��-�pʿ� ���}�?:������3��S�o��QT��S��I�s��Ф=u�y�cN����s6�F�N���J�U�aLI��{��rE�o�tZH�t뾻��V;�wiU�Mf��Q|�;���ޞ]8��������A]�?Ֆ���x�)�p�V�t3�3��{� �OtXv�4I5,=DL�4]]��v��cX���BJl�ُ���pZ��k���b�bZ&&��}� �fvn��ޞ]8I[X;�;58�����޹ #*$��(m��<Z7��F�a �Z��oC���(0)�����&�oxt1v]E�f:�ө�줖�E�M�f�`�5jѣ5��ێ����4Yj4�2! �ᴴ$� @�w�Ot���ko�  �p �`$��   r�  URhx���ôAon�6&�G,p�1a׈1���j6��K���ʶ�$$,,�;��)ʝK%r��ٜ�͠�u��9z4L2�T�D� �I -� p�H��   ���%�sYҰ @@6ٶ�[��n!`�/m��jF�l��`�v�۴�=�Z\ٓb��<1���bu���<]{l�&�����q�����ّQ
x��=Tݭ]\���iu�X�(�Lۇ=����t[-����<\��Tqj˸mt����m��u'a���%�vgl,�gμ8G����q��f���g��vwP�ʰ[� ����Al��;!\�Q& 7':���!]s��s���+��s������Dv������3c�'�w�������H��'5�׍�N�HLK�Ib�`,�7m�����45�PEX�5Tk�r��)�7P��j(l!<�U����l��U�c�ܜ���<ڀ�N�����LL�������d���]o)z��� -����F�a�˖n�±��[��q��WV�u�q�T�J�G�V��٫�����m\��NK-E�+��-��	MHi"˯C��]�!�Z�vD�t��6�и������DqT�/Q��Gu��֧d��UT�Z�^q�n�(j:���gGHH�Ĵ^Vn�ҵ��UKe�]�ۆӮ��祓��v��s]� ٝ�c����^�=̇
R]�Ȅ���ގN�1e�*=���jGwaNr���|���ݴ4��4tw-���բ��7Q�`S' �zs�i� ���v��(!�����ܽq���uW3���;v�͛�kKkrlm	����]Vx��U[:��̚;v��ʬ�vi��b���iS$�Lk+��:1�-��Odkyӵٺ��n�Ҷ <������g.sOO+�W �m�H�ݲ�n��ɱ^�۝�6���8�G]��n�m��`��a�3�a�D�U��������n�_���n�Ɓ�"t�YC�b�l�&;�1ܼ�+5$����d��s��z�z;p����[���t���X���銈�86��r��ɮۧ�NĻ�M�����n���Ok�ҙ)�⮶9=�Ŭ��_%��A�ٸXv�#ٶ�ph�c��grn�pv�f�m۵�:m=a}Lwn�c�i�u�*�u`�r��:J���k����JT��I�c(�Q!5'���l6�����zY�.�j�Ʋ��A�Y1�ʗ�����ߟ����6�J�8I[,vvx��� ��jR�I�����i5�}��:L��y,�jS|��ߡ�ݤ5~��J��*���������?w����{V`
5)�7�����u������M���ga��=����wM��ҵN �+k��Ҍ�V�ҫV���E�o��-t�X�{��:]*IU�'b#�J�uޝnݍ;����+��mɺК��4na�E�F��nƝJ��5%��~�4	�e`}K�����'u;�ַFu�]k���9�׊�PNa^�ڕ���ݛ3J��0�"B&h����Iƌ�%�[3F�(b"�0M[\0SHl��2���0�u1�a� g�?�g5�_��q%����ԗ;="�=:�c�PҵV�7X�{��
SgC;4}����;���|�
e8�TU�vR��@�$X�/H�	$��>��n�q�jS�I��&��i5�}��)��֥m`}���F�6����ߖ#씮E��ʵd���+�����i���4Y�ڍ�r%N�:�n� Z���６`
5)�fw����N�d�:�j`����k�y,����ޞ]8���ZF�Ҩ	��ZUj������S��UV�(�^��Yi�!Jƌ��֝`;4P:�19�t>*�x��(�s�{��_y�9�t�D�D�����
���Ù��=��Ӏ.=��f ߝ�gu�����B����Rǘ�	$��=��n��}+T���h`�����������m��6�CgR��^5�����nϝN�������qV���P�iՍ7_:��$R^�J�,�����������`���C�����K�7�:-��X��߹�����# �����WIkJJ먩��=���N�+k�{V`�(�1h��-Q4Q4ԍY7s�3�3�˻�����T�������1�-S�{�t��J�YNݟ�n�}tIE��J�8�����ﺺ i�"C�<Y�GV��s��m�e7D���շ]qK����Z�ƕ���a�̷��2r���T�3W�;���}))�5%m`{�՘ ��LDJx��"��*j,�RS�����8��3��w�߭��~�T��'8��@��aW�1h$��=�t�����I�'KWX�T4�{-淳�P2+�}�?w�\���׀o�H��e`]蔧wi���;(M��Ix���@�&V�{��WK�၊�&K�8,�I�.f$3D1I ��1D�ꪪ�;Fi���E�э�Ʉ2�tlWe�@XlU u3�x�$r`���Lq��a3ۼ{qȻ���.���=1��p<]s��n}�ޱK�m�k ��8y�z��Ϸ9�+����q��[	r�m�\��c���W/Ss����G\˻6�.��$9��u��Ri��Χ[	K9�Y*�z�p�w07"3:�;�TJ4�Z���B�3�f`z�P	*�2�EB@�
�JמY���g7!�8)��u�c��j˯X�f� ��p��r��n�c:F亭��v��5OwN�+k�������|����J������������5%m���� �G+�����t�E��JJp�[TT��05E@�5M`{�՘R�Y��zR�$��~/l>��j,�5�U(~��Pwqݒ����һ� I+k������ 7	�H�爊�*
h���>�RQ�33�w���������)J,o뿮<c��+i����{��ݷ<�ׇ�3�i%��=��7���������-�_|��I&V�zM�$R^��H��-Y��X++�U�MI{������f�������n��óa�NtX	OwN ��X}G�JN�Qv�e	=�$R]��Ғ��ۘgh;������ �zԧn�Z�j�;�>�I�$�X�H��zT�j��Θƕ�ɻ�RV� ���{U��(�3�I?����������/�nL�B��������hyp[Z���,����&��y;:s��Gje;vSu�wt������I��L���Ҏ�M!��X��T������3��C�?�~��~�m`{��]�\��?]۲ݎ��x����tub���1QL���9K.
FH1��+�']t�n��Ix�"�wj��];�l*��N�fwx]ݍ`n���5JQa���z��pˢa��������
���=�j���JQ`gʒ�RV�������ۭ��ˌ�v��m�#��n�u���M��/.��uveuv�A����:7j{�tR^�G%�$��=�t� �{�_��b���ଯR\������3 l������T�52RT�D�QCT�5F]��U���{V`�ߢJ��>������K��*e;vSu�{�K0S�,�T�`S3�7������~��t���'�.J:)4�v�!7��� ��|�(�5j��=�j�Y-s����1˚�:�v`��n��؎j��]���u�'2�-Z�Z��7��F����3�IF�U���{V~gw�t����+�"bb�j���h���V�k�vv�wWf �WE��*J0M�&X0m���m��=�I�E����K�:t��;��܈`��e�؋opf�:��ĩ(�5j��7wV`}�N�4:�nժw�l�K�?��ιv5��]�������332UU�ݧH]���d�le8866�3u�Q�ٹ�����a:U1��j� q�k3��n����5(��A��`��k�f7MU�u�
jj{�Yݍ�3=v��$Ld�K��gж�]���6z�����qh�,Z���M�][�)�V��mu@����K��n������^5��2:�	`m�`��ka�;s5:!�����{�ݷ;p��g�&˶�U���n\�ۗ�93�:ۅ6�q�!�˝b�k����j��1�t�s/@��+ �t]/ ���}Ivۥ�ANݍEU5����9���٠]+������ ��+ ���t���Hv��V��K�6G%�:e`��t��\���	�;[N�*�#���2���\�K�v��)�+aV�2����+ �u΋ ؤ�@;��?�$�����z�F��Ӊu&�{>��g�Ϯ���&�v�]���:����W�X*�����Y�l-S`b�����[Xͱ�MDDIPIY�l-S�J��]���;�us�s�����+�DJv��`�j�;M`�h:e`��t��`����r�S�U0Փw8���ιv5��]�\��H���.�t�*���f��7@��I�Ӝ0	��߾{����Xē[��y��h�f����n�ζ@x���>cZ�R߮�+c���.�J���@��I�Ӝ0��\z�QjU	ն��I�b�-�8`��t��e~�\��v��r�	�����5m"��n���2fjt{d���٢N�}�&@���\m�1����;�ǯ:�Klɍ�Ua�ۺ����\���6&��8��,X�K(�s
ɥ0
b"��* ����&
�3��<'�4����! �J`���J\��dX!4m3Eo�����z����ь۵m(���v@�$�`a`I�����˽�-��ty-�oɱ�p5f4)���C��.��f�pR �S�9ۑa l�M�aD�JTf���ߞb�ꀈ%� �G,'��Wa	�î���]�_�Zj��֎s��;�
��آ�$"� &�?21 �"Q	 ����x�!�:S�/`���(&�> N�\@S�?�<A9��>���$^��ZJ�%yn��J�%@�f��Y�l-S`b�J0gմ�~m�P������j�H��픢��>�}���q`o�V`ӰȂC����n���e�ma�K-m�4l���뇷����0�OV{3���z�B&��m��������p�'���~�>�%������%5U1Ee\`ݤ_3�Aڗf�=�x����}ʺ]��~V�e1�`۫0�R�g�IF��E��/��	��ժ�i��)/ �s���~�|���WB�������^�(�*���V��x����W���p�'���r���qjի��n��n�7%cV}SZSS�5�݇��m�nN�]8gmWr����o�C���e��p�'���tp�'����D�-�ۧt�X*f�{uf�j�X� ��>���)�t�ӱ��tp�өN���q`v�ـ����)�������"���gq��;һ� ԫ��'���tp�=�WF5MR�SSe����m`s3��j]��yuq`s�}�k��M@0Ĭ�S�� D����s9��3Y������/%��#��y�x' �Z�V�yYK�W2���ڧ�71����}�k�\�=�+��N��en�ɻE��#��yv���ø��ܼ�sk�<O��4;�v�GN�2��k$nb�V��<�Kr˦�t�+2��]�B��1���9�F�t�
j�;�c�>���k[�'�2��g��g���,�b�e�s�RJ���w00�3���ĎTۊ��e!`��;q�s���ݒv��G,�r���#g}�)���:��Um5%��}��Iw��>]"�=�2�	!|](�M'v�-Z{�}�� �.�h�X�j����	�%3MSTX����镀OwM�>��K�m+������@�t��'���tp��UD�t�@�qQ+�lM�T� �u�OwM�>��O��h�X��?1��VUF�� ��vᑸ����f��l�cp�j݈9���jև���IY�}��`/�%8�U�3�;�@rK� ��sMMM%D��E���9�w��H�Bh ���gvw�:���]�ک�2T5M~��i[5f-��+ ���t��tp�7�$Zܫ��n���[���`��n��G~�K�=�2�	8�!�PQ-Q1$�U�ک;;ó�����j]m`{�K0	f[�!�B'�4 's������cq�e@�İ����H�z�"�����m��:��[c٠}��۪�����9�ٙ��������;�q31LD�Wf��mn��훠}�� ߤ�h�*%��v�j��5M`{�՘کyٝ�#�%x`�X��w�R�ڤX�V=�?~��8`����+ ���t��D��Eӫ�V[f�I��=�2�{ڳ �U"��gvf�#��:����&�rp�� %�ڸK@<ɇ����ŷ]sTܚ;N�YT�9`�u;��������}�� ߤ�hu��St���7wLi��{��tp�7�2��V%.��;L���ot{�V�I��>��X�u+T�P<E1TTDU5�;���G���0ou�U{�s���?*��cfh������N	��k�4�ȿ(;|��q`([<����a�b�
�� ��[X{ڳ ���`gڭ���1�
���]���'n�@�C�\���-�G�N����/�]���V��Jg��Mw�m�~�v`��,�U��;�}�>����H�{�{��o�2ޓ+ ����Uv�B�"�϶����j9���#�{V`�\X�R1�7��;�+cח�}�2��{��o���^�J��vSu�}�t�����zޓ����z	�H�%œK$ 4��ߚ�	ح���m}�*y�={N�':����6+��Ԥ�:Ypjv���)���rsn����ŋy�eN���s�pb2�n��Nݞt����Տl">ݨ-��ZqH(ո�mzN��-ݠ�hM��4��`,"�*�Ys��q��a�uo>Va�nm@���������w]�Ղ���X)�L�OZ�m��tӖ;�(s�õup��0n]�z.,�m�e��v��mgb�]yNu�ĵ�M�\���:^�^"�v�۴Si��ws��G%�zL�Ӻn�IµBR��um���0�9/@��e`��t{�0�E!v��0wq�}䭬-՘s;3Dn���^���!���T�UUK05Ma���Ѽ�}�n���ߕ%�S+ �8�R�6��VЩ[{�{��w��zޓ+ �{�ګ��&�8�s����a�[���Ih�g=�.%�մj3D����Es�ۣ*��~�����&V��7@��K�$��m��r�H�yu�%�~����0�f��U6zv��=����9/@�׺�!�����P54����ޝQg4B�W^������$R�4��H���hݥ�`/uwF����<�V`Z	RJP
�&�v����K�>��X�t��]/ ��z���"���t�}u�x99�����y{�I�ʘ�V�0��A;�g8%��O.�%n���[���>��X�t��]/ ���Ex��m��J��� �{˥��r^�������B"����i4*V���^�I�.�`��w�h�T3t!�N9�J�iN�Z���$��N���*��M�j���gxwgfx���k�[ـ�����ik@;VӼ��!�}�2�N���^$��)ZwE����}䭬-՘�:��ߒ�`��,�7����&��p���;c���n���E�c���f��ɝ8�Z�rs�D��ly.�ޝQ`o�Z0�����7�d����j��j���=������u�{{��-՘ ���L�a�)��ݤ� ��hzL�Ӻn��.��m�G.�%n���L*��4�&V庳 ��TXS�;�o�b0jM�v�݉X4�`��tyt���!�}�2������ƕ�����'k�5��mɬ����]��[b�<:GkWfG����馿+Iա&�@��K�;�2ޓ+ �u׺!�l�$��x}&C@��e`��tyt�N���U��C�Ҧ��}�2�N���^�I��=uv�O�C
cN�N���^�I��>��X���R
�4���Si��.��w�Z0����庳 ������S��2��ZD�H��P�}�.0&�Oa�,$�N�)4yo����]E�\("���񶁊w�G��)�#R�&�I��ol��΍ӽb��vj,2��tA�4�TK%խ�ZǮ ���������#���P���2j&�zm%�P�`5���͈�A�T�h�Ȝ5��F���e��@vx�'K U*AM:]�-�Iы�����s]^��dE�QF9��&�4:��tk�Q��N�1�[�Df$�)����6�m��m�� pk��HH   oP   T���+n�Թ�Z;7j�e�]���ۈ�^��	�U[jYdĉ� �׃N���Ω�n:k.�v�ri��mc�Z�i݇.3t�4؊m�m�À	�  [E���   F�ے��m0	� ���ZeMV�UN��8�v�U<c��iC��1½Q��6^�m�br�jLP\;�x	5�:��Rni^^N��qی�H�'@�k�;�c;N��Z��l��X�x�[��d'88S�)���OON�� \ut�Fk�3���Iؘ�Ug�28���3��lTۓV����[7o]��ѹ�.���pl�Q΍t�ե�I��sS۷+�.��-�`G�����֢��!��g:�=ɑ�+�P�L#�vI��+j�����cפ ) �v��n۪�#��Q� ;L2����
�me��Uk��f�ѫ����F�zl�(9��^u��N��4�.1�gO�� �
�bA��AN���ȡ��Z�r5���v�H.o*\��(ӎ�����_=uV����k��݁jP�k�u���ɫ<
����TA��K`s. ��vl;-��C���c��֌�rΛr� d)ӄ��1�F��i�Xpݨg�G㇄l���pUUX�U=.�,��6sU��Y��Ӷ`㎉8-�|�����]qU,��Z�XL�kc��<�s�r�i�E����tp.�=�Wh��b�۰h�i�F�n�1��2+��+�1/2dL(s�<q�7�g��!a3	N,l�]��ӌ/�87ió{mǴ�ʼ	s�;q����u�]-�4mv�&���=�y�x���۸�]���F�p��f���6�F^j�������eXn1�M �h늣m�쇶�ݘ�l=��Zի@�n6���m�3���].���nە�u2��!�x�Ya������n˗K���=����.x��Q�m��ʈ�X��M)m��m����s0ᘿ��b� ��E3����l�Tjj���d����gv|8{Q,tWFW0ث�n�ۈ:�Q�h���jI9):�y�Vړ�T���JM��mm�\V�gp�9㋴�rf���7�;�ܻ�B�\�8��8����!����Y��Z�����nF��dC� ]���0�<!�s�n^B�ӗ>���l]��Wn�u7n^�`�OQ�G�U%rֲH_ `t0g8�=���M��f�ƽ\�h[��-Hl�뱀��k��g4��hZ���y[���t�'�C@����=;�����H�b�n���L*��4zL�Ӻf�JQ`o�Z3�� �~鹚�����&`*j���K� ��(�7���V��|�J��봆�V�����L���I��zwM�:��շE6P�!6� ��h�L�Ӻn�����o��Wŀ�&զ$:i�&^��{��9(箲d�t��,�t-��k��N�%N���4{�V�}�%����K��i�)!�1�XW���w�a�;�@�)1q$1g�D�@��g����c�d���E^�^]/ �t�h{�V W���iYn��Ot�����!�{�2�N�U��J�R�ZC-'x���t��=��tyt�o�2X�N�÷l,o0�>��X�I���^�!�p��5n��ub7w���.l�.�܃�lfՋ#����رJ;^n�ܴ�M6����M��n��)/ �I��=�2����D���Hh����R^�!�{�e`�&�u�j�)ۺ4��x�L���I������S��,a$�8�`ı#�����������\^�EU�5=134T�������ư5wv`��vf�]���ڢ:J��ի)�BN�t�tyt��&C@��e`�u*��2��e�m6[��xg[�ka�t�<u]�^3N1�Ļ���N�ǣ�6	�Wn��otyIx�9/@����=�M�:�_RT���vZC�I��T�g;;����kWwf�N��=���bvP1��3/@��e`{�f�������ګ�0y��j%�ղҰi��>�t��$X����`؂�S����:�Þ�ڵp�l��&��{�H�r�-I2�t�t	~���Anۺ.���oL�=�j�+Z�@\�נ�wK�[����]s��[c�j�	5m�ܤ�@�L��$� �G�N�m����I3q��$�+ �I7@$����=��]�;N��X¬I��n�I#�=s�z�e`T��`�Uv�)�V`IU���JU�$���3��B��� M	�Zfyƨ"d����е*�J���$� J�g�d�46�ݷq�ݻ��e���RR�����1��7� +���%en��+6�����_9hݝh���9��:e�{6��[vw+ӈ�5�>^��=�-��qm�ۯ�̧��.fC�����r�vc�b#��uٶ���~�1���0�N��wcO�s���R��d#�nhz��\�n8fx�f��c�|��a���c�5�.
���Q��T��V.W�ϋ����j}��r��"y+���y�<ݖ�@�2�ɕM�.;d�y��U���0Rq����ɟ���TPE��ת �7V�����:G�I�E����v˫E��`�`IU��Z�`	%m��� ���9�悪 �h�&fk0���Bԫ �L��$����[c-�4ն�\��$�XzI�$� �5MUQOQ-LD�V\�� �V��-�� ���u)��82�"$����H@kK���1.��k�����S ��W3�٩ĝ+��hv�4U�
�'XzI�$� ��H�	$��>�?z��4��e���u\�9��&�`���1?�&���
1̌F��D�Q��LđI�u�8a��3h�6�T�3i5���h��4��)��(LrWlQ�#�4"kX����Mj���Mx ��B���9r��=�`УZe�e5DD�SQUV��(�J��x���� ��Д��)�
*("��� I+k�If�$�X� I�Yi���l��[M��I7@$����=I2���X��%�$���}���$�,E�$6v��n1�jݤ�Җ�]�C���6�$���<��!�I&V�I7@�tCV��j�5m�ܺE�I&V�I7@$���D�n�v���i3^b�$�+ ��s��ti|��	%	�FX  ��\�# p�3!�1�ĄHeCS� �a�fgv�_U��RS�l7�
J���"������ww�.�� ;�����H�	$��:��_@T&�4�)��@J�n�Q�$������ �~H�c�a��Ff�;����{��9�.�±+z��Y��Db��׷Ar򵍰.���K��$����g;;��� wwU���"�`�ha����j��J����t��H��ό��r�V�M˫E��`zI�$� ��2�e`S��D�-SjГ� �J�>��F �V����,������0��D6�Lv�ݍ5m����$�+ ��M�	$x��/�Kwwn���[e�;�L���+��W]pn���C�ud��u�t	6�j�v���4	$��>�tI�t�h�D6���"�h&i��R��I*�>ԭ�e`�~��
�Ҧ��6���<�!�I&V��7@�}IRJ2�,Hi�o ����	$��=�&��$x�"��j�WE1�f^�$�X��� �G�}��z:�=n�� ��l��l\�l��Lv�9�Z�yjVjICA��� ��{�N���wλxc�d�,�tq��C���3[`x�K����X��s�gq�b�������xe��:�7n	pN�.�'�y%rm���m�`�2;5�Ʊbۊ���qd�=���:��C������&���S��������#���4cf�H�dx{�r_�w}��/��]��+�۰�m8.2&��:��mv���g������`�]��Sp�,p�k�������0$���U%I[X�cfa�YM�ڦĒOtIPtr^�$�X��������wv������}��z�e`�tI=:6�_�Wv�ZLop�$镀{�M�	:<ޓ!�zY�v:AnʲӬޒn�I����N�X��~~re��\Y���,����/G
&t\����4��-�c�<y+g����otN� ���ht��=�&�W.RT�F -%m;m��������;�ȕ+k�If %���wwx�c����� *��
�� �]m`{�M�	:<ޓ!�IR,�ӥm	�V�i��=�&��<ޓ!�~�L�g]r*�n��:i+OtI۽���w.��=�`n�KDC"jsr�g������q��ѺK[�["�\��x�=QE�tc�uL6�gT�}����2�2�zI�'G�N�敖�$���I�+(zI�'*�=����� ��:J��)�"�h"i���� KUYm,�8�ð�0w/�"y�;zx�&����h��`�F�z�ּ갳B�K,8����W{�z(p]��`=r�C����� �� f	Ĝ�
�v�r�`����Mtu���f�xbF�6j0ѣa��Zr@���ゐ�T�� �Bw#�4f�0�i
J@@a��צ�GY����ZMc�BlY)dF "j(�t��-j�՚�+]h�m�ƅ4�ā��	��4��ٱ<Ӂ�ˬJ#L�@n�кA�#���[鷾�b̌����%`!M�(=�i4�tB��� P4+��D�	ګ�@��|�,�\��e_׆ �V��BA,LERAI7�'G�{�d4	:e`Q�I7@�r�BW*�����{�d4�[X�K0-U`s;s�&�h���c�+�3�d�F{a�y}�MOl�ݭO���d�wVGu�I�5�Ė"�������?����tI��!�I]SC���˫E��`�&��	$x�L��$�X�u�D�);�T鴭=�	$x��I2��&�u��VӡZhm�M��H�	$��;����_��_I��m���MI�e\`���9��ww}����0�.����sD�tDT��Dĕ4�q�{+��;���U�9�qۡB�-Mֹ�Y��7v?ʚ��-:�:I7@:H���zI2��O޹P��mU��@5%W�ݙ�h�]р.5$� �r�E����I[CM�#���e`$��$xEˁ���.�M���/@�&V�$� �#��wG%�����ۤ&]Z-�� ��n�jJ��IF�+k��ݙ��#S[[] /E��9֢�4n:\d:6+��Ԡ,U.ǚl�������iգ\��ͻ�C�����u�!�.�^_O[�[3\u��p���R��hu�Dk������|SE����*%�]9H��9�Tx=�Zܘɸ`��]1g<�Nգb�r�p����zG���,�q�]�0�g/kgt���N�{O,-�9M�������*�!��(=i'���EjN޳�(�ɮƮ6����z�ۘ{n1r5�����s��n�K�G�K����7����JрjJ���If�۩5m:��ڴ��&C@�L��I�$�?'tm���j�t$�kp�$镀zI7@$���2�!����SWubN�I&��*��Jр%������5�1EID�f %������.�>�u���n����.1ڤ��G�T���Q�ܬ��A�$ml@xv��;��i���w�f��*j&����h��m`|�Y�����@˪�]*PQ<�5A���\����f�$E�@��%& @!%|z��>�}�UϹ��W�}2UPu{�1[���L��[M��I7@$��wL��'L���Q�5DKST�3Y������V���$�X�$���ғM�N�i�����n�F ��V�ڒ� I*�>�U��e
���1 4ēh��Cl.��Su��M�㸲���<]r�i����"�&f*+,�J���u,���w|��]|`4i�����h&i��R��fgx����u�$���34A��H\��Q$U���V�}ιwhu"A2H�*�=�ݤ���>�%��(֙��SC12T�UU�3��G��� �>�K09�ݢ;���]=((��hb�����0���>�K0$���uZ0fo?�l��\]\gjq�N����q�c��ϋ�6X^9ݛ۞)i��Wr���/a�ST���� I*�>�V�ffv������l7I'@�PD�5T�5� �U�}�2�e`wI�]{�&���Z�cM[o ��d4	$��>�tI$��m~iX[�I[��h%m`}��`IU����;<���� 8�D6�X�&"�ĝ`wI�$� ��d4	$��=!ԿQwWv��k��Z�l��OM���!S2�8�s����j���:J��ʶ���<���$�+ ��M�:�_RH�JTR��&��>���V�t��}rE�t�p2���MV���V�t��}rE�}�2��Ɠ@���D�ST�۩f�$���uZ09��]�`|����i�%���j� �S`f�`����uf/���Z��R��R�D��lX`AܜZ��u�Q�ۙ�Cq�.�v:ON��Q�\�
��N=r6�!z�"��[�ڸ����G�a�� tt��kt�d��s���n��حqv�s/gG'AĻ�V�x�� �؍
���f��7S����8�7�8<;q{)�Z!|�ipn��Lc�W������#\q�FnӲZ�(�\ ړ�S�w�����3��P`�Ѽ$���u<�QM������n��3�;:��yn���t�������_�k��Y�}	)�IUUT�J���V��wL��}rE�ot�h�H���Ք���u�}��t�H����V���}Ю�t�ʶ��\�`�2wL��u\��B�R�
��k ���;�e`wt��,�݌<������<�b��8�釷 7m���yW��]\DQ�g�����G�h�2���n�����!�x����dQ�j��vZjK�}��s�������ٮ�F%6�V�wU����h�K)�T��&�@�� �t�h�2�	��]{�m�&����k �t�h�2�	����,�����ҫb�I5op�=�2�	��t��X�L���"��*2�&�JBZ^.�Ɗ���wgع�T��WJI��s'B�vӫVSt��u�N}}"�'�d=_XwGLT���N��i���[��8�'t��'v����h�MLO<%S`w��������+�**)Hf%h`�	��!�[믺�}��}�k�=�]�eU�aj�a�{�e`wV`F�6������0���US$��c��V��'wM�>��`����+ ����bWh�ؓ��T��.�yn�K�==���GV|u�gc��ڍ�)`D�H������U��@��E�O���wL�wt���)(�i2ڧcC��>�K�=�2�	��t��X���ؿ4��I�s/@�t��$�~w��.�;�]р!)�������Ih&i���0RU`%>Jp5ޙ����hwf����M���
	 *�H�Ot�� �zE�t�+ ��n�?���]�o��0Gs��lo�4�h�'\+�&t[#n�usn���:��.�y�ˤm�E���L�N��G�z�C.ܲ�Ӻ.��-��X��t�� �zE�J�q����e�+v�`wM��<E���L�g��+%����M��7�H��IF �V�����ܗ}�(m���vҦ����"�@�L�N��u\�9����;
�`�
$`�O!M��zc`b/Pc���0iq�֌�Dc
CX�����0���"�lFU�:}f��#��E�hwo7�����	"&�`�LIȷ��Զ��
8�DGF�403!C@]�0K3,��"���n�jH&` 3t`K�M��	�j3�U��q��V+v݇,q�{x��ѷb@P�$H@�B 
!"U��"�:�Lt�)��fk-	���MAE4Ve�C&(��2�4DS4R�QQE:7�S�6C���0���!HdC���kF��������kTֶH!6U��3{�wH@hX@��	hJ���h
���!(F�d�(,("g	�uPDHT@�M`�n�A��!�"�A4��ս�{����` �O����8h!�   �   t��e���i-<�;vݚ��!�TC���gaݔ�b�<$C��O;Qi ڹ,"Zh�%�V�4�v�����,�6!���:j���;$a"ډh�E�  [E���   f�ے[A�ˮ )R  ޻m3H�V��ۺ��8��)�j¶���||����յ$�ۀ��X#�f�2�6�+��<nE�;�sO���`��˨��;rn��i��݀V�v�������r0�r;nݳ�	��Q������m��s�9���xF�8j�:4��M؜���v:�m���-�V6����:�hՂ Bh�p�gl�ȵns %�-�m�1ϳ$��3=�[���3��:� sF^�Fk��x��ݶ�f�X^�=Mzڝ����O9t�=�/g�һk $��Ka�H�'P���h�K(��;hˉU`H��Y�y���Kʭ]1�st8c���P۲/$���;rgя^-g��l��g�(mΐw��qJ�Ų�S[�{n\�܂�]8�+R�]�:;aѶ�ק����`��[
�[2�F�[�^��$�t�I�k��yWg\�d^I`��cf��ڪ��wP U�=����n�c]*m;0p���VԫV�1��|�Ms�;c;Gf�Ltx*���')��KS�Y\K�h�8l�e��M�n�8���֔[�t�]�J(M[D5�26�[��u��:��j�^z�8�ݑ#���b��vb۸�&C\�n�;a�	l�yH^U�=6���v��>�䗧���Vw\G�ݭ�v��n�n�Lo<��b�v˲�S"Z������v��A���b�=���z��)�g��B���ݙx�"�OW�5uG�p��=�5[j�B^�S��pQE#��@mg����n����|=��q�+�z:Z���ոZ�1z�j�:��s+�%/]6���ݫoX��>�X��a��]j��p�m��v�|&CUu&B)l��m���`L�9� �(�_��j#�::T�ff��w0�����cq�Z��m�/-��'��^p����-^����\�:�(��lZƸ�cnwF�Ӥ��n��n�۱��6��]�n������o�v26�]�-�-�	�00{���/:s��sѭˣw	��ݐxm���\�\��Z^�NՆ�p;�Z�(Fn��[����ɲ�P5�k��q�;��@�]����n�8�aqѣ�8���Q�{�����}�}�,�r+��m�s��RL�y=������e8��F�3�+�Z���^��
���]ǀ]���Kuf I#�$��zǉ�n��c�*�'X��$� ��K�$�+ ���:E���[��@$��y��I2�	=�t���hWjR(BCN�x�}/@�L�Ot� �G�z�C.�?U�t]�yz�e`{���<O>��}���������ب;n�<G8�\��h뺛T���qdS=̜���>�����m�I[�L��nۭ�����IU���T��@.=��`�?7wn�Zot�� �ϥ�$�����fwx�����j&&��Z������;��� ��m`%�� =�U��m�/�QN��L[�z�L�N���y�zǉ�n��c�*BN�	;���G�I�%�$��=^��@�J�j���SI"�h���qܥksSq\�.^���\IΘs]�Χ��d+n���e��=��<O9/@�&V't�U��+��(BCN�x�r^��+k-՘�*�gv�7���("���j����wu�����5����!�I��5RfiM1M�� bQA!�D-�,����C3f��|�T`۴��)%n�2�V�`wM��<O9/@�&V>�\���c.�&��{������o�>wu������wߙkJ���K�8qK�b�n��n�`4Q�c���ر`*(�<�Nn�1/N����I�%�$��$$x���ڲ�ӵi��I2�	;��I'�C@8��ݫt�պ�U�:�$H�	=2t�XT��}�&�5wV�=�I�{ιwW���uW�,��3�fc����x���(�J�R++��	yZ0%H��Y��U������S��%=����=�קc�R� ^�&;$:��pKuf�\[�����p�$�<OL�����m4���˺Um3 ��n�wH�	=2�p�6z뒲X�eۤ�D�f n�V^V�9ݙ�9uq`w%�����1ZvҦ����'�C@�8`wM�	$x���ڦ� t�Zb{��$p�$H�	=2U~�&X�v46�6�m��p�5Fs��$��\��) 5���})\ea�����5t��a�����k@y�`5�����~M�>.݀䮍�q���aسH`�}�g<;����Tm��炳�9]:ݠh����6�ln4NV��*�s8�A�	ѓ�s��k=�	�n �Ѷ�Ŝ�흃��WV�q���ژ��>�8݋��a+����\v]#<��x��C�&��d{7js�Ǘ;1�e6s���r)ۡB����뎵����DESLA�r]� �U`%�h�����@wuq`&�6#������*&� J����W���Ł�f�r����(BCN�xw�C@�8`I�tI!&:��*�"*��%H�<���IU�33�%�8�9��ꩩ��f�"b�h�<���9�ݚwV �+� ԩ^w~N�N�nx�ܼ�nM]�V���ۓ[í�l��of��0=\A��moF���~��� �:G�t����1Zv�16��L��W�?W�f�ٙ�ggg�v�5*��3�V`��$����Ұt�Zb{���8`%�0�vw�wU����(�UPSVlj�f��7@:H��L���+ �G��*��v���[OtڕX��m�G�j����-Y�{Q]�����Ժ�{��7THr��v[���x��lf1��V=2 ��]t64�ѡ��w/tZ�p�6N���<BE���)�;��ŠzGd��#�;��-WsQ�m$�.�5L�`%�Y��U�336�0���@J�!A%(.��k��G{�rUr�t˷I����t� ��K�=#�'����Ȍ�b�"�*J�&���m33��_v�f n�^�ve���K}S�{Z�e��83 �%^n$+c�6�6��,\�qri����Wo�����������=%�N��˺���뛷m ��)��OI�:G�w����>0�K�J�tݠ�;Ott� �/u��|`zM�%�_U�M6����xy{� �s� ��n������+UՁ�	K\PM)�j��tp�$����xy{� =��;�%���tK�B�؝p��Zl���f���$��J;\�&����6[`zM�	�<���w��N�\�\��2��h-7�:G�u�ܰ�>0	=&��܈�+nݪi�e���{����'�� �#�=$���j��mi�tp�$����x_�� �����v�(Li"�l�$����x_�� �s� �����~c���Z�������q6p�1��ɸp����n��As���ڎ�v� ��OF�2g�$�׋wQ&��:�]�咞��ո����̵^�'Ƨ6�nx"a��?�ˋ�'9Q�#�)����B�n۫��=�tæ+��/N���m����ڻT#F;N��݅.Z��zz�x쨛�v�\�[��v���78��nw�A �9��Tۮ��B�.�W���=��x���ڷ ʩ�z3gO������t��T/$�ϵ�g[*έd��v��D׼��V��ٰ7�ZX	{V`�E*�&�����x_{�����Ij� Z�_�v�9u�PEsH�5wS�r���K�f y%Vǽ� �{�sj�i�$]�bL�$����<���{���'�W%W(wL�t�m�zH��{��s� ��n�u���,Anۻ������Z%Y�#hmmt����vh�hv4U�<�:�+cjƝ�[o@��[�y��'{� ;�� ��5wc�٩��NT��vo;�����"[�0jU`l{ڰ��뛷m"��i]4ـI�7@'H���^�������N�I�iʙ���fw���V���kK�zM�%����TӡP���xy{� �s� ��n�N���qe�W�~\��#͚4��Q���81�n˝h�Tsv���Tqɱ~��~wr�h���m�:8`�M�	�<ܽ׀u{�sj˵��˺LI���tt� �/u��|`�W%W(vʶ��[ot�s��>׿gW��P���fĲ
Ųk�l�^�ք ��L�q4�T��-�_���H�5�yG�V�����;faI��� W����:iS&K���0�2�:M$��-�`�03�|ѭ�	Q%�"�9$XZ�AC&`S`FǠ:���Ǯ�""&4FQ�&�H�"�,#&̈����BA�.H�lنF�ZCXEf���٣F��Ѹ���Ob!" w�5���-�B�u*ǇY�m8d�0a�S5�VRm�h�F�z�Rc�f��3Η3z�=LvAD�h �b�+L�d�u�8�k���z6oqj0��¬���,Y�a'$�̪�Ɔ�IO[��n&,��K���`�C�[��R�2fi�&30�&$ �����ޔ�Je������;����� pD4'����V@�
���
�������/�}�����{�;�a�Ȍb�+t4�2�xܽ׀w��N����x�H�n�S�e��j�[�tp�'zM�	�<�^��=��{n����+!q֗�D�6l����iꭄ8�����f��\�uDK�=XJvـN����xܽ׀}���=]�t鴨�;Ot�G�{�u�w>0	�M�:��I�mP�Hhm�ܻ� ���N�n�wH�	�&;`���&�w�/@��9�u_}�o��>�)P��!d&!&Fd�_�� 6]ߞ��==>�4�ʣM��U�/ڒ� �J��݋����������������]���Gm�b2�BrX�>��
�=�����זF.�l�-��v�� K���݋��әٲ��� �]��+b�CN�-��w.��>�|`I7@;�x����ҧJ��ѩ5�zGI&�t� ;����]sv�
��v�l�$�n�wH����w>0�]���*�;Ot�G��� ���I$�~��w���~~���4*JUU�h�5;s����W�m�Q++uU$��*�\t�Q؎2�uvHڥ�v4ooKa�v(�z���X�4�ώu��$�WF2���aKR�i�R�UӜ(�F��wO}Tvs����ն�6�ڟep������Ql�y�g>w�$�>+n�x�s]M�؃<����­mݲ��ۺN�:����JW�&sL�!zԈ�hGk֡#�r�����ɫ����ꇭp���^�7U�KwW1ֱruGsx��n��{=�v&���<����:M��8$����Bj���z�p�$�7@�� ;��?�]�\�F��k�Q2USX˻0�ڦ�7۵`g��lwr�U��m	����_�, �w<~�e`t��z�tLv�n����k ;�� ߽�X�&�_�,}�j���ڶ�;T$�'�����v���`N��ؘN��Nk,�
�S1�pE195X��m`%�f�{T�;��:G�u�]F��HM��ݧX�}�w��4)% BL�2HD�0��U�:��>��]Us�y��>����%��P�ҡ?ô�@��"��s���<N�tU�_Ji�mP�TҴ� w�� }���t��}~�`�L�jR)
�e�c�{��$�7@��"��s�>����]�:�Xi�K����l��v�fx�!� ���S�)���uʟq�T��g��J�[o���0��M�o�j�>����1��hT�Zot�H������<N�t���m1��,M5�}����}�}Z��$"�*$e�"*`��AO����;�,�i�+uwn����z���u,�>���~fwx�$���j�UP�ڰT�n��x�t��z�"�����w<k�@Xu	T�:�I�}�6�^8��gqSqV�$�m���Gq[#]���E�n�	�����, �w< ���OI7@�p.Ji�mP�T�SS`��_;;<@{�U���ـz<���'vԤ"�����{�<{���� }��}_/sh��_�
�i*&��^Գ �{T��ݫ�ݟ����%H��@�R�!��gwgk�bU`w�1�(�*	������tX��� o�� ��7@��8������8�jrd�6��Δ�y'f��"t�Kں�L���*l����K׈dT�Ѣ��X���}��	�t_�XHH�n�[��I5���ޑ��&��#������u�ۻj�Se�CM��&��G�}���}�V�Q�"��%��
��wgv���V�H���V$�`	�$�-Ӷ
�N�M�������	$���<�K���Am��m�Ћ����&]=�@�8�Z
Z�yh�\���kE۞(;[x�3����G�\A�1�'�v���r�i�&�vB\�yr�����nm�5��S��؛�핝��F0=!�4F����Ƹ���@�Z���x:v�@�s���ܖ;�x����gA�Lw9s���������z�����=�V��-x��ja^�g�����K�`f��@omT�VI]�nґ���ؓ�6ݲ՜n�����r�Nw�6��j4�HB-�/�	?��$�n�{�<�����6����E�t�i�I&��G�ws� =�s�'B�训��+v	���#�;���s�$�n�.�]��[����o�~���В�X�U`rIf y%V�:4ӺWO��I�/Y��<I&��� �]׀}u೪��[N�J�#X�^SnD3;��m�͛8�drb����I�ݧlm;���S�ƛ�$�7@=$x{��w<�u���v�B�
�� �J���gvg�(����=��I�n��p.J���S�m��ό ��� ��� �H�	Jʩ)Q$�1AD]���������ݘ��V�kK���j��"^�Z����KR����R���E�g�����+�t�%eN�I��ٰV���v���n�6g{7l���P=]&�3��wN�݂M�{���� o�� ������M1��v����]׀�s�$�7@=� ��41CS�4�L5���-K0�3]�f��ճ��R_v{�.�|�V�ݕh��7�OI7@=� ��u������gD[��	����tx��� 7��}$��wA��q�j]P�<:��!*F�4��n�9-f^���c�$P%-4OF�qU�c�B����S� 7��}$���G�w����RWJ�2� ��<�$� ��<ޏ���{��]��WV�o �I7@=� ����s�$�")�ӫ�e�ot�����}�Է�jx��!0xBa	Ad3$#xG��L� �#%`���D�V�LCI	R�5������kN��336n(�����i���QPk{0�L���3s��
w�����.� �c�+t4�;I��)׀�s�>�&��#�$갾,�w�H�������80fەK2��ݤ�X��:n0�Fk��Z�u���3����l{�<g�� ��x�y� �s�TDQ5IAQ5V/%������`{����۵i�����胺H�*(�&��&� 7{����+k ��ڰ1y,�:�д�.�]��m�}镀}����tޑ��%chr��f���� =���fv�{���h���~�U�W������"���`�*����T����Y��b��!Q@���B�(9* "Р*�����pߙ����hQU����������7����������������������������������������?����������U��g�����`�*�j����*����'������������a�������������w!�����w��?���(��w���@��k�J "� 
�%*% ��  ���C*$)"0����*HB��� H!*$� H$�*H@� @@$$��*�B���� ������*�B+(�(+ H! $!"$�(�����!*,�2�2H�@@��
���! 2#H H� �+ H#!� �! �! �H*!
B"���"�H�H@,�
��@!
���@�B+ @�(@�!( H"H��!����	 J
�"���"��0�����2���0�0�
������� �*�H J�( @$!  J2) B�B! J� HB2���0�
���B��(@��(�0�(�0�°�B�(B,�"��*�!��C D�`D�$F�BTd�$Q��e� $A��$dFRQ�$BRA��d	F��`eF�!A��`F��d`XA�	a@��@�@�@���	$B%%!`BY@�!P3�͚�O?��x ����ޏ�3�����?������ࠊ���������l����5�� ������g�}�_��("���U�r?�o�EU�����j���������_��rS��#?���c���曂���?�������DU��G��՟���Q�=~1EU�����U_�>�.�Qt��3.�������_=����?��U^���?������Z����~?� ���F��5���s3�/���������u?������e5���$]� ?�s2}p��fH)�TUHQ@H �JR
EIM4"A�RT�!
	
)�z P   @�PB
�(�I@
R��� B��$P�)@� �R�  QHUJ�    � @P *C >���n�#�b� i��o}�Ūz�:`��� �G   A���i\�D=�-Q��=�"���z�:>/��ݴ�c^N;��_|@@(   %!�@������6Y� s�� ��� �J ��((��P)��`R�3��J� �z�̠
#JP
 1 �`i@ހ�g�zR�: :\Ƃ���R�3e ����@� �R�OG@��ΊS� � H  
�w@΀)��
R�}��;���v�s:S�� `��}�ݯ<�jNov�ɪ�w�Ԫ���^����9�� ;��nWZ������@����O=ޛ�㻯n��4�{w�\��  ��罔�i���X��� ��R*��  UE����q�ͅ��o\�����W�� �+'����r�y%��|� �Jd޴�3� .0on.��<���Rǻ��w�u��R��v�< S�^�!�dc��\ ��J P ��cb��|صL�f����:[�ﱗ'�J��L��ϰ� Ӟ����S�� � �7�޺7� �;��!��[��o������ޏO�c�{��Ͼt��    =AM���� ��D�IT& CAǪ�AQ�4  '�T�h�z�`  ES�Д�U)JQ�  DSD5%I��0�҅�����(����>����T�:v��P�D%��w�DPUqUO򈠪����X���TU?y�#�^��
��Uk�HSe����|_9MYy/�'wm�'_��Pv_�QbW{{t���~��uj{�ex�@�
uR��@���H��@%4Ih��w���ͼ�g �p�0��ʐ����<�|l�<��>bH�	����dH1�!�I����b2$ؖHY>&��}iB�I�!$�!��_cI�Hb�b�W�`� �#�w߼�MهP�A��=��J�ww��������6H5B%A�$*I$�T$F"T"� ���Q�"�!8#��j����=���&��y�zmdYx�h6�UX�P��s�Nl��S��D'v_���� ʃ2��h�4@(�~��[hڏo}�'�e S����%�2�!$E{����H@�d�.�! D� ����cA��#b��Π�4�k�
 �DD\�v.���C�Bo|��9
h��HF$$P�7A��p�;k�\������
pٷ��r8xH,���WAcj5�@4p�� ��E@t� �ĸ�Y�l,h�!U��7|�N� ���=�	�����]�ُ��+$0�>�V/�X����x{�
������]����
�O�j�\8o���#���^n8=pGeT ��=�y��.��vD����H��,��B�w��4��G�ݙ�8�4���#Q�����A�9X ��@J(�IhQ�)�HXI�P� � �F�h���|�Qb�8�D�I���FH��$#JF@�$"0�Y�Op��O!Q����=D*�H�\wy~�UcE���-_�=�u(�xs7��,
h�h �A�� (��3����k������t���7P�n��-�8������<���mm��c*S�תQ�1xFk(�Ã��V��e�D4k{=�����xB;bG���|��d-XR�.��>v(x0
��$ �ti!H�b��J:0p=���3vk�z,L*���*ߺ�x=3��4l&��>�6[5�Sj�+5�ܱ���t�/����h4<0�L<�q��,�N�aMNy7�
y$.�q1l�-N�M5�wk�V��h��0�y̜�|֎<J�1(Ə���&���y)�%E�A�i�e��X�"@�=fĕ�&J�����#X�$H$H-u�����
B��B��
B��Á���D�h�,)��f<Y]lÆ�P�,,.���F�͘B�׋��.��HB��rӁ���t��0�B�x�ÉJM6Iy��ѐ��!� �X]�;!P�#,h�BA��$�jA�H$F�E�	 mUP�lh#A�6��w�+��2mv�KZ����҆X��@� ��@t� $�"B�.�F*@b���@�@bP�PP�u+,xz�
��т����w����JfY��s���Ɇ���6��J�@QK
�`�8�
�:^x]�%Q[9p���`� �kN�tR�A�<<	S��&#E����=�8l���Q���>Q1�ȱ�X� HS��p�9����OO �5��xxS֘$�Z�D���N%L�����6z��������&)���/�#�=����n��@؈���xA�7��u� Ѹ�LK�J�*�A݉^{Ģxl��Y����Im�2������!�,hں  Ļ�)�v����O��=TPr�co%�4�~�f���V' 
YB�X��)�P����$!�<{����7�xiD�*qT��Y�rzp�0��W[P�k�B!Q@`� �b^.B��0 �M�͞Ml�,,�98g��?�������`5�B�d�ULAxr����l3��y�M����=<)�\�$V0%%>vx�ͩ�B���.����I���u>�9��/������) �D K�&h���
r�c�@�����I�vތ�v�uD(��1�D �mf�^��$0�0

� �WP�E���6�` �E	f3������y���P+�@N����J�wuxP!&X#W�j�O��ە�����@u��բH���aH�7��5!�
i�d׬8q��LH,�$�sf�bm(E���j]���7~���7���߶��Y@�7�w~�zp*�D13������q�u����%&,+�3�`�J4	$� 
��
}�{zz�X��4�j�LW^$�
�Vnz���oS�F����h@�iF%@� �F��k�,aMS7z`��B@���C�M@�0�x��Ԧd.�SŗT��L���ٳ!vp�t�¡����&�\B�q;�R@I B-��H	��	��$	 �E
0$�B���ώk�7��xp��!bqB,]h@h�g^���v@�5�q�	�N1��*B.щDcM=4g	���g����j1h����E�L�4�&��!]\�o�(�A�%��wn.��Nhç�Q	�����TPr�����jǨ� �G��G%�ڢMɄaY�x$c	����)���4������R)���ћ1�#]l9�f��d��$Hȴ��%�H��M:cL<*Y.ɭg�������B����Ը�l�"Qd!X�$O<,E=�c$&����۲l��΍���:�ǣ*,L���A���%�����2Kq$6U�yX�ދ�Pb�Ky;9�#�<1�:0F�q�sN{&�!a�<2TA��1	y�2s2߭	nf�36�]8l�+����I(s�O� �A	 ��D��G$�뎨u�.�kz��xxJ�`E���1�2����S���%�!�V#�}��xc��>�3������#]���N��}OX<���! ��w�!/7�8|�%4İ_��]h$��)O�����l7p���ǃ�ą5�)���'���]�Y}!��0��
	rf�`+�p&0҄mm@ф�燃��~a��r@$	�T��@!M�Z/\~�4A��)~�rݛ�y�牂�n�lߚ�1��(����Ѡ��5�.� ��A�HH���S*�Ayyj���b��x4!w����@@m!�đ#M9B���A��$�,����A�91�d�4z���E� �5�0K�2�1�[�qk�	X����zK�٪h��_f˺�w�!2��¥�*{C��0a�L֏fؚ5ɪa��Gb@�
��z�r������ � �����0	���`�i5��8SZ�WMCLR��H"Q�
���Mq6m(��6��&�B0��0X�(]˼M�*{�H',�Ng�в�m�EY�`4!]�E�~(#Ρ
�`��*e�!&����b@�Ѷ6�t=��ٌ/8�ga�C,�k��[,�X�#	��$`2, bF (@>�}��=�.���ʳ��Q���L`�E��(��ϼ6k�<Z�c-ц�*F���B���(�LbWJB�O<���j�//�%�
hčv�lh��]H!"Jh�4Y�a��g)�#3r�ɨG  �N�m8 �����%�<(��y���œ���,+�{�g=�w��
h�w8x�d0���F@6J�B�//tu��y�&�<7��=<�Ĉ��VJi�3|&lY~�!�A
�u�^��(W��A�މ���>>u����H���xm�`�('<p�<��g��@��TPv"�~�� B~�����	�y3����! ������3B�Bʞ�@4��`�B5O8�/x��)��.�0�J�F��4!�#����^�(L��9�/UQ �B���Ŭ�V(�"<�(�%�/(1=�Z)1,g�>Z�4�Bd`�� ���	 ґ��h=|�!J��@����ʪA�/�{�9��L�;w�*	bƠ6h��:#i�`b��H��=4�k6D)ĲCDB'43[F��0�E"D�Me d�D�����m�ߤd]��!�\W�b5D�#M�	�_>��/�^<-��plP(4Q���w�����������~�:�o����    � [@  �    &���Y��n $)\m�\���Љp��f���mm���m��l�f� �ll��U&p�`jT�H m�]z^ݰ�d` ��%`ڷd�m���a ���L�m�ζ���ڶ 	 -�ֲ� 7m�� �m�am�$��� m� kʗ:� �mXaΒ�-�  )�m����&л�I�$6� ^���W��r�,����	äԝ,�J�m��V�6��   [@	
P6�                   	    ��+�>     �                  $   l            ��                    h        �>    -�      ?�>  ����                   8p                     ~�             l                >�o��ͷÀ ��m����݀A�-L���(k�gf��R�e���N��!�ŵ��6ۯ[�l-66ض� H   �F� rKh-�� �� �pm�m�d��ll�H� �H��{m��#GW�q��$�� �     H$�ֆt4�mSF��0X�7ki�v:B�o[W�4�j��u���4�6�z^�ધ���@��)�Lݰ�ƾi���H�m�n�g%�. �V��v�a -���p m�ϭ[��� ]��L�����҅������q��h浀 H'Y@%d�,�H�6����Ѷ\]p�ɭ`,2��!5�{u�N��On:;j��S�X[fZBnU(�)s�,@랳�.�<��np�a\�܍U����+�++q�\r���骶�����9��I�)ok�z�[R$��'95^h�  ��Kh[V� ��8p6�Vv��֦mUlv�5��$ոt.��R]�#
����eSPY�UUT�p�"%���٠A�Ŭ9�P)ݙ��ۢ#J����ZJ�/��ֹ�5��'�N[�����\Aڦ-�73��  $����Nځ7i�iҝl��c�t�h �l��^Yݔ��W��n�����ɥ���� m�$���Y���m�����0�$݅sm���r@mz��Z�`[pu���i鴘7n��m$�ݒ[�t�p Kv��qmky��%pl���r�ft9�_��u� m�ݜ/Xiv�'J�s��r�*��uѫIˢ6�m^�2�^@��a"��A��gaPoQۡN�:V�LVj��vvvyG5��TUR��i6�ڐ 
[oj�Ksl � �V�ɫm����m<�;�sa��{3�)�m���0;f�I$�����k�@�	��Gm� l��[���[K�UU*�\��A�HH�� .���1�Ēr[Bn�d�ܨ-3GP U��mƵ�P�X ��қ*�#�=����DR�u�C�K]WjyF M���iV����9L����q��M�r�"z�'``�����@:��<yVݹ]��RZ��B̫��E1��]�+uT@� ΍��1��t@  6ӴԷh*�Zl�$]����W(ݫ���������:H ��W�(UUR�8:B�q�m I'  �   ݝd��  H�2�p6٦���[@ �������M�i� ��ڥ�]  	��� -���m�@m�%���l ���   $�+[��p ���Z[:6�"[J��T�R�����U�[h [M�H-��l�� .z�[lN�v�u�K��s�`�p�z�Z��[tR�6�v�lHp˶� �dĽ��Ŷ�ɝ� WUV�m�ɢ	Pڥ@棂���uU��w�cc݀]hD����-+>j�7T�Q,HI��u�o�l�I�  �彰͵�� ��t�s�wU*k�7����Z�]Ѓ�ڹz��w;ca;$;u�]q�(��v�tn��޻��S���� 8m��d�9ċ�e�N�Dn�2�8�Y��ŷ� �R/j��<�ʲ�6�!pR�'6ʯ�����*�*��6�*�@^�;\&���k�J с� ��<������I�ܯl��i��M�-��h �]ԓ[[f�{ ������H[v�m� A���`5�W�Y�� -��Yp�H�&;Y�si�u��9���RI)�Ò �ŝ*ܒ�$�,��mNZID���pl��C�b[m��d-�i�q���2U@hێ�6�j�2Qب��/kq;yJH��K6u�rPm�˼[3����]���z�c���0�\x6�]˥	�:ۤZ�m�&-��-�n������u����  ���:2qf��/e[Kd����6�Upml9x�;t� (-�v�	ĺE��Kd��  I�����Ix�c�[jՠp��d2	���ul  6��ٵ�d�'M�i� �`  N�ȍ��f�l ���r��睕^[�sN�Q�j��s�ҭUTKp �Jආ�.��r�i.��6�oP �`4Y	6텶�,��h��:�X��N�
���8:�tf#Z@�]�Y=H�hͫ`rI9�n�]�p�m٢Ѝo[�K�3������M��{�[����cbVSl���fu��9~�?}ڪ�(��:��,t�Z�wGm$DX7Z�ܠ���G)�f���ǀ�W}����mqiF�燰U[Gj�;j�x� �`H�:ҁ����o 2�#@����e�)��6ͱ���a��&�t��U}���El�.����)V��Q�{*�Gh�%Z�(��(�5�֩�vsAJ��)l>�}���x� iӴ� �e�L�Z턀]W�  6����V�T���G$�t,RFճNP8  [F�:l���4�;$��u�0Ӄm�ZǧYF�	 m� [N] (]U�h1p媪B�-�� sm�l m� �o�  �����0[K�v�-�  h ڻie	�V�j��K%H���&פ�,� m[	b5��BA����a 5�pWUUJ�
�J���T� )[m Mm��L�X �l4Si׋c\�O��|6�Hm���$�XK���"��ٺR�oe6��m��7m� ]�&׷`�@X�Qݜ� �UD���]���� s��f�3熎5&��,8hVMۊآ76��FC���h�v���[v�\`!��Nm��4l;��8����-�l��M��w;e��z�ۥ�c�V�R���үe�|�祷W2!�`�CC�G7�,"dWv��$pD�K��  � ֽ�/����3l;
�@�m��7BMJ����7ѱ3�fGF`��tF� ��m��&e��a�jӬK��   �i��A-MD�mV�    �4f�S���unYYV��z�b�evq��U����t\�t����n��m�$�  ��Kzܖޗ��Չ2�F�iZ���ݱ��A����Tv�L㗍�df �v�<	�7L�(E��m�V�e�8�+�"�J멶��s���٤rM�J[�8Y�ݷBjzղ��rgMNR(�#GI��Ԓ8I��H춀��F��-�m�D����T����P��6�����m��K(:�[p��-��zt�M�Y�쓆�&�鴇��{(���ЪΥX
�j��&�V��	]��j��
U��ږ6�p3�lIe �XY�&��5���  km��Ŵ]*�/[mh @l#��Y�j�]���=!m����m��  7l�Y�  ���p	4Qm  IҶ m�  � f�[i�I��1� ��m��xEj�8   �8  	   pm�6m؍��"[�� �    m�$�   [F����ݰa�����h��̸  ����z�&�n�� 8 $  m��O���� n�t�J�k�m�     ��u��[#Fն��C�m��]�Ya"�.���$��%��e06�ְ � ^E�[@,2S�KWg[y�®��Ë�C�p{'o2j��=�`X�M���k�������[�^�o\���(�+��p�l��l��.��U@\s�u̗�t-�̗-T��v�5��AU�l��ꖪ��Wi;ם��a��.��]��mM�����^j
@��(�-�,�X�Wd���m�s6{=�wQ����o��� 4����f���]�%�I�j:��Y}�-Mb��M�������
6
�FVV�n�eZ�P����
�Π2M�  ���{��w��T�"" ����v�� ���$X�R
�T�*��?��?q/�������z�D݌(UA6+�D�Aڧ�!ꉠ�b���SWF�$�!"ĂE�$"�I#0�aF0�>]��DR*U_R���� DVEG�`�����B������}E����$BE! �0d! �A��#BB�X)�FA ����� ࢿ"�@p�DD���T�� `��V�Eq �B�.��D<t����E�t��B>�+�HBX0@�����v�> ���
�"EB� ��@� /� x)Au,ĉҼ�8�!�S��<UCЈ�/@��|��!��Q�=���D���",W`����Q*D
�x	EE� 6��� ��S�T�P8	�:A�F#�����L b*����'��W`��)An�S�T�P�C���&�ث�Z  ��:������AU���H
(1TH�w�_��i&��{k�m�n�d��K9�vΉ�dq��I�]�V
��ͦy^�pv6���kc�p�{m�l   H��    l �(   ���m�m��   �l   6� �`H   ��Z��5��������X֌ie��H�0"`imUR-A�� =;M2n9X0�͐�fv� �:��Xz�v�gPJ������7a�{.�^�u�OiK��ܭ�k ú��\\Qp\2�r6�ݪ9�r��p(8]8�N���GcK�:Fk%ï���d�e�[N��69I���7]�2;���m]\�m]Yy�b�Y%�Gs�;��S͎���d�I�3��,�V��L]����Mm�x�{\#�;sH��nQpDT�� U�۳���g6 �%�f�:)5�;*�u�Y2�T+��Vǂݬv%^(ȳ�W�ޓ�!8�n��ӳ,-���!�M\\Ml��]u�v�N�s�ZTM��Îr��6��1��5ʑ�ix�a��y`˸���'F6�uɷeԓ������콯[�Nt�����h�ϛ�^%Ú�d�6ˊ\Һ3F�8��C���q����pr��L�B.���A4��;M�[��[�Yx�''km׳�6�	v����L�n��C˴�pLU��x�'�j�]-T��g4r�c�n�,��ѹsM@uUc�t����[��K��bک24l��������'����˸!�y8�Ս�ۭ.ܭ�Sm�����:��jӻA7nم����/F�C@)���_.�x�X�/�n����ռ�rvҬ��=s�dʓ�]��a���m������Sv�m�GL�ter��ԑ�"���/k'	�ě7e��c�+���Y���Ͷջv�0��Ӂ�vi 4w[/
�r���X	<Rku��!�;UuWe9�����nl[�Ti1g7l��]\�m��=��.��x�vhru�[R�*���!j�.�n�k&f�\ֳ�q��
��ڡ���ȧʄ�hMl (? �U���'�Z�5���4�.|5t�K;m��Ci�U����ι̜*�\p���#ɓVn��<t�8-�c�簲\0�td�;��7n��G��cm�r8��ۛ	6�D�+f��[l�m�]s��Z�wh���S����ͭ���ۈ%�Ѩ�eɼ�OF����u5ڪ��z�k�6��ᨷ.�j�S�t��g�!��� p�ɵ۩Rt;V���{��u��f7��+݌��M�"m��ra㷲�{l��vܽ��?���c`6�m��'���^� ���=�Jh^�uł�bq��M��
�W�r�T�zS@�v�ʬG;�#Ps&8�^ꞁoJh��@��z�v���)�D�zS@��ZW��*�T��,�'`�H��p�/;V�U��
��=ޔ�=N��r7�4��*F�;���v�Ъ
���v80���ݥ�=�vhF�=I���m�����{�z�)�^v��P�d�Ҍ�b2Gd�^�N�U 2���(�Y)�^v������X�c�R��U��� ��0�����=������= �KA��Q�ԐI�@��ZW��*�T�zS@��c�,J)�F%#mŠUz��uO@��4�ՠu�q�X�`<��+:c �ݸ���9��ϣm���	��wC��r�i8#��152`ӏ@��W�[Қ�h^�@�Z��Lr`%##RB=ޔ�>�ՠUz����@�R	�v�$���@��V�U��D&�GЦ��>� �� ��ӑ&#h��	���
����vI�~voY�}]�@���:�1�Ly�#�9{��޳@��V�w��~��ݝ'�� xM7Y*��f�f����;�d��u�Ty��# �i)�Ng���HG�^�@��V�w�����@3�Z5"n(�cn=��� �u�.� ����ݎ��QLRPM�U]� o5���:ñ�N���=���@�������ɌrM��� ��Z�aDBDD$"!B�^�h]V5H�?�H�$C�@/u���� ��h�[4\����)�6���n �āӞM�Ux�n�ql���ù���kZ�5��y�Z}l�x�4�Y�ܚvD�FА�H��٠�l��f��>�@���:�1�&?�2I&�{ų@/u���� ��h{�V2D�8�ds#c�@/u���� ��h�[4>���R&�F�j� ��]`I(�������� =ޖI�(4)�>��	�$[���ێ�]p�I�6۶�I���7n���q:)���g���}��nuU[vH��ʇ1\�1��\D�*u��ևc��Өp�0r��B7=<�&0�y�>λn��n�\��;-b7�����d�����;b1LkOd6y�"�������мGiR���ݫ�7��2ۂ�lJ=�N��<�/Om��g`���9��s<��P��B����ȔmF�h[}�Fkv{S�&x"ǋ�ɰ����;���Dns�x#A�,S�$NG��u��� ��h^��\��,�MA̙E]� s�w��	)��}�g_k ���U�X���d�㍎M ��h^���٠�l�/�A1+"��$O����� ��h�[4�Y�ܚvA86б�#��f�{ų@/u���� �%� z�i�p'6z�NJ�Zy#�׵"�^H@�����ul\�i.�$�2��7;x)~�Oϋf�^�4/uz�h{�V1�`q�c�6\�I=���� h�(	`XA�F@�B#.�Q0�T$�&w`ݳ 9�����\N
F�QH�NM��^�ץ4ު� ��h��,S��)#�:���{�Y�z�����,G;�#$s1�h�U���W��>����ץ4���:��#z�����з��i�ۯ]!����{o��m�e��z�u�BW���JW�m���~_��^�ץ4ު���Ĭ�s3%����<�Y؈S#뾘������@=ܚvA86б�#�8�ـ�x\$�� �%v:�o ����Pu�Lm�G ���@;�����ץ4�ѫP&8��H���l�9{��=zS@�z���e��(�l�Sm9!���5���ֲ>Ӷ]ٶ�:NQ���v;I�tO����I�'Mɠr�W�z�����UV"Oo�K$����
��I���)�|�J��l�9{��<�b9�Pi$��9��W��f���^��Қ�U�Xړ��L�(��w��/uz�Jh?f�a �!T y�vI�jD����$��$�@��@��M��W��f�ה�q2&�@�@Y#���5�	�9�`�v��]r���㰽x��L��5a��Hs��^��>^�z޶h���PuULM�G��W��f���^��Қ��Ս��1��Na##���@��@��M��W�}JǑF)��#Mɡ��R�_k ޻�}<c��Je�{xW�?�,$X����>�@�z��޶h��������q�Cq���igmjj�@keZ��b��l�ꖲ�W:��F��Ƞ���d�lF���[�����v��WO09^Ϟ��%���O���%Lv��uk��8xe�4d�p�x���D�r����ֻcDRdn�X��`�p�71l0�����T��;ڋ=v�&1r\☶R��l7��ٽ���!o�Р������Qn��͔�[b�:�Գd��ֵ2�7;��uڷh���^ll&���u]x�����Gͽ�8�qd�&㦣���?������������}V���cV1��G�9!�}�f����H���w;�h/R��rA1W#��$O�$�/uz���?%�ߏ�@=߿M �ri���I`9���]��Z��_��}�f���^��P����1�H�q[I,���1$�[>�LI%�{瘒[���> ?���Θ^�Q!�B�p�e����7[zvԎv�f��[^n�xYJS����ƣ�I#�ܥ����瘒[��+I%����$���,EP�7��Z���=[DP �j�Ѡ% �G����N\�H��)i$��� QRq��1$�_XV�K=9s�I#�e����瘒Z���h(���ZI,���1$��q��K_��bIn���$���te�F8�q�y�$}ӌ��[鼳Ku��i$�����I+jS4�q(d(dBD{-���ڃ/���p���nO\�-:��@mq�HʎC-$��o,Ē�}aZI/�*��H����I{�4�pm����"�I-�����N\�H��i$��yf|*�6��K���P&�CRi$�����I#�e��^`�.��f��"��3Z��ze6Zh ��J�DX�Rf�K�)	�kD�<NS�F�v���.�$P��d��]ш`m@��K���֑i��V�Vh̈́��-ڮ�%��	� D�� �XP��P�P�e%%�%aH��`�".��j� ���-���itѪh�ՓXˠ�)��	H\
�b�3@f�]�ںB`r7WZ4�ք�i�B�tgE.�ٳ��#,�)4ի�ĊLt](ib�My4���a��I�X]].�5�B9��!��n��d�)�sZP��.���P� M����!
ӗ1�H+VԦ����4h�ֵ�K��� B��@JJ
���5�nPO<���]2���� R���c Lm�aw�MW])@��'���E�R��1QqQ�>
����� �� uP(��z
���U@z�˛�1$������m�q� ���N�Q�$��N2�Io���I-�����N\�H�zy�"��F��ZI-��Y�%��´�Y�˞bIt�-$��xD�AanAG������h�L�s�e7]E�γ�[�T�Ӭ�:�@��$��H�Ku��i$�ӗ<Ē>��}U@m%�;嘒\���!�F8�V�K=9s�I#�e���M嘒[��+�
m���L��.J1�$�ȣ�I#�O���[鼳Ku��i$�ӗ<Ē�ԉ�s�A"IRH����M嘒[��+I%����$�zd��"� B
H�	�E*6�A|U�y��7m�﹕��I�\GbIn���$�W���H�MI%�N7RH��M�"��S������v=��[lC&0m�:�<���ݍt�>�#8������> ?_��<Ē>}�ZI/n��� ��]��
�I{��!"p�1$��r��K۷�1$�_XV�K:r瘒DW�cȣ#�n)�$�ݴ���}aZI,�˞bI>�-$�����I�HRC$�1$���;I%�9s�I#Ϫ��K��O�I.M#�ő��i'�IgN\�K�(��SIo}����|׿oSv�|0�Ű Ą$$VIIT��s�5Z١i��+s�Eܕ*Ɖ�\��n`��1�kvctIU���؛;[����-r���LIƜ>��^Y)���r��뭻�;[���p���q�@X3����{�<ݗ��v�[�,l�\�Y�R��]�U�`��4!�u��v��vyv� �����=��vb͛�^vN���*Ź��H��b8к�N�J���#" [J(�1	�ڠUP���m%md�pf����`
�V�[[�.�N�v䓁����z��stP�*�{L�*Ey$���;I%��㘒^{�ͤ�Μ��$��$L��	HʒH�$��o�bIy�[6�K:r瘊G�yKI$���}!N�H�"�Ē�ް�$��U_�$���MI%���$��8�W(FR2��IgN\�H��)i$��|sK�zô�Y�o�e p����y�$|����_�U�Ϗ��Z���IgN\�I-Kz�HH�� �.�ѧDk��0�Q�m�d v:Ů}��l��ݨΚf2�Q�ɌȓqKI%��㘒^[���Μ��$���R�Ik���S���IbIyoXw��%U@�� R�iT�$ZARą(�Z��Eh����H�B�U]��|��H��^ݾ9� ;ܩ�!��;�KӳW? ���>y�$|����^ݾ9�%�a�I.{Ï�潦J���~�����~K�{�㘒^[���Μ��$��$L��	J"$�KI%��㘒^[���Μ��$���R�Io��m㑱#h��V�mý�ݵrm�	�˖��7�� j�%��=�)F�6T8n�����?��s�I,�˞bI=�-$��o�bI{�qW(Q!����Yӗ<Ϫ�m���MI%����Kˮ�Ԓ_^�\b ���N#Q�$���2�I{v��&�lTZ)�_/�l����{~�9jDk�̱f2c2$�2�_UP����$���ô�Yӗ<ėª�޿���\�|� IpĄ�$9�%�a�I,�˞bIl�-$��o�bIs���/l�mvz�n']f��a�^u{o>��6���"sqsst�i5��y�C^i0��I,�˞bIl�-$��o�bIyoXv�K��es��F8ԑ'Y�$}����^ݾ9�%�a�I,��1$�� ���L�	DdrRI{�i��%��q�I/��W�$��KϹ��p��	�p�$����i$���,Ē>��ZK�
m�Ē�%�Y\�E�Hː;I%�ֹf$���2�I{�i��%��q�I%�J����Q~�زU��Ûs��=�q��+'���0Ͱ�i�ƺ�͆�����/�|�K۷�1$���;I%�ֹf$���h���̉'��^ݾ9�B�mj�;I%ﾵ��I#�e�T6������K�$$��!�I-]��i$���,��U�ޟEi$���9�%��u�B��Hͤ���\�I{gEd9�l��%	N��� �ʩ�ګ�.����Z{�4wJh^������0U
�wY<�%�Lq���@�h���v��$Z �[p��<s�����*�+���������v��,cu�f{���5���)�swF靻b�x�<�C`3�b���۲`y[k�rWG8a����*�]]�E�vGקu��`89����*�����ܼ�7�c^ΆM��T�;����w%��9��L㤻F��X��B�8�J��;ٯl�ە��h������zy�?4�Nv7�6R�m�;��g�N��wa5�d��@{Wa��mqU]"#��/Y��>�w4����Қ�si�pM��̍�h^����V���M�Қ�!���!���s�.VI�l�g�P��[?�_ۚף�3ɋ#�s��@�t����M��s@�ت�;9�M�(�0��$�{�S@����>�*��Jh��,I)HbQؠݞ��@x#��� �u�s�x�F&؝&8ic�2D���BI��s@��ՠw�S@�t����:�d�!��3�>����}�"�$���B"HƁiQXQ�(�V, �TE(����_~���>�����]� �,���9�NH��-������;
�:�� ��변}.d.+$�$@�dr��4�]���V���M˹�쉸�hc�#p�>�w4�Z{�4wJh���l�_1�k��l�F��.�xc��l��]��7��V.�H�r�1�S�u�$�ɚ����Қ��4�]�$�l|�!A��(�N�g��Q2kw� �_q`����k\�P\c�FH�p�=�)�}z�i1fg�̠�
�{�+$�vq�N�	%�"RHI!�}z�h�:��Jh��=ZG;�&8���I3@����;
!�Ο��L��U�i�s=���q�Y�-킶�����ݰ�t�˸�Ճ�[�(ɷ9:"�n0��Y��w�S@�t���빠_X��>U ���L�(����M��s@��ՠw�S@��m;"n$��Hݘ�^,^ܹ������`�}0�T@B��dŌ��3C�+�����gf�}�}7&�v 5`�(� �1��H2�7{�}7���q��LY$���QE�w�S@�߮�>߯���EV�Ue��(�hc"�B]��5�������v�˹�v�NQ��a���D����O»WN˨߭����t�>z�`���R�A뾘e��긐8dJI	$4�]����e������Jo�H��"��Ɏ"d&(L�/��w�S@�Қ׮�{�UT��'$�����W��4��L��Ы�]�����]�ڻR��]]���`������w˷� �m� P��Zʻ�LB���,�|�Y`)�CSo<�.`SXm�٭��݆���a�t������D��^C��a<��cR�A���she8D���4��o0CbEbF����	P��aO	tF�i�H�4
�����h��3Fm�5��@�ɣёcBjR7��NGG�^h�5�&y�!7�ˡCO$���R��.�IH��of�o5�8(m2)�0߃ȜZ%�]S=TA��,1E�f-�������k|����I�Y��6J!&���xF�5��c��ItM�+�$�|�||ׇyR0��&�]f����������f�ZK.��ܹ�'�4&�)�TS��)���z��P8��?�А�$�d�Һ�eV�Q�9�6�Bv���f ����#d�ҨK<.ln�rV�I�q���   $հ  �   ޠ       n�   6�    ���  [-V��"�e��\M:#C� %R�cLs,�3�����'Q(K���\=��C��;OU�ͻnUL{1�7_�W��z���5tK�.l��՛=��oe�-���vK��F+E�=&y��h(��aN�v�nӶ'-��y%��ݳ�˹���I�񾛾��&uf⡺�&�Ν��rS���b�.� v�Gq���J�X 8
���"���a�.:���T�� 2s��9+�YNV��v���#k�Tu��<�z�md��x�֋�V�Y&�8������ǅ\=���J�����k��;�������U�����8�1<�v��XRk���O�S�����\�]	'L���h��e;�`}q�n3L�۷)���C;����uu@���-�e济vܒ):N��ӫVD�݌=������,�ݩ�-�p@�����J�ơ�ֶ�Z��!�4�[���n7�ci;3Q쒘6��T#t�nu]3��9ڠ|�3���B�cG]��Y:�S��a���ʁo���Kr��4�T������6�d��XF��ɼ�
��U�^xӍ�7Wm��Ge���셓r�ql�u;�\MGB�dZ�'K�GWc/������ݸ��Ɣ�೓K��G���|��f�B}n�+ێ}���cq4ʺ���!I�������Pn�Nڙ��:l�v���,�\��WvgE�]�iმ�ɽp��w\lj��v����f�n�t[$mcI� I�^lZ�� ���]��L
�%^{2UPm�R�lI���$.��2�e蚭�,L7i�Y�݋w`f�ˋ�m�d���LXP�ͱ�^rF��U���V�c/q̅���n��
]������ڶ�R߯{���{�{��^�� �P�`����GP�Ңz�ӊ�����~��luj��W���"~��f�- [{m��lUR�粷<���a�iJ�����爞��b����m�b��<�̓3q9w<t5����p��]Y��cg(]��"�90�[��۞�{r�Z� pg��=;��fW��p��'g�v$�Y�N9���<��v����͇Wk����<���o[�v�خ2r�y��Y7 ܄8��5�)Ւ��6 U	��jl��u�e��%39n-�Dm��6�n����GK��8��ѻ;Z%�wu�m�r&�I���F��O����$��`Ͷu/�]��9��,$�ͩ�jUuUf�m�;
dz� ������s�>q���	 nT
Cd���`�هaL��`��LxmӚ��tE��՘IK�Θ:��m����y� ��uWU��U����.�����'���=w� ׶��-�fF��C�$$dN8����������:���lX�2�b~.�#.#0�������S���m�K����b}߷ٴ�Kı<����r%�b#Ao!��@Ԁ��B���4��X�{��6��iګ���,�$DjBFEu.�
T��4B-��$ND�;����r%�bX����m9ı,O�}�ͧ""�F�4���D���A B0Dr����bX�����ND�,K���ͧ"X�bX�t�}�ND�,K�~�fӛ�oq���~?��� ��m���,K���ͧ"X�%��O�ٴ�Kı>���m9ı�>����r%�bX�t훒��ԸaML�kY6��bX�'�>�fӑ,K��߷ٴ�Kı>����r%�bX����t0�F�4�缗�8�6�i���`l����ѽw�X���;/W�� �*����P@��7*!�h#Bı>���m9ı,O���6��bX�'���6� ��5ı;��x�_��$)!u����P]��Us7Y6��bX�'��}�NAVı,O;�xm9ı,O�}�ͧ"X�%���o�iȖ%�bw]:k�e�k!2�k&fd�r%�bX�w���r%�bX�t�}�ND��z�>E0Q��G����*���@��5q3����Kı?}���ND�,K�����$�&\�36��bY�
AQ;��?M�"X�%�߻��iȖ%�b}߷ٴ�K��@[���M�$R{�;{p��$���̔�dؒ	"{�bn	 )����iؖ%�by߻ͧ"X�%��O�ٴ�Kı=��{���cn-�8��";#k�0�h�nm�y��3�9�Εڱ�im��:�t3Y�iȖ%�b}߷ٴ�Kı<���ӑ,K�����ځȖ%����A�F�?����7M;��fk&ӑ,K�����N@Kı>���6��bX�'�}�ͧ"X�%��~�fӑı,O>>�rY{��E535�ͧ"X�%��~�uv��bX�'�}�ͧ"X�j&�{���6��bX�'����ND�,K���w3T�aL�5�r�j�9ĳ�5����ӑ,K���w�m9ı,O>�y��K���
B�"B(��(�� �X����]�"YA�����M�d
Ð4�h"�%��~�fӑ,K�� }���O"X�%�����]�"X�%���o�iȖ%�bw^��nB��k#l��xn��\�'e��{vs먶�n�tT���]�ss����2Hn��F�4=�}���Kı>���ӑ,K���ٱND�,K���ͧ"X�%���w%.&��[u�ӑ,K���o��NDı=���m9ı,O;��6��bX�'�w�6��%�b-�>_(���HS�����4��{����r%�bX�w���Kı<����Kı>�w�]�"X�%�{퓶w3Y�n�%��6��bY�@(�'��~��r%�bX����ND�,K��}��r%�b���o��a��h#C��m?�M��M3�CiȖ%�by�{�iȖ%�b��{���9ı,O~�}�ND�,K���6��bX�'����/����\ɚT�۫T�t�`���86��I��ͶR�I	4x�N�&���뭱�*�%�N���]�z��U��_ ڳyٱ=��7�b�'j����g��dU*�ظ�+<��6{&YE��5�nּ�1�3p�zi��:�)��<v����]���W���cl��vZ+���Aj����$@\��֍H�2�7���ѧ�<-h��LZ��%7L����v�=^��p�A�q��u�p]<ϹwF���d�aML�k0�>�bX�'������r%�bX����6��bX�'��xl?� yQ,K����iȖ%4�߾��F��$��QH���A%���o�i�
�%�by���ӑ,K�����ӑ,K����uv��F�4��o��&@�,In���ı<�{�iȖ%�by�{�iȖ?�����L����ڻND�,K��o�m9ı,N�Ӧ�k,�Y��S.a��K���WQ=���ND�,K��o��ӑ,K���ٴ�K����O~���Kı?~�{��L2L�e̶�ND�,K��}��r%�bX����6��bX�'��xm9ı,O>�xm9ı,{���?����V�Ϯ��-�c��B����3�'}�rI��B�D������z��qYj@KrG!NF����F�4>�����%�by���ӑ,K�������A"j%�bw�����r%�bX��"#�GF$%)!�h#A��{�NC�Z+��6&�X�o}��Kı>�w{v��bX�'�}�ͧ"�Pꃑ2%��~֮��+f"[."�p�4��hw���C
X�%��{���9��Q���j'���M�"X�%������ND�,KϏ��f�s%�
��a��Kı;�w�]�"X�%���o�iȖ%�bw��fӑ,K�A�O{���ӑ��h}�[�#AA@ܨ�j�a�ı,O��}�ND�,K� ?�~���%�bX�����ӑ,K���uv��bX�%�����ZfY�	fN�R2Z�ZX;6�t��&�wg��us�{m��6���2�p�F[��a��h#C﾿�ӑ,K����"X�%��{���?A�&�X�'{���ND�,Jh~}��#�$\ �"����Aб<�{�i��-��,O��o�WiȖ%�b~���iȖ%�bw��fӑ,K���/�2ɆI��\�na��Kı;�w�]�"X�%���o�iȖ;���_�.
��j&~���iȖ%�b}���m9ı,���9}j@K�E!NF���G�����D�����iȖ%�bo�m9ı,O;���r%�`
�B��ީ�_��$)!O�����]Z�)�$��6��bX�'{��m9ı,?�(�����i�Kı?}��v��bX�'�}�ͧ"X�%�ߤ����iz����h�N�㶮N��xymcz�lmu̓�����2�U����&�FkSYf���i�Kı=����"X�%��{���9ı,O��}�ND�,K��xm9ı,O:|n�5{�.W4f��"X�%��{���9� `���b}�w��r%�bX��~��iȖ%�by�{�iȟ���3Aw��H�P@��7*)�h#E�b}�~�v��bX�'{���r%�bX�����r%�bX����ӑ,��h{�[�6�p�@���a��X�X��{�iȖ%�b{�{�iȖ%�bw�ﺻND�,�S��Kt�(�0 �$b��B���E�'lN�?r�9ı��������d�CCh#E����"X�%��{���9ı,O}���9ı,N����K�q�ߏ�����l�mvz��^n���,�c���s���v��3˥u_H��Sg/����bę��̶��"X�%��{���9ı,O}���9ı,N���D�,K�{�ND�,K��}{��R[�9
qEt0�F�4��>�]��B:���'����iȖ%�b}���6��bX�'}��nӑ?$�MJ�_�/�����G��A
%���p�r%�bX�����r%����������9ı,O��߮ӑ)��hk��o�f"�N"Ӑ]4,K�{�ND�,K��w�iȖ%�b{�w�iȖ%��'{�xm9ı,O}>7e��̗+�3Y�ӑ,K�����r%�bX�����r%�bX�����Kı=����Kı"cb��,H�)�d�V�jEH�@��$T�_7��K�a�n�]��t��$�����Ͷ<sӑ�.^Amq�Ӹ�n�{=:����]�w�va��\��]�i�u�D�l��we�[�ظv�:��dW���g>�I{F�û���j�j���f@�]�؃qF�璝]�u��m�\�NA&���e�z4cG�d�7�g���P�.x�֍�>��q���D/�N��	�{[#jy�i �:N#i�@��͒��&�9�9[Q��7(�����0Ͳ���{��n�h( BH�Q]�F�)�����r%�bX�����Kı=����Kı;�w{v��bX�����p$�)��A�Q;߻�i�#uQ,O����ӑ,K������iȖ%�b{�w�i��QD*!I�w��U���7w5fk�"X�%��߿p�r%�bX�����ND�,K�s��ND�,K���6��bX�'��w%�fL�rL�n��r%�g���9���_��Kı;����ND�,K���6��bX� �]D��߼6��bX�P\��ˎ\�)
qEt0�F�4,O}���9ı,N����r%�bX�����r%�bX�����ND�,x������Hiz��(n�l��E�2t����ʎ���l1"`q �*8
h]
�"�c�����
G��h#C��`��Kı=����Kı;�w{v��bX�'��{v��bX�'����H�1�q���a��h#Cw��r:cA>+�R(VC����	0�`���-���T���:���֑�.�*"xP=|O��2%�����v��bX�'��߮ӑ,K��~�� �H�Hj&�X�|tݖj�̗+�3Y�ӑ,K������iȖ%�b{�w�iȖ?��D�O߻��ӑ,K���߸m9�#A�}�H�PD��Q���A��D�����}��~�ND�,K����ӑ,K�����ӑ,K�j'~����9ı,Ozwg�Mf���k0�2�9ı,O��xm9ı,�	 b }���O"X�%�߿n��ND�,K�s��ND�.����c�JH��(�c�8��$��W��yܼ$�<��)F8LZ�u�9	��Ff��r%�bX�����r%�bX�{��ݧ"X�%���݋���"�MD�,N���ND�,K(k��߄F#R0dI8.��F�)�����r+�����b}�~�v��bX�'w��"X�%����"��h-<y}Q���E!N(��D�,K�s��ND�,K���ND��p�#`��� �00t�����z�y�)�p؛�@�O9��b��À�4�Ѭ�p�t.`\��tʚ��<�ּ��<4n�tl�Iu��������&�>��D�Z�k����kD����RX�{��
�ٶki�%%'5X�M �P!A"SN;H]b˦]�BXm�śf�ݦ��p^62��j]��(0B`����
����LC�O@��	tiiC��0���>t�Ip&h!� �#���֎'��9�Le�)f&�ӿTSV���tDK5��c�f�5���K.�U�]��d֣�3H�RTb@�a��!�
|���&�P3(��'�.�up }Q��(��>���@�)�0M �_ʤ��L�p�r%�bX��۽�ND�,K���[;���L,����]�"X�~T������Kı>���ND�,K�{�۴�K�����nӑ,K��]�Zֻ���E��D��h#A����C%�b}�w{v��bX�'��ݻND�,K���ͧ"X�%��~�}�kB��[]�R�ӳEӎ���ݍg����t���[�V��p#��ޟ�0�ӈ�;t��m9ı,O���nӑ,K�����iȖ%�b}߷ٰ���"j%�b{���6��bX�'�߮�\��\2��5�f\�ND�,K�s�ݧ"X�%��~�fӑ,K�����ӑ,K������9lK���흹d�j�	��	u�iȖ%�b}߷ٴ�Kı<����Kı>����ND�,K�s�ݧ"X�%��O��5�L$�ff]��iȖ%������"X�%������r%�bX���v�9İ+��aB ��X ����5��iȖ%�b}�l��D��B܉)��A�F�o־[ND�,K}ϻv��bX�'��}�ND�,K�{�ND�,K��+a�~Q3
�d ���eHC![\��Y�y:w;�8�u��cM�v߯{��J.ə��2]e˴�%�bX�}��v��bX�'��}�ND�,K�{�ND�,K�{�۴�Kı/}�ճ�����ɘ\�˴�Kı>����r(ؖ%����"X�%������r%�bX���v�9ı,Ouߵ�k�(�E��D��h#A������,K������9�K�����iȖ%�b}߷ٴ�Kı<��Қ_FTQH�G �h#A����nӑ,K�����iȖ%�b}߷ٴ�K�[�{�ND�,K���n\�.Mf�3.]�"X�%���nӑ,K���o�iȖ%�by�{�iȖ%�b}�w{v��bX�'�U$GI
yM	 w㣿��dZbz����i�$Z �n�a&� ��H"������<u��K�Q�3(��i�m����k&�ۮ�֋��<��*m#�'&Ën��Y�o4�p�f�!�n�<�<<���Nm��k�db�0\�;Z6�v:����Y��vU�agY��ݍ��:[�j�c���;�&��V��i{$�����cv�vx���ב+�X}�����w���*��ӐVb.�ۚ���|k�f�M�۳���i�
�F�'��{���]�26Ѭ�.��=�bX�'���ӑ,K�����ӑ,K������?��MD�����r�)!I
H^��<����feљ�6��bX�'���6��-�bX�{��ݧ"X�%���nӑ,K���o�iȟ� �j%���Y��Y0�u�K��na��Kı;����iȖ%�b{�}۴�Kı>����r%�bX�{���r%�bX�O�D�f$�B�Q]4���
5H�������Kı;���6��bX�'���6��bX�'��w�iȖ!�_oŤ~���� RH����b}߷ٴ�Kİ��@"@A��߼6�D�,K�~��v��bX�hn��]4��h}�+g�\E6��{tmOa��u붹�Nm�m�X�#�fxy�؛��YVb4dF6V�{�[�ou�by߻�iȖ%�b}�w{v��bX�'��ݻDS�_"j%�b���2�)!I
HZ��ML��f˒�f���ӑ,K������9
��D��	,(��RM�th <dMD�5�w��r%�bX�w��6��bX�'���6���?�*0�dL�b~����sT�e5��ɬ�r%�bX�����ӑ,K����iȖ?D�Ow��"X�%��ߧ�m9ı,O=>�ۚ�rkY&�-�]�"X�@?*�����W"~���&��	����A$O<�}��$���s�ݧ"X�%����m�I���0��a��h#C�}�ND�,K�
��~���yı,N���v��bX�'���6��eh#A��P�	2)�:^z5� %�<vv�r��=m���M��?}��a�鍣%�5��K�q<�bX�'~�?siȖ%�b}�}۴�Kı>����Kı<����Kı/��>�M6dRF�)�.��F�4;g|��D�,K���ND�,K���ND�,K�{;ͧ  ؖ%�{��V��[�L,���̻ND�,K���ND�,K���ND��	����{��ݧ"X�%����nӑ��hk��o�d&"�N�]4X��"�'����iȖ%�bw�ۿ�ӑ,K�����iȖ%�b}�{��a��h#C�֊i}R4�"0��ӑ,K������9ı, �ϻv��bX�'���6��bX�'��]4��h|��/�q6$m�d��.�.-������]�`�O�]�ܩ��C'G5պ�>�~����{��{�v�9ı,O��xm9ı,O;�xm�Kı=����ND�,��h�(�P�	�Fq]4��X�{���r%�bX�w���r%�bX����ݧ"X�%����nӐT)��h{�y��Rd�$L8�h(�%��~��"X�%�����r%�bX�{�v�9ı,O��xm9�F�����D�
pB܌���E�b�X����ݧ"X�%����nӑ,K�����ӑ,K !*B(� b9�<����Dh#A���дْ9��WC%�b}�}۴�KıP~����Kı<����Kı=����ND�,K��oNL�5�e���� Fc�l����d܁���<�a)9Ǯ��c�@��Q8��"��)$WCh#A�}�ӑ,K��w�ӑ,K������A�&�X�'~���ND�,Dhs��m�fBb-4�A9��A�by߻�iȖ%�b{�w{v��bX�'��{v��bX�'���6���@��L��,N��캷�5.f�Ԇh��m9ı,N��w��9ı,O����9ı,O��xm9ı,O{�xm9ı,N���35�\2�a�j�r�9İP�s��ND�,K�{�ND�,K���ND�,K�{�۴�Kı<��geˢ�ֲL2�3.ӑ,K�����ӑ,K����@@��xm<�bX�'�~��v��bX�'��{v�4��h@�p(L�8ÒH�a�@�J����5uR�5��WJ�F�����s��
;8fy杋���9���X��m�b�l/��[�6�<����;=s���B��';ua��Q�Mt��(E�smH�;.�M��2mJ���M� �z6�������M)7Vz�mY���[d��v���p��޴��뭹����dAa��ѷn9��n��d�4�m�,^�f�k����ƾ�-�1������踻M=��s9�ݗ���m������E�-�2��m���ˣY�=O�X�%�����iȖ%�b{�w{v��bX�'��{v?�D"�B+! Ț�bX����ND�,K�w���rɆK�ɭfj\�iȖ%�b{�w{v��bX�'��{v��bX�'���6��bX�'���6����"������w��������E�4��v��bX�'~�߮ӑ,K�����ӑ,K���w�ӑ,K������9ı,K�~���Y&h�i3���ND�,�3� B`��H�?w���iȖ%�bw����"X�%�����r%�`��N��߭��A�F�?�6��d&"�N��r%�bX�����r%�bX0RDO�����<�bX�'~�߮ӑ,Dh#C��]4��h{O|�ylILIwa��NM��[mb��pra.��s��	]��鸷rj0�8�	�x���~���bX����ݧ"X�%����ݧ"X�%������+ �5ı>���6��bX�'�����֡p˩��fe˴�Kı>�;۴�>�"�EX�,D�� ʃ���6�&�X�����Kı=����Kı=���WCh#A��>*&�M�d()%�r%�bX�{���r%�bX�����r%��!� dL���n�]�"X�%�����v��bX�'����u.d�X�̺5��iȖ%�b{߻�iȖ%�b{�w{v��bX�'��{v��bX��.�w�߼6��bX�'���[�DL�'!nFT��a��h#Cw�_-�"X�%����ݧ"X�%�����"X�%��~��"X�%����?Z�J�����w%B��Ғe���5�gI؋���z5a����ݻ��m��Ⱥ��2]e˴�%�bX��?~�ND�,K�{�ND�,K���ND�,K�{�۴�Kı/}�j��d��-��.f��9ı,O��xm9,K���w�ӑ,K������9�F�4;g�+���4��sm�̄�5uu�.��"X�%��~��"X�%�����r%���|��E�����*�V�ʩ@��

�6	�)��Y5Ȟ}��]�"X�%�����᠍h#Cw���2�e4DaI��Kı=����ND�,K�s��ND�,K�{�ND�,K���F�F�4>���dHbf	BH��r%�bX�{���r%�bX��"B*w�߼6�D�,K�~��Kı=����ND�,K���u���6�]�ӑ�ڑ�HKc,[��7l�C�g��m˷m]cv���bB�V8������%�b}�{�iȖ%�b{�{�iȖ%�byܿw[�	|���%�n���_��$)!k��z��W�΍f��r%�bX�����r%�bX�w/��ӑ,K����nӑ,K��w�ӑ0��MD�=�j��"d!9r4�Ch#A�/�=�"X�%���ݧ"X�%��~��"X�%����"X�%�~�I���s33-̺˙��"X�(�� dN����iȖ%�bw���"X�%����"X�\@�U"�S
����m9ı,B�~-%��"H��t0�F�4N��xm9ı,?� �Ud$N����i�Kı>����[ND�,K�s�ݧ"X�%��}�k\�KԦ݌	F5�^�4��\���u���=�Ni]�[ܬ�n�׮;�w"X�%����"X�%��r��m9ı,O}ϻv��bX�'}��6�4��h{z�M/�JDSDF#�Zr%�bX�w/��ӑ?D2$ Q5������Kı?}��6��bX�'���6��bX�'~����h�l@�jH�wCh#A��WG"X�%��~��"X�@�����߿p�r%�bX������r%�Mhv���6blA!AG��A
 �D��xm9ı,O~���ӑ,K��~�bX��SQM�}9����$-vv�Q7b*ູѬ�ND�,K���ND�,K�D#������Ȗ%�bw����Kı;����Kı=_2H���GaB}��dԙ�%�(w��H��M#��#,�(=А<T4��$HG�q�98�F�,���)�0"� ���H�L��	n�:�:��%`]0#	@���"��p�:�6��B'�Lk��+����)#�H��eg�������O� y
���S~�i��zu��pHm� 	,$��6Fٶqǜ�̦�*��ltB  �C �ɵVm6i��d�I��.�6�   m�  �   �@       �   ��    6�	   i5�kx�[vQ.+lP�5�"�*:F�d��D=UTy��ە;[c]�֬q�\Ւ��-�{�)2m�ڇzu�-��e���LMX��
E&�&zm�iV�t��nmɻFsg8�n�gƽ![h�ͥ�3\��s�+��nz��������],�n[`t`�+���1�'p6��-�	I�d�eِ,b	����r�d���w�T�ca�ͺN9/O=�h�r/�z�u4h�ę'd�+6�%�׋@�=]�����5v��5���`������]�\9��6�g�	���<�7���ӗ��%��x�K�q�Z�Ę�ݳ�`a����<p�cz}��<�l��ء���s��9�0e�5�JK�����.u"�ӻCθ����d���Q�=�'����Xw�5F�[��6%x�uӰ�ۢ��Ղj�ś�[q t�h��)<(�5e��y�[�}��xGm!��v^�Z,��$qm�Y"�j����0v�Y�Ö�ƚ���%��gcӳ�u�Fv�MU8Ұ+�=���N/(���J't)n��TY�	�����S"�;ol˺�E�q�rg��綝�<;l7d.����t�-��,�;r^�]��esof���UFN�Ci��y�we1m�4�����j�E͞ۃr�����󖱋����nh-��#���kd�98��b95�wdm�Q�Tv�jv_#L�M��� u�CmP��[uR����\�TqT[���e%�)t��e�x�\����&��m��pa����V�Qv:�s+ѧ��<0Y�!�z]���N(M�J���:ۛ���pǳKZ'6�m$-�=������@�"|���Qt��ApG�L�.>*��� �x(: 7�
�U��F���rFM�#��I\e�V�q�j��P���a_L�Ɗ��z˒g�B��,�t���n��[p�::+\��=��W�ٞ�����p��v΋d�Wf�mqp����{G�m�{�w5e񫥞pi�s�ю
f��u�\Vl��$�+ŻN��s��"��ݮwg�+c^��*P��u�y��뗍�I�0��s�py��b�j�4��m��^yc��mvz�ݤ.��x��C�{��l�{nNk%��hi��bE��Κqa��%�bX�����ӑ,K�����iȖ%�bw߻�b�Ȗ%�b=�}��a��h#Aq�~�4�MI$K2�.f���bX�'��ݻND�,K���ND�,K���ND�,K�����r'�B(��j%�}٫o�d��-��.fe�r%�bX����ND�,K���ND�,K���u��Kı>�>��r%�bX�k��35�̓.[��!u�m9ĳ��Ow��ӑ,K���^��ӑ,K�����iȖ%�bw߻�iȖ%��oZ)��iH�h����4���~�bX�'��ݻND�,K���ND�,K���ND�,��?����Γ��}���V�6	��=z�n@���G-^�73�m�����_L��#b3rE#�h#A���Rı,N��xm9ı,O;�xm9ı,O;���ӑ,K�������l��&B��+���4�����t2}0$!���"��Td@�P��D�(Z� ��"2�B�� �#	�+!*�D��!t��F*��&�j%���6��bX�'�e�u��Kı>�>��p�F�4��3�*B�c��C"X�%��~��"X�%��r���r%�%�by�}۴�Kı;���t0�F�4���_(����1�ʐ�r%�bX�w;��iȖ%�by�}۴�Kı;߻�iȖ%�by���t0�F�4���?}n6��%"sZ�m9ı,O>ϻv��bX������Kı<����r%�bX�}�������Q96�M�"l��Elf.{W �2e��y旎��B�z�:ղC�&D�E2)"�?w�ۚ��s@��|� �O����:�癩9	�&Ӏ����}��g����변q���m��>��M+R!4dx���[c�@��{���S�|7"I�F+1_��"�4 �(H�B�� /���<���>��ٹ'�{�f�e�"b8�r8�P�ӾVI߾����Ł���+��n��K��.j�$#�@��s@���h���>���>���������+�W��kpm����|��}mnw)���p�✺qYp]RU��7�Xn���ֹ�UV"w����:����Lj4����ۺs�}��p:np�^,�$�z=�r���6���YJ�(I���������hw]��Z+������W6�n�p:�"'{}��o���|����\�d�/wIrM�0�H��n���ՠ{�)�Uz�$������bn�EB`(6�bHJT<6$��Y��p���h���j�nՑ���2ilb���#�$�����{�)�Uz��[��^��0�"�nIuu�s�l�yBQ��J.���߫ }���uנ{�L�i�&�H!)���z����@��S@�3�Y*�pZ��M�`v(�
!V�{� ���?��=��*�^�U�U�25$l�f��uנ{�)�Uz��_�nI���,bEB,��MD$*E����r~3pұ���jp䫥�6i"��ێ  yu����tl�ӬK��F�7-��ܕ�<�Q����N�i��n3IuL=����z���W����1h�qmP��g��͇[
n�x��v]q�C�MmoW`�mvm���Ǔ��ӣr׫@�F6k�o[$�Ų�W�+ƒS,�ٍ�ֻi�܇:��.N	��z���n��fJa&��sF�f����	�@�� �1 ��Q E��Q��Q@���A)"DRB1D� �y����Mj���)J�/Ut�l�[����<qs�Ɔ�c��;GW=n��٥\mH�����/���hwW�}�tP�>���vI�����d�!
k2nI��ߵ��'�TH �A�"B��5�ذ�O�X9��g��s&Ej@�H��n��jק����0��w��sX)-E�R!��'DO�Q$D�R@S^ww��Ϸ� s���DO7��`}��]Qf�"ܑH��l�d��@U
5BD%��}\_�� �ԷX�fu4S*���%T���ٮNV|���v<�Ѷ���"&D��B4�$�A	HhwW�}�w4��Z�Қ��edq2f�s5�'<���P1P��DB���Q4?�}��5��`w[�*�j��&F�䍑��>�Z�sm�v!$�����O{��5�ذMciƔ��j)��t��Wuz޷s@�����Pj'H�ȦM�ـ9��:�Ds{ߗ�s�/��s�l�?B[�9GQW$�U�]!\��jh��î��u�����w���8W�fxy4gE��S7L�&ԁ���������W�{�)��O�{�d�}�E4��)MRAd>u:�;	(�BQT7��z_}X�ws@�e�62aEܑ8�{�7$��~ٹ�}+� ��(����b��D#�w �O{X8m�]MQsUavI3v`z(����o{� ����Q;�:`����b-Uқ�X�o䒎v���u�L���R��"DX���1	"rG%t�<X�Ã���'5u������?|�݇6I��dq�
9���_�wt��}n��������JD�5�@��f~�J��U~�,}��|�\z���p$�,�b�C@�n��v�:�$�y�}��w� �u���s&Ej@�$��e4������ܞ#Ad!��@�m +;ϼ,����|ґ���6ε�`���o:|_{� ��fߛ��?H�J`M�FK�,pv���vcu��mu��ls�sn�φ����s��ձWwwu�n� m�X��<�(�C��G�ZY���a����4m���D/(IEQ����7��]`�l�7Y̬��&Lq�&h[)�}]���)�[n�U�U�28�I	��0;���
"���]`�o� �y���h�Ӎ)���=wm�䒏BK����~�������������5SD��MH�O^�Η\ٚH�m�Vʵ]UP�$mx�CpA�m��j�]=�T3�:����z�!Y�e�*(]C˜(i�u���a��)� s�V�V�*�k�Fp� �<=]zv7���Y��qn��n݋��L|I,� �d^���=�:v��v�M�Q-������7-��MΠ���Y68�wM�&�N{J��.����������[J��[�!Fb�l��Ո@��k�q��m��q�g]���f���!��D�E1G!�[w4���>�����>^�H�2(�R)&h[l��
^�P�$$�E��W��X���`۹�}lBi:ґ��#�4�7u�n��)���ŀs�����ۍ�`1�	NI$vO� �hP �@*o=��=�{�;f���m24�F�8$I�m��������~�G�{�ՠ}掰A,q7�h{<7Dk�����v���l����/��]����J?
^Y�}E�av�Z��������>t���Ss�">��{�X'�*{V�GRB���'9�Gn� *���& 9�np���9�l�%�P�ۻ�v������倡�X�~�~~?���-�s@�����vǠ|���8M��.sYw'�� �������������M�`�78���L�&������{�S@��c�=�j�-�s@�ũ��F�FГG�jMfM�k�m-'&��9�a���mV���������oUG��ideH�h�Ďw���;$��ՠ[n��YM��5dȞ)�$���h۹�{�S@��%26;].��.�¬�.�p��ŀs�ه">x���JɪD�(HIP�
D!�y��$�WO��mN�a�Lj����٬�%��3T�3���s�#�c��MRP���omcp�Mhʋă�a�s %��y �X0XB�"@�br�SI���!H;1����4$/�t�7��C",�lBPӉu�1��¤D
_85��ň@ގcIfq@ےnr�%���Ӎtf�GJ4�f���!*B�I#�F$H�H�}|�F��	�L�KIB�2� (Ѩl���bX�@�x6-�S�_���.��1�)�T�*���]�: 
�Q��:�P6�QD +�
 h�}��;$�_r�N�9���$�	�5$�޲���u�s���uD(��{ߖ��J���+V���r����;V�m���Ӎ��~_0�Ԅ�]@�m�����Ht'��{�n4o���wi/nCt�ZT.�cf��%�8��I#����h۹�{��~�K�B��Dr�}^�����*�j�UrJ��sus�6�,�(Jd��q`�w�Z��Z���s&Ejd�RL�=��`:n�B��B��$���zp߿~�d�{�)�ѕ i�cH,����`�78m����IEB�*Q*�f.�74�,j4�"h��I��Ss�v!z P�(����{�\�~�d��ϝ�N�-��҈��(�h=1�l٤���9؆ ݏ-�&d��&���G���o��8$I�o]�޷s@����=�j�;��VF@�c�I3rO<�>�蟖) 	� B%Q��W� n���׋ �[*]\��b9�Cd��ϝ�}�ܬ�
�T��_ۚw���8-�n$�G�)���+�U?��b�Hw�~�8���� �� �ӧXܦ�i�S���G�{��Y'���n����k �)��. I(��I*/����l�3j˺����U�s�ۉ6�9���eٸ�%g��	�;^z��� [��^.�:�����
�Y�g͕ۖ1O9�����	���ָg��aŅi���s�\���+g�1˳̎�r/0�ru�+r��(/&�sؤ�Wc���:d��n������b��n6+c<���.��a����B�-�D��QFZ*�U UxN*��������(��/h�8�\��n\����%:Zd�\.��k�/�"�A4*���e��DڂR�$����>t���Ss�����ےjW��#�G�8hW]{�#�������7$�ϳ���HDH5�������m��� '$�=���-޻��e4�����H�xG��2]���ŀs�ـ|�Ӭ(���$��!*o=��:�����`jI��e4����v�޻�\�7V6܉)�Ĝ��0%n��<$>��l�����[��w��ױ#�cn�c�\r$�tVI��r�N�u��K�K��B�����߮��&Vf��h�3.�y�~��:�$��Pw��X7�� �����+e�uUtM]��m\�\����>�a�D(���	;����~���VI���GEjd�RL�>���>��-�}V��n��X�ұ�Ɠ�G�}�,Z�K�B��B]���:���,�;f s�?��Γ��{k����ڰM&���Y� V�z]�l���=��n�\��餕��svR$VI���N�u�$�q�X���~�@�K?����D�h���BI~"Q��� ��e�9Z� �g2�8�p0��RL�>���>��eܡ��+BDd�
J��R5
fQ������X��R��Aq��29�����}��'u���=��hz�h�'�G�	ݘ9Z� �o�� ������w~��~􆗠�&�t���[qM�%�68�����=�����B�����w{���Ҹ��52(����ۚ޲�޷a�{Ϫ�>V�#�dȢmL��I��v��7�`�k�u�Y�IDɳߒM�щƓ�G���߶��������^�z����]�Wf�BJ"wm�p��X�v�`w�a<�&�� V�t�J�KE��4E��XGWZB@����X�a�V�z�
�� T߾�6Iώόi�c��fK��u�X�B��:|7��0y�Zy��ģj4��cmțnpv�1s��/2<u�[�gr��x0�F'�WV���E����X�v��7�`�k�(��~��<�~�D�pqdrI���3�L���8o���M�}2Gs2�i��M�I���N���Ig�r�O����9站���r$Z�sv`y%����� �W�88�Y�n�@�[d�9�F����ɚ�ڴq�� ��f���j�$L��۽�n���~l�d�iwb��=_l 6�'M�m��A��lx�#�����#�Gn,�y4В��'%���\�q�
�3����77c�v�>۸s��g	���{A	՘�RΈW;)��9��-ٚ崝����u����,k��9\��1�p�fwg�Uu"$�<v�<��1�SNy/7 v���m�n2�`4:��|i�:݄U��k��f�@��_1�%����tV�Jbv�������E�zۆ�v**������ ��p�<B�)�����@��M�n�U���,j6�Lx���i�4zS@�[��Uz��n���:R4���Us5Sv`��`^���B��#��}������qѴ:.�TՂ-U�wk�DOk���k�p0�ـs[ŀ|���c�C#�m��u��Q����8ｋ r�������I׮�z���Ďt�SY+�;A�����u��7:ݢF�m$)��,i�17@��4w]����u��uVD�E9-J�Cd�n�������@d�K!/Dx+O�� ���0{l�>�k�IH�Q�������ˆ�ץ4w]���I��IƓ�(wX�D~V�����{���su��6_W�w���ۄC��cNa�u�M�빠r�^�����Q�\�S$U1�%L��d��rv5s�%�1F; �T��dL�l=le������J�m�|o�۬�v�З�_�������;?�?�����8L�RL�9[^��YLe�X8�,���9=a]�Su6+����� ����6[u��9ԵG�1�FMb�4�+R���CB
4 �J JT�0�T�҈�%иA�A�����ۚ�~�~z�uS�X�Dbr+k�=�w4Vנ{�S@�u�bn"����8��wX�O�����߿V������۬�(���r���IV6�����q���k�v������@z�e^�R���҉�+1T�H��)����?~�����9[^���s@��M;q��
q��)��3�"�߿=��� �m�w���"������n����*�j���=?�~��^,e�Xz�hqґ��'��#jG����۬x�$�(��D/%>��� s��=E�sWs(�.n���ڴ���9[^���s@3�܈��;��`�CR�űn�j<peZ���oF.7pj����f�-���%�k"��b����9[^���s@��Z� �L�Ba��r$����
�4P�U�ذ����9�l�7iӢ��S�J)�'��[��uv�?陟�w~���߿=�mqI#�D����s4<�䠂]�{Ӏ7��l�� ���9z�iؓQ$���N-޲��n�q�X�np
V�&eB�RTaH�� �ޡ�Is�]|��'.�ƛa!M�,.�]M����I/�u<G�$!d'�f�1%ȩeai*����Ć�GL�hQ� �M3@ca)
K�n���)p!��-��%4�a$w�ѣZYMV��lD�i�$�$	MD�֐(��� H\��f���� ^Cd�{A �)�P��b���2<( a�'�������Āf�h�mN���\�I�v$ m�m�T��Rvͤ�E iƶ�&�<��m��"W��6�  �5�  m��  �        �          H UURJ��]jOeXJ����U�Z�]�qAo,�m)v@,p�G;u�(\c����s�m ՛@佱�On��ֺUݦ;Xe݌ܝd��g�Ÿ+��Jj^m8	ٳ� �g[��X踴 �)'>:�W�qlu����&Y7.�4:�ݪ6N�׎A������X�n�Vx�v㛳�o2�Ѱ�<�;Oi-6�g4�q�Ӱ�ݱ3[T��Nv�v;U*�Н�:Mٸ�bܝt�JH�<Qӥb�n��T�\�+\f���`X�kj�:����,�뫠�*����\;HM<�������:mq�%fj��nzm!��q[uX�p�۰�R�^�Lu'm�vq�A�.xpm�rAF,�$^���������svE3�
�KX!z�ݞ#mF�v�n�F%��I����tRn�uǚ�YԾ�q�-���-і�v�[(�9�x.�n��'nK��+�h�q��= �85m���8S����M�;;�l��|c�c+U��6lI�-��B�zc<��\�����EX�v8-Td�ͧ�5�^9�P-!8�\UP �����r�	� zb �!����:ٓGmƞ�:�IG-���.�X�WZ����aL���vv�1h�ۄ�'���<���w^70�-¹�D#&�j�[���pi���Μ�W8$9�CpUsɜ��D�X�ϋ�Q�n��ڸ�+X��\c��f�oR���wk��ˣ]����ԓ��&
�.��.����쭵U^1H,Q,�6�5ur([E�B�&n�@�L3�j�U���tE[Bh�v��d��֮زdv",��h��a��X9�v��v�[��KɆ4��xє����vէh;b�H���{�w�|���|x#� 6�UOWτNw�����~�V�p��Ռsm��H��ݶ�N uU^y�AZ�����G<t�VF`��]��@�ӹ�#<��]�HE��/1g�m^8�$�n� u�<뷖�p�������;'Z�Mq�sV^���CR�s�azra:3�Ѻ��!�틆�ÜV�7Xgg�ф֞��U�6��8:��tv�s�{ I�.�n}P��vݮ�m���nW������߾�{��}�ԋԦ��d���4&6v�F��\k�7g�ȵ;��*�$�J��9�8|]k�=�w4���?�¨י=ߧ�d���?�b&#,FԎ<�o����v�e�Y�""�r�Y���8��BFԙ�_��Z��{�$�"�������X��)�����9��@������z�n���Z�r����<�NC@�z�޷s@�����Z֥sI��ml����Qή\�$�@v�mv��hܗn^�k��������߫���t,@]�w5u�<��X��8�k���~����6�G�"mDLN9�^�ފD�@"��`��AE�*�a$*�b���@� ��m��n��x�ߒ*��� ��dMē�j
8h�����z�]�ץ4���[�M�(Ɯ4^���w4^��/�S@�)L��c��G�^빠~������ ����6x�`r�n�,R��"��h{*LU\S����ݹz�u��m���k�a��FG�K		��ץ4�)�r��@��s@�Z���G�rʛ�0�l��P��;/ެ��`�)���qc����r_>�[�}�l܃Ȍ`$��(�/đ�"k{w� ���`iR���I8bR3#q�?
�)}��$��}0�l��IDyDWm�Հl��S뫯�Dڈ��s4^��/���޷s@��M�����H�h�MH�p�!��r�a-7/`��nڮeotR-��$��PQ�@��M�n�}ҟ�;�O��}����n�M�Te��oyB����w� ޻�>m� �)L�y1���/�S@�z��DBJg�� ��ŀ9ݡ�v\�D�"�'�f.�/�~�?zݛ�@�T@�V���ܓ�嶺�S7d]]�5w8��0'����;�~4W�h�ԁ���7��nqvμ�I9�w�:���6g��^܆��u�`탊b����>��ۚ�Jh�������g�@������!��'3@��M��Z�Jh�w4�VՎ?�Dڈ����=_U�_tf��{���;��`y3�3L�������f�pͶ`��`�l��	DB���Z�?ͥ��4�71���4�x�Ͷ`t���l�*��L(Z�Iia*���B�[�$d#!F�R���h��`G_s�\搂]A�i�\ �v֦��x�U��V������~��^{26���v\f!�n�b�$6�m�d4sy-=����<Tt�\c�:�n�����ҏ�bsp4��<�M�ph��'AVqO6.�g\6:ۅ�٢�����v�5�YvU�ݔ�k=GccL&]瞻G;[<ظ�9q�Mv��ut�7Vv�sў����&�gD���������ve�6��B�1uٶjH#7X�b�pe.��ǎ�L��uk?����Aћg��J�Luߌ����m��x�
��Y2B@��&�p�=]�@��f��,����)��ޅv�L\ݑuvT�\�]��7[Ň�g�w� ޿ߖ�{=UŒa���ru��ץ4Wj�;�)�w5k�m]�3wE�լ����~�zx_o��n��[z�o$m	4`����\B��mN<\��#ն�=�����p.f��
���"mDLnHh�ՠw�S@�s@����W�䓣Qē�(4��;�s�A�>0S��`�]JhS{���1e�!�� ������Ep�`meGD��MbJ��;�X��L�����������Ĝ��4�[�����M?٘�~�-�����A���<���}zS@�v��Қu��]̬�! B9p�=]�@�=y���q`=�`��U9UUTɺs����.ő;���s�Rwgw)9��`S{.�v���z+zk"��o���~m����Қ��h���\X�bx�6܆��n���M��h��;����4�I���}z3 �v�)�$	 P$�H��)"�bAV ���M�Aj��%E3/��>��{��lY'�mtqё3!��!�U
[���^��w[��_t��|>I:5$I6Hɚ�Jh��h^��=��,��/j?}E��(����A¤3��4ݛF�M��Қ���P�]7a�a���<I�R`Ӈ�[�����M��]�I(�A�>���USE�V��IUk ��5z�}��>���V/y�ɒc#ȣp�=��s@�>�@�[��}zS@�Z:�/�?��suk �V��7���>{l�Q�q$���^J���B��UX)�ArE�w���>�)�z���;Ϫݷ�����/A؃5�����n!��r�96ygy��O]m���#���ٙ
ؒA��h^��=z�h��h�lY'�mtq�P�!��!�O�z��I���߿nh^��/��'F��'�s$�����n���M׮��s�u�4�'1I�n-�n���M׮��z_�@�g�m�D8$Ɔ�h^��=z�h��h�w4�2��Ƥ#�RE�L�Kf�K$����mm�$�`���ӄ��N�{k���wV��1j�1�F�'`�q��AOPtnX�jx�7k�`�`�ua�3�j6A������݄�dy���'��n%��pTc<��v-���Y����l��bɭ���qw=�kGn^y�dwL%���V�űl�����1��s)���L��RQ����slV����wK����$W�L��'ډ��2/���y����<����@�<$�u�Ԑycn/߻���}V�޷s@���@�Z���?�����y�Y�u�����q�Y�)��#{=S�'�#nH���s@���@�빠[Қy�X5#j@$�����X�X{l���� 5��������ӑ��w4z�h�w4
�W�}ܣ.����L7���Ekt�E۶�7+�UG�u��N��V3 ��q	���3@���޷s@��z�]���P�pi�Nb�"�f�oTJ���I ��� ����B� ���E�p�$����ǯ ޼X�X��ɒB#�MǠz���-빠w�Ł��u��Ozڵ(��������Xz�`I�{�����=x�����`�qø�KLGj�=�׊ݞ�c�k������a�f;k2kv�۳N9���i����n�u�4^��^��y�X5#jC	&6'3@:���]X�x��x���L��ڙ��T\�E�h���z�� ׯ�� !%���AY�WF����p���(�h�4���/
����
���2�Lfk$�$�iW�+�
�
$(B��
���)	��4��TB4�(h���<�t���|��,G�!ÄY燏�5�ȾH�	��"F
id���B��B)��S���$BF� �"��]�a �d�!$ q����}R��H�5�,f�@�]$T��M�L+����#XeR�k+��k[81 5�i<TM �B&*i�!`�����i ������?
m�h"�C�E���(�p�C�IE���1`z� |+�N�G��i9&hz�h�w4���=z�heu��$�)2+�X�X��8�X�x��w{�������Ԫ"bk6��9�N�\�x������øNjn݁�v)�ln�-	���<���󿖁��s@��s@�[��r�edd��A�q��Z�Jhz�h�w4���>V�W1cQŐrF���׮�޷s@���ץ4 ��X��C�cnf��o���Ƕ�
������� n��-Hڐ�$��N��VI�(��>���4�]��r���M��'��\sv��mq=����m�ƍꋵ/X���WXXL�K��+\-m�_���}���s@�u��:���x|�u�#I���f���5�ŝ��G����}0�Jheu��$�)2(�h^��>�)�u빠{�*hmD8$Ƅ�hzS@����׮��빠r�eb�29�ym'��^�X�^,^�0Qp�go��`r8�@���2�:��I&�6�m� lqΉ^4�k�Y.�7F��ܱ [��g���U�Uy��:���t���ezt�����]�t�I���OM:�.�'Kx����<n3rg�鵕�E���J��$ݟ��;s-���C�R-�q�:�n��M�g]y��=Z��1��g[��k��,�A��sk��C�|�؊M�ks�HO][O���;�����s���lt5,�[c��lʼ�8E��l۬����?|���ٛ������_ξ��7��`�ـ|���9!���Y&��Lm��;�w4�)�}z�hz�o�H������ L����>��|���5�ŀo5��vV����5!19!�}z�hz�h^��/�N���lr55wk ׯ�(^�︸}��|���m��~��/R����d��s���K�ڱ��Ռn��3kI��.��=�l��H"�$﷬Y'{g$�oX�*�W��/��s@���Cj!�y&4'3B{���߈9�*CJ'�o훒|���'}�b�URD��ɧ���j��}ŀl�u��I)�����$�w���q��H������\��X��X��`=x�H#��J�D�E�ڹ��y��>����nhzS@�Ԯi6�4d�/.�wW.K�țz�pe�Q��;p�u\�"N0jDԆLlnf�ץ4�]�^�<�G�_q`�ڙ��T\���-M]ـ|��Τ�%2>��=}ŀw�q��P�M���I�iEM9nH0��� |׋�PB�B�%$�	/���:٦�m���]C����9�Z���СD�_~X뾘�XQ
_^t�7�ӳRUM�V��I5k ׶��^,^�0�x��DB�l���n9��Wv4<"F��jV̺S��m�/\�vz㦋m�rv�k�l��������)5g ��`�ـ>k��I} �女���� �cRH�s4�)��L���X뾘�X$�j�U�����Hh�)�u�M?�~��s@���h�Z��R ���!�u�f ���m��D$A��K��h{+J���Y�����/��hzS@��M�Jh�jo\��2'��SY�ۥ�vۣ[C�\%���<�ϣs��L9C�f�&�M5$m� �O}��_t��ץ4�]C����9�L�Hh�)�u�M���ץ4WJ���cB��:���}�s@�Қ�Jh֕4�L����������}�`��`�l���u�l���_8�.H�RH�pY�)�_t��ץ4�wdY�|L��zӅ�]p�I�6۶�I���7nSfN��)ivK����ں�ыa����Tl��ki�<M�y�3�qi�Yk�f�;5�<��cp[.C1"[�F�V�`\���wş�M�-�N�}^{]`�m�܇kb��nu�$��7fyLW��i	�c���m��Z8�ֻm 
��vX�n:la�����\�w{��u��I5���l�+vGs�pt��4u��o�}�"��Iv��4�;��ݚ���'vk~��}���`��`�ـ>T�AJDԀ921�hzS@�빠u�M��4ݕ�do�,�HLNHh�w4�)�_u��;�S@�>I:Ҋ&��8ܓ4^��/��h�)��E���@�~u�pi���&E$4��;�S@�빠z���{�_���8��ԉ��qųVl\78s��q·o<0odL�F���<��g�W&4���/��h�)�_u���94��7)�)�d�������C"!B�Q��}���5���7�ـrm�$BI"���=zS@�빠w���}�s@�_�u���Jc�awf ���v��^,����w����R&������e4�]�����R�֒7�6����1q�6��������ۼ�9�L밡���_ͥ$o �%1�C@��M׮�|��g�;����I֔�7��ㆁ�t�}�Ɓ�t��}қ�L��g�Q�&4�RL�9�~��o��q
����+�PV�� ����=]*hC�PI�JC@�YLx��X��w�:`;ӳSV�ʫ����j�x����/�޻�w����|�eX�r$�4A�$�*^ŋ��&'������<��&5 ����9*9�&ܒG!�z���=zS@�YM�e4�_�uŊ �9$�h�)�w���޲��]��ڂ)sSv�VZ���0�`�l��z���ŀ?v�`6L���d���J���x��X�0>Q�^"!-CZdB������ܓ�M}m�un\��In8h�w4^��;�S@�YM ����dk�D(i���$43����ѓ���3�@ʹ݆��/Lf[#rdQ��=_U�w���޲����ϐw��s@����4!�($�(��;�S@�YM׮���� ��i̙�㍉�@�YM׮�����e4
��$6�r7!�ԧz���7��8��0=�){��_��[�(x���y^�@�YLx��X��������+ �0�C.�h�!	 "�A�L#,d�A)�
 R!�	�jA� PcUeF %!
BơH�����FB2$#
	MMCAU �HƤ�@IV�T]J��,$`�"@�!$�($a���*B	HNh�۠�0���"����&aZ%eaHT�i`c"�4h�R�d�$� �M��3I4EI��]�F�HB4i&I!� IrͥH�B@ּ����3)D�9\��J�5�vm��ml�n]�5��#��f�cm�*�Jm����1���TQ�.m�  �m��  �  �      � �   ���        ��m��[b���۷��mx��YY�n�
]#*�f;$&�Sj��5�7g�[nТ�e8F�6��rC�3������@��XT�p�����-�kXm��m͵�k<V\Zr݇{q՛y�'���"�;��:1�kv��r3/8'��ڸ�챷��� l��u[l�Ǌld�Gm�5�c�o��v���l��2�T�J)Fy�0�v�������v�\]�� n��cE�oN��߃uz|��;3�i�<��\�c�4VD�$�Cal��˲��'/N�-��ѵ@u��1���,	�q�۾G_R�'<v��P�ŬCI��uԄ�����t���qېG
�(�m�a��P�ɱ�NeyC`�h�fu�-�h	��Z��Fb��R�3d���Z�#��|��K�_Nl2�۶㖰������s-r+i�0���|�}�ukRh�FΉ�vSv(
M�o0p�9�Np�[��������[��i��[�q�WN������Z�t\v��2�<^�72��A�
��z�ͻV���R���挶�3V02�����Z���8$�ki�\址t/8�8:�rmP���!8N�Q�@�%g����;	�m��v�U<�Wnq��c��ޤ������<�#���^^�id��\����
;�6���q�u��\�7PtdvK\ݵ�S��ӳ٫��� �)+u��7�9g���pb��έ�MIm��ev� �rkz��A�5�ۦ���oPm�M���a:�4�5H'1m��J:Ls=%���2�<Ks�۬�4�ś�[j�nȥ�-��,�$9�������X�]K����x�̻.j�e��.fk31C�0 ����C�?o��
m ����'�����5u�j�ZL�k-�ͦ��f�v�uR�5��WJ�C��y�ꚇ�n���K���dԆ���1�v��7�ݤ��uŤe��i��I�Bn�]�c�R3��{u��s��lQ���݉�������7\���mk��vKjls�Gf�.�6(Ixӷ;���<k�Ig�6v��F���#��q��]@շ=��\ ���fzx�%����n$�&RJ������/NF�!-�Y�[�t���\s�y�<�N������[����8�(FI�8L�)�ߺ~4��:���*�W����v�ȔǑ���4�w4
���zS@�>I:Ҋ&�r9p�:���*�W�u�M��4���[ɍ�RL�9�}�hzS@��M�]��Ҧ�N!@y&8ӓ@�Қ���Ο ��� 5��D���$WӑJ���mR��l���^O/<[�܃���3��M�D�#u��̠����m��x��]�(��뾘�zR�"A!n7#r^��}�h�ـ>m�;
ɱ07�*l	�Ww`�� �߿M�Jh�S@��s@�v���a�$iɠu�M�Jhz�h��@;��'cY�(�9!�^�M�]� ��hzSC~���w�gB��mltH�Dl6";i�����J:
3�u�[m�7J��I��Ғ)p�:����f�ץ4�)�}��:�Lo�rdQ���f��m�ݶ`�ٝI(�7�ӳR)��l)]�����]����	L��� IE� `� �!�$b1�BF��d$	�,!$R����b���;��o^���nI=��rC�Z$ә271�I�@�Қ^���f�ץ4��VD�B%N���5� �(��������`w�Y'Q�w��ă!�AJ8�	ڶ�x��wc����k۷[����m�[�<�Tl[a�IHh��@�Қ{�4�j�&�L�'&���M�]��Қ}l����v�YI$4�w4�Jh��@����|YZR4���H�rL�;�)�����fq!jR�D�$$%��E����������8}�����Lo��d��@/��ץ4�w4�Jh�J�q7�6�i�D�O5+8�9�N�!���[yv̯>�̎�N�zge��bz���c�I4�Jh��h���f�{�i̙��F���{����M ���ץ4.�VD�B%NF���Қ��4����y�}0���D��ԩ�WSw$� ���ץ4�]��Қ�P��p� �ץ4�]�y�� ���ĢB��76E�%j\e�
�bx��@h�t�kn`����t��=; ���kq>�&"��m�M�^���Ǹ���r��jz�x�s�Y�v�x���t�!����Qyls�=Zs��筺�p��\��^,/���e�G^X�ڱ�	��Bk�s��0��`5țu�	V�L�����t�v^�<���`�gh�\�ی�������*hմ�Y�+t�X-�[[e�҇%�7�sln4oV��k���r[/Z'�24�� �
0�Hp��恼�f |�ߡ(��C�w� l�35�J(��ȤrAd���7��D���Y'�Y��;�w4���[ɍ�RL�8h׬�>���;�w4�Jh���4b�%�I�7&��}V��빠o6ف�	)�u�������V�j軻����7��`��!�Ο s���}_U�yvrbDX��n�ț%��؋<ql��<l��E�u��c+ӷ���v}��Ù��H�π�g�@>�f��}V��빠{�a�qb�q)���}��f�Y* @Yg>׿]��s@�t��}�����2;����Z� �kŇ�L�w� 9�٠q��� �	�@�u��;�)�^�@���@�|�n��&���n���y������>���M �����7�6�g���;�M/�L�=;���<.W�u�x#�=�z�Ĥ$�"p��Y�}_U�w�S@�t���[��F)Y1�#�h]�`�l�7�l��w�I)�o�)4�L��I#I�@��Ɓ��M���AґB#W%��rO>�>�˨Ց s"Q������M ��4�Jh�)�{�a�qb����	�� >m�Ԣ:��6���fԡ$������,*-��{/L:�'fB�"�n��§^�(<��p�u\�ӡ#$1�dqI'�{�����4�Jh�l�����"�S	$���Қ{�4��h^���&��l��ۊI4�Jh�l�>�)�wt���WP�y1cD�p����3�;��9�}0ݶ`R�$��SvN6I��Xi��!�$�>�)�wt����M �-�?�����cn��9#\�4@��n;v�m���p��'m&�R=2��Mu#�4����Қ{�4��h^��>]F�����H�4�Jh�l�>�)�wt����uŊ1��I �-�ץ4��;�)�_c�"�d�<�"��M�ҚwJh���٠����0�)��C@��M�Қ|[4�g$�1B�݄�r�j8�M� s�����f�- m�m����n�]�]�f�5�t�GF��:őlb���c�bt\5������]H�|uv�:�nŧ;��M��cBe��<j�V�\���'[+��Z�V���ΨS���!7WH�nlA���nոE��F���ܺ܊heq$�v0�O�3�F�C�&Ş\�l���o]�u�q=Z!}�U]^�(��7��E���RF6�ݴ:T�n��]�m7	��0�³������#h����g�@/�f���M��4���[ɋ�$pq8h���=�`�l�7�l�(Q
d���q��R$�c�"��@��?wJh���٠֍52L��I#I�@��M�Қ|[4�Jh.�VD�̉FG$r{�4��h^��;�S@�o+��#R�nu�ve�$t�qץ�4u��c}�����N�'�&�]�w��qŻr�ݚ��m�����ozq�{ψ���@�c�R()2#��%�s�q�*����
�B�"P���[0��0�n��hN����I$4��;�)�ų@����w�4݃dm��q��(�/^t���x�m��m��]C��Ńɒ88�4��4�Jh��;�)�������&6,�j�f�͹هQ�p���]�#��2�7&4ъD��dP�h^��;�)�w�S@/��@;�jd��rD�����M�Қ|[4�Jh]F���Dr)!�w�R�'�{����R��T(xhy�K؆��P�2 @'.�s0ܺ� A�D�1(�������d�g��8.�au�^?FC�x) ؉˦y�	u����.�=@��bnB�.�tK�SX��k.���!Ð#	�\�HMp<�$�#�������),!
�P�Ť)Z��!�6��0!�08@�<4�h��ˬt���!b��HU��'�䳜��9�6+ H�M8�4� �X�D���D�Lb@�6УBJ�{e]R�
�DR0`@�@15���$&�؀�T�#YId�#
��@�R�jH�	�F�h�-Rṷ�"��*QO�����".��P0=E_Ec�DS�� �{����}�S@��ú��1��)!�ų@�����Қ{�4�|R(FL��29��>�)�wt����M �-����5��䍡&�,��7Q�4g��-��W������7�'Xq]�aN9L"Ja$��;�S@�t��_��Қ�ɦ�#h���{�4��h^��;�S@�+�u���y1���_��ҚwJh��;��4ъD��dP����wm��m�K��B��
��@*? /����srI��٫����rD����Қ{�4��i';g$�*���ɦ~A%"J����t佛bɞ��<\d�V{���W��G/b1��"@�DG"�z�ƀ_����$��m�Ld@��M��������٠}zS@��M�җ��C����F\�I��>4�Jh����>�d`��&
"H�w�S@�t��_f���M ���v�0Q��sm� �k���y��DG�K��ؒ�1n��4�� v֦��x�U��V]��f��b q\����{]A��t����S����p:�]j$qiz��ˇ��sGD�y��i{N�Δpt8c	�P�q�ڧ<��vv,q�Gj��`cs��.,�vm�,]Z�k����K"N�O��㇄ݎ�mݧq���RC��y5�W��u҇d8�^yHU�-˸&s���L1�ՙ}��΅�{\	͖#VJ��<�؎ݫ"tnH@0��x9�[�Ӱ�������������4�Jh��;�)�}l�\f'PI�Aɠ}zS@�t����M �:� �£Jc�6�$���m��m�zd�s��`��VD��"��H�4�Jh��h�)�w�S@�0/��9�9!��Y�_t����M��47������ph�B�ۊ��#���ix�<�N�{qt���B�|Y��Q��K.��� |�f�m� |�gb!} w��4~��0O�0�QG��f���b�� �*H�B+���M�CR�k>����r�@��M �ri��<q��7$p�/�S@/�Y�_t���t����u����Ƞ�p��Vh�)�{�)�_t�������$ȣRh^��=��;�)�ܬ�m��q���REwm9�[���gg�u
����Wbݠ�9N{\�c�6.���!sB�qē���t����M ��f���M�Q�"CSQ�����M ��f���M��M���.(�&I�9!�ܬ�>�)���3#	BBHD!��� ~��ߧƁ��M�)&9�R"9R`=�`��0��0:�B������" O��$p�=��;�)�ܬ�>�)�u�pdM��[]���h#b���Zq�F퍮ڙ�u�sx��ݫ�)0�t<���So�������lܬ�>�)�{�)�}A�:�LAV6MMY��.�!(�9�}0�$�q�����?�f5q���(Ԛ�Y��=��;�)�ܬ��G���DێH�p�=��;�)�I��߳rs��D�A��D@"H�`1T� 4�"B�UU�-v|l�����D���J9#�����Vh^��=��;���Һ�;��J*�m���v;[��{muk�O��bv�ݰ�ڵĜsL]�� ��f���M��M�Қ�"�� 
DG#jM�Қ�Қ{�4���֤D	�c�!$��Қ{�4���ץ4	��i�0�%)�8l��U.޿��?u_����M��M����,p"�i�@/�Y�}zS@��S@�l�d� ��Úr$�FRD"��Kf�Y'0pm���m��l�㬯SE�v�vݮR�o`3�b�{Zy�<+9���mt �
�5G,E^��a��uD;�1��mA:]��ʏ*��^wS��%Lu��h���Z(7m׮��p]%��J�BJ6�.�;{nWlj��cc�φ�WXzI;6�W;	�U���սG����	������r��`���b��wwv���t�.���U1�U,��6ѭ��Ӷ�۲�\���	cvYfH�c��dQ�4�g�@��U�w�S@=�Vh^�)n9"I�@��U�w�S@=�Vh^��9u�dX�S�(�NE�w�S@=�Vh^��>��hFqr<b���]ف�Jgu�o �]��>��8��4yґBc�"#��&���M�}V�w�� ��Y�{�)�q	�6��p[�DGl��Pڷl^�ͷѺ���nON�4�GLJ[dt��"�2}$�~�� �u��r�@����{�4�Șq���6�VI;��d@P������f�m��>��hPu��8�Mɠ�+4�Jhs���hz�\dj1ǂ�2(ԚIBJ{�:`t�8 �����w�xT��M��N�Қ���_��� wU�h�)�r�:�H�:�o��j��v'���.�';�盤�:�Z����ӿ�_���jM�!2U�[m��~~��r�@��M��M���\Pi'2c�@=�VhzS@��U�z��v���)��4'�{�M�9���z��U2@"�T�Q	Z�un���w�6�B�4��B&94��ZW��{���)��M;�8�'ڑh^�@=�Vh����}V�|w&�"^�1k�I�&:W���m�d�8�κ�c�9R����B;�،��#j��ު�ޔ�;Ϫ�*�^���:�#Q�<X�țRh����/;�h�����U��֋�E"m�$p�;Ϫ�*�^�{�Y�[Қ.��D��J8[�Y?R���;$�ߗo om��D("B�	�B,B1!	52��LQ�����	I%�C�� �\ P���d�^A|���p@ZwX�9w�w�y�����^��7��}��ck&�4����d��n���׎<.��'���-��j�B+2�$����4zS@�>�@��z.ꞁ֥��1���G��[�?�1I���`[�� ��3�!%!����a�$�R-��=�q^�oJhWj�>�u���A"JH��k���f�M�b��u�����q��&8�O@��4	�C�ｾI;~��'��{u�'�EW�Ȋ
��EW��EV�(*��AU��EW���
��P G�B#���� �@X* ��@R*�`�D� 
� �E*@��AX*X*� �E`�DH��@�� �D`*R
�����T*Q *U��`�E
�A�� *
�E *��H��A*U * �A�
�EH��E �D�*F�b�E
���DX*F���T��`*R
���E"�
�H
�
�H��*D *��AR�b�D
���@�H*R"� *X
���EB"�*  *A`*PX��U�@ *TH
�QX��H
�QH
�`*E��@�B�B�"��R� ��E��A@��E�
�"*V� *X
���A
�P ����@ ��ET��D *UH�,R�V� V(�B�B� ","*P��E��� O�"(*��(*������AU��
�EW��_􈠪��"��� �
��DPU�AU�AU�ي
�2�ΰ#����������?����G� Q�*���	 �{             4� 0  ǅ)M,m&�Y,���Hu��&�-���gs. @r�Z�Ls5Ђ:͎�u�tt�r: Et�td�1]4r4u� ݁�i��-�w	�h�
 ���v��#�b�FF�����F7  C9"�6WM�6QN�����Qd�]g.  �:�ٗ]f�4R��R�V�Aڒi��)��p z   P���S?�SQꞓjmC��A��@F��R��0&F�`��&��Ѡ�~=U$�T=@�h��L��5<j��UH       �A�ɓ&F�L�L$@I"i�M5=#MF�z�Q�G�=5=���|+�~?+_`TM�?}��AS�?�0�(�KS���L����?�~C'�����eR/�A��I'�0�����D5!Dq*H;��7����\״���[e|�q�v����
��(1�w$$v%�v$%݄��D@���e
!�UHɔ0�(4c"cA#&@� �3  �	1),a($$�+BF45rPH��1��D3)��F8WVF�(�"
�� '� E� �>EU�q�B�8� K�c/# �p(5v1�
�$'B�	�L$D�"�T^�KG�X�cy��f�xZZ�,�Iќ�.e�(�?��eZJC�N��{j�ΐNY�B� ��%�Ǣ�#nD�8(Dr�l�ƴg��W�j�"ȫ"�-��sjp�U�H�&([��<]O0n�@���x4/�'#Gc�B`��a�a�P��B� BP���P�SB%�Q"a�<!8e��x�uN�ąX���`�����b
&$��Y62�f�$a��Y�hR�� �\� �hCZ�Wڄ�\��-@ˠ RؘL��g2�Ug.P��$(��ZB�9��"E�Q� Ų�m!VA+s9�aC,i�Օ9dȾC��h$FH%���T]-�`���� ��,�Q*QF�1")#Wuz�������p��B2	AdXc&-��7x�Ƌ�oMܓ�ٶ�� �s@�H�x�T[�� �42�9��E���e��!���F��zm�Ad��޲(b��s<�l�����9F�v�t���4�N52&�|ͳx��)n�eCB�RGhA(A�X� �M�l@Qf27��@#l�e�;��]�ɭ��8�ك)�gA��`�kzvÆެ���ζs}ѻHaV^�٣d8   �MX�����p
l�м�;:@�  �T�c4nU���)É�vÀm`Qq��;6�4��&MJ DS��D��n�L�c[��;��[�Cp�=����;]���Jr̦�m�;=ҸmsC��&��3�F�s*��[�jUhy�[�4�&��΋nؑ{����e���Z7��l�li�ٙZ�s��Y�XpP��D&�Js!�vjs��|�Gk���y����v2+b�jR=E���MO���g�b]<���e�[�(p�.�U.�-++��Κ���9�[g�?@           6�    ���                     �                                                               C�                                                                            �z                                                                             =@                                                                            ���                                                                      ����/{���_l��d��\����D��ne��:mH)#Yd� _-b��[CN�y�m�h��m4���� ��"��MײJ�l$�Kj��n�n��kn�W��FCjؖI��mH�e�"�!�l��xi۶�&m��k���M��m�nѭ^p�$���n��-����} � m� �  h��[@�  H�\�^�I�@m��h    �m�v�h�K4�I@[A:#^����T�F�ݷ6e���$��$�E�n���KgO������kkj�L�mu���;om�m� ݻH�mm[&��mf�����?���g����nNKҋh�ۗ�Ci6�-�[E���r-�?�{�otP�G<ͫ[%ݧIG;ia�[v���趀[@��e�m��l-�m��� �&�\6݀F�e�6�#��E�N��ãk],1�N����:��8�zS�[�fk}��6�& �YF�e��Y����I,��Y�U�:@ ��$�m���1-�.��.E��	���9[H)M�Z�0��n��l��oHnܮl-h   � m���kv� .�  l �$ݶ9t����zk ����f�Ӵ��_Dov�;[$���l�m���l#E���ScM�ٶYg����L��	:Lo}��U�Ȯ�'G[{:mu��iz��ZA�j�rV���3�fwV�	x�$F����+ct4����ŗy�U�ĳ�����{�����ׯ�UU;�_g��c����(���������zQ���!J�����8}e?�Ƿ�ہ�2^~�g��:2�l���)[Ʃ�4��T�ӊ�PN���CRt ����I���`��3
2�e )�/R�E
�
�T��8�
lV�!��눊XeA�dJM����\��S��aI�drtwe�nm�q��܀@��u7��Q�EL�(]��A'8���
��c͜
eW����,��7V�X.B�J��L'u��"$�[5bi3�s��2��n����}�
��H�~�l�J���� �P�2bW�ݻ������'tQ"\	4�4������w�ǿ��lm�  �            l              ��              l              ��            �c�{�.�k���In�[y7-����'I�aZI����[m�km��nn�:M�l��)'i,�W���,��з�s4l���ۥ:YJ����E��սj/N��&ݭ��[;j6���&F�Lt�,�X��j :F��ؓ"���f��ur�n��]zT��l�4���'�@���X/u^��ĵ�W��?����$   m� m� m� m� 6�%��k\�4M��D�霸�RFdXFG*���Ꙛ�5T� P�T))m��m��%�HA�Q-4��O���h�_|54wov��������ܹ��4�U��K��L����]Гg�H �IB.k���t�_u�w}J��}�D{Ѝ���'|S�����Z��)f���j��SGv��`�ʿ/�  ��Z��5\V�fSv��=	���9ݔ>ס2�j��`��z���u����*�[y2s�������  :�6�.F�2ܔ����ױ;^�-ڻ=��'ÓGv���ҫ�Ŧe�;�"&e�����fo�3�U���    5?���H�t�R���6J���N�;ݘ
e�|/��y�Am����V��nV�m_1��N��������Ƚϣ}� �               ݹf[�y���]��rj�ʙ�D�,��t��u}��=�믠 �d]l8�dJe.��UՅ�Wk��uN���ҽ���ͽz+v�=����S-w]���;�����  	��$;�����6·w�;I�٭��='�B$@WtD�̣Zݬ�,ɼ�U�6X�9��f��vW=����~�    :HK�e��fms3��v�	��W�u�� �^�(x �}����h,7�s��o�f�ֻ�g�[~  L˦��8���-ٽ� f;�M���7����X&��[{�Bj�o'j��Ʊ<v*{�\������    ��`��D73 �^�n��R��q�e]ɞ�ܭ�>���b�%�Wv�h@���98���3���ɍ����@               m�zK�ٺ��!+-dr�&Ylr:��W--�rڈ����^K��Io���P  t	���K�i�%f�ʝ���Bh�� �����L�ʼ�g�ւ�~u�nߩV��?__>~�O}�  <t$V��5�L�fq��.�N�����w>o˱��x;�5篋L��[��3�|U�y��������  �5��8�ܹ	��*��{kAL���~��Z����g��*�^=k۾��ڑ���0�L�(f�4���PH��@�DR���
^U���bØ(!���+\@3 �n7��;�c��0ˇ���|�{/��<(M$���(G�D��=���xo�gW�}YŹC�绰�^�2l %��Y����gϗ�  &�[wK��%4g���~�"n����I�����˙�ςk���;�7�?ʿy^k���8 :{t< 1��϶��L��k��7~� �cv�I��m>�՛ys���V���N״�j�UePג�14y�gu���I��������_��w�'����$m              	%���^��n[���˼m54��_�Aq=��C
o{ZI}����  :&#[���3��ϟ��>��ס2�E^o!�����_wٕ��zo��}�?;�o�-���:��Q����  $٥��dݭ]%�W����[�G�&�{ހ1	" ;��{�DN�����5w��������Y��g;�}�~ˊW8�<��8�?~�    ��
�+9]=��/{�{���[{��;�������r[�ݓL(��@���}��_@{��� n����U>��Z^��y�kM�r~    "�`J�f��d]�y�,�r�=ӝ3�|+{�f>���U}�M1�,����X,����gs��W��  s�s��&�2�뾫�sk�\�[7�k{���G�����}�w=��/��7P��t�]���{_}�b����.�a/����              v�ѻk��vw�z�Z��6�E6����v�t�5uĽ��,р ��{e]u��R��h�
�A��!��6�ڡ�{�4� n�9�OAm��,@�[�Fb����nU�1Ʃ��l�8B�k�\���ϯ��S�ﯥ��� �d]#��c{^��X��ƞE�߹�*�x3;!�0�&� �CX�@��fN��.��̳C�v���R�#&|܆��N��ƛ8Q�{o�M��܄ʕ�#����ߚ�� f��������km,ɶw�[�~��M�k�D�=�l�K�.Z�;�����@������aP�Q�h�1o�[�SO�*���R��=�*�o��p   $�%������4��ww��c`�>�Α{��tQG93x�H�{k�M��ܙ����}i�-�>����tyG'�yň�`���ɧy��;I���4����EǍf��䓀    !���D�-od��,�����TF�"@y��&��' ����	�e�+׬���h�F�Dn��Mw�2���w!pUy��7Q?#�7�;F�������ؙ��Z�c��U�����<�0^L����PȰȱ(���n!	�^F�J+ܣXѠ��E�5E��`/� ���PB�S*X��aP/cL�$5����L賥0���h   m�                                                                        ?�z � ��K�U�:����N���F�q2(�ۊM��lm�k5����Ҷ[e��O$t��xݍ�9�^�zx]��m�����uv�z����XV�k:b�e�4���u�H��V�nAV�IcH�ݗ[ڇ �Фh�Qc9�W:�#�hN8V1��%\n����#��/߼��}��@Ã`;�Tv��=����E��'��|�d���  ���           �$���݋��j�,�4u��Eh4(G[��
����ޒ}w��p  *����O>z���K�����|CI�l���-��N� �i�Lv����:c��n ��)�ל���,�EI�Q��9F��]q�\�L*��8����E��3  &�[��<�u� �@���դ��|��4<G���dQ0y��۩� �wZ���r�x�� #��ڱ�� cH�(� ��g�N��qDo�2c��^���{�=��  <t$V��� .��r��q���Dn� J"i/��h� A�I�u#������+'w<�!�f��.U1��
P� E��swX�T�{k�*����7$nw�oyT�����r�Oƞ���՟Mu�s����    )]	]-�-�[��������5>���MP�Y���8�܅�Oz��ۍ(ɏ��ܸ����?�r�xDJ���>yF�����QX����3~ch�����&�Df�t�̀ �m�\�Fܻ����{��8� #uFz��ӑ�qP"��3�_��hq��g�G�>nChYϾ�O�!�QG����v��T;�'`@ďG1�!5�$�Am      ?�=       �tT�K�W6�t[6Mom��d�%��Mі�ґ�wo<�g�� �%�()�r�Jd����{�X;�f�~�-ʡ� DT�TI�m)����@V�5�T��������@��D����ϳ�L�1�{.������[]�;?     ��e"gDD9�t�6�q1�` B[������;��� *x��E*zZV�=z߄��Τ<��6N��~B�;,��b��㈒��È������my�4����zk�����ɰ    �UZ;d%,K2.�\����o��+%���+�%BwTy ������Ӛ#�6c� 3� �pD\��l�����h|� }#��T~���>K��/[�ڋ>�@��8�'G���~o� �$�6k�wy�:�Sj�QgA#����{���r�q���}�	���
�^���nU&J�^�<\������`/|�s�����=&�Ƹ�ª(��&��>}��w}}^���u�  Q���R�L�S)�1�]�7~�$n����̳C�x@ ��c�F���Yٟ7A�y
�E�f��ܐS,P��;PF(��z��[n4��P��uCB��O����r ��         ���  ��H��׮(�n�۝��m�&r�V�}���l�Q G��s��  �#n!!��y���}�/�~��(�K�\�b� w�<�#y	�5���Ѧ{V�� n���YM9t�a����~���hl ?w*��j-i���    ���i�N���@S���'��!x��a����r�s����b�M%"CS���"!o�:2�qc�@��܆�����U�T@<�y,]!�p�I}��C�=�<=3�<G�QGzկL���̀8�������{����wϺ8A�a?_2�st�u�=�̳CHh����T��k�T������c*�Pʷ%J�$B"� B �D�H��0�� F'���ޫ�K��ъ� �=BZY����'E)���q6���b���U��6��"r��Q�xr���Uwkޚ�g��ן�/ܳ�    � tl3{&�����,��*�����%�T+�Hf���r��[� n�V���a_xrh���B��",E�@��j��L'1�(���ڏ����}� A+]�dl�k��}�0yU��6��_&oiG�2��܉u���[m�	 f!v�n�y�.��m�Cڈ����v���ԛ}��             �nY���4�J�s#Z�M��rC�v�l�5V�M��*�^� �K&��55�|��+q@U��47WD����p˽6�4�1gu}��G��Z�lt ��=*0�!�~nCj(�sg�79�w�������  [1�\��U@�]��G��C=i�7wo&5��pRD n�h���xC-\+oG��@v��G���8�Ҟ-IQ�Z"x��EG }��Ѧ{�w��_4��,�<     ���NJf[��L�aAhfh 1����>e�E$���� Uy��7P�AX��@� =�2�z#��11������ێ#@�@n������  :+Zq�������&��[�9���^�r�i�$kqF<�M�/З 7J��pi�#�q@�D�A����V�����5��}�l�mzMc_;	�    )]	]{Kf�nժ%��5��������]�a@�_G�}��ێ�J$��d���7*�����'�qW�@��:Y��O��y[^q�J��>����~�>6ٶ�             d���5�9WE�n�^:mn��ݓY���/f[mL��G�q7��  S:ۤ���%�}�����w��35�{8ژ��P�] ����Y��
�xr�#�TېڋGr�4�� �����~2��l��� �أ�O���  2뗨�58��iHٹ�V_��C�a��ޢ�S,��U:�]W������C��|F�9���ͅ�?<�w�n��S�bh�}��zffd �������ǻ�4����W�Qd\ϛ��H�b�>�q�qA�W�t7T{�+`��gDE��� ;Zw�>��<D��j&�G��@�ӻ��Mc���9     ݢuUh퐔t�,ȎMg���_<�6hw(�4�v�~���4�1p��3�|�4>z �@�\~�2�F$�5��D�����@v��� f֝�;�w}��?��  yI)����.����Y@�B���ی>h��,N`qy�nU 9\#��Q�&��r��&׈�8@<�qM��>��7��y��ާeY��-�h�DD�;���;_4�7,Q���L�\���m�߾]}�[@                                                                              *���M�9M�m�����J�.:�jK�"N���km�6��m6Ӟk1��m��;]��u��z�$�^��WȽ��n���ڙ�2i&�l��泵�%�ݹ�%n�[�i��c�W*uK�)��L��[k�M��:Nm��#IgW�-�m����TVXKh���W5���m\�'@ky�Z9�y�{�|s�<�]�mm              	8I�F�]-ͱgL��n���5�G4�hűu;���  r�oh�����zm�ϐQG����W�̳Rx����Q������b��i�=�&�!�d}�`�]��>��4�7P��<��aP�]�?�ϟ/�  s+np��y��&ʱ�(w(�8 �isR��[�Q���AHH�<��x�A��P�Ey�)�ZN�# n��W�St�u���o��Y�<c�Tj��4� gy�w�g�|  <]5�l\]���Ȓ	"w���Ln�I�9�$�n�A$O<�J�yMA$��A$<�"\A<���I�����T��c�.��aPI�*	 �����}z��}_K.�;���.	 ��ؒ	"o^o�U�SPI=1,��j	"kt��O<�D$$NĨ$�^.�v^.�� �g9I�%�'���,I�;�K�H'(�$D�{��\�1� �*�a�&��w�A<��B��%D�$�yEb�D��.	 �~��]�c"H�Z�ȕ�MQBH$��R\@�&�r���$����~\���A<���I[�� �yv$�H��PI�s��6]A����\E�w�X�	"v%A$
�L�:]�l�$D��	W/)�$�w�bH$���t$�v�D�J��R\N�w�w�<��_o�  &L�e�36%�PI�����D"����$D�i.	 ��ؒ)"x����WYMA$�R2	"c4� �*	�݉ �'"TA/^v^.�� �'{CpI��ĐI�*	 ����I���˩��ODG��ĐI�*	 �QBH$��R\A&�k����D�I�*	"��w��A$L���	�]��Q�&��������jIo��	               �sn�tvg[rHj�f�yW/ޮ�'jil��;58�����K�zI%��_��@   6��ei]}��ZM�/�k]z�IvR\A=z�b	S
�ȕ�Nc^��wYA$N���� �q�1bH$����NU �'�^k�U��j	 ��ؒ	"n%@ �B� �t=��g�%J�'bv%A$Y�	 �'{IpI�!�ŉ �D��s�U�^SPI�I����`�	�ݩ'b�*/I�i�4��� �a�Al�cXļ]e�Z�H�yIpI�nĐI���$�n�I�;�W��S)�$�w�kykQ"�m*b!Q9�
�v�A$Nf���J�M��	wu�� �'"TA5E	 2'9IpI��ĐI9�ۗ2��H'h�$D��.	 ��ؒ!$����M�>]� �'9IpI�����D�.	 ������<��y��߫�@ *�e�bc��9%Y/!��$�y�ؒ	"b%A$�(I�7�K�ȕ߭�8%\�����|��=$�����I��.	 rj�I�=k��U]e�7�N�BH$��R\'���XlT�4H1�� @�oh<j	�݉ �'�*	 ���^*�� �D��K�H&�v$�J��K�HH<���I��y.�SPI�˱$BD�J�H<��(I�9�K�H'3/�w�0 M�ۥ���z�{�nՑ$D�J�H&��$D�).	 ��ؒ	"g=��r�SPI��>�S�$��R\A<��I�<�PI�9�w��2$�H��%�$[�E$ND�$�n�A$O^w]%\�����w��$j-D�J�H'h�$C�a�tׇ<=�;t��L���.���j	"r%B@$4P�	"s���M�����_;��}��� :d����J�
�����	�$�H��%�$�݇�@�PI�*	 ��ף���"H$���\:D*	�]�! 'bTA9E	$��9^��S)�$�w�bH$�ȕ�Bv�A$M���A&�l�]LdI�;��/c�(I�/���*��A$L�_n\5��I�$�Hz<��i3�9t&��ĐI8�ZM�K��I�|ݻ �           �    m۝c�kV����X�u�����+pH���kZ��-��  :s:��9�5��hI�;����H&�˱$D�%�$�P��TO=y�	W/)���A<����M�$NĨ$�z���I���$�k=�IW.�$��J�ؕ�MQBH$���\A9˱$D湿EU�SPI���A$L�%�$��A$MĨ@$@r׆�HP�7P�Q�N��{��\  c��K�������X����ql�����|��@P Ui����U�|�5��@f��|�'Hɝn[RE��rhq$iﶴ�Ma�[��[iw�q����   ���,L̩�2�L�G� ��=[zj����܆�;��/
r��M��9�O'�s��c=��V#�E���]�%���bF"� � �5�`c+ܺl�`ŉ��XƬ	Va%Y�YX���x�%�D��R�Z�8Myg7`�&�j�8�mmA�n{�h>[�(��u���9f��>�[�ĵC��G�'1��cS��5�%ɡ�E�k�nr~    Peq�B���wu׵�-�*y?5ֻU�rh���Q�,B����4�
�qg�7P�u�)�XG�
 n�>؊��[�.�4$Ӣx�^���l���  M��d��b\�b�X��$a�/qh��] ��q1Q�54D�y1�+}�=Q3�>e�>�j�"�~nd̠3�3�X�ZWZz֟7ߛ�[i$               6��z#��m���m�qV�hN��VPgHon8�z�:w�N�|�>m� yIK��.�˱]�0�#��T~�z
e�E�Y��W_��܀�C�F�^�(�wVJ��0��������;�|���>[��  ��ț��W2i�5E3~��^��Y��.����Qddϛ��#u�Gځ#~��*d�C�E����+�汯ˑ/z,ɨ�~�'�    4R2�`
K8��H���Lc@�K�Ru_����0��4�hf����j"+.ГYcSFG�q�܆b��y�,�@��;�i2���$ ����J���[;k����V�#�GH����^X�Q�q1i�k�S)Ƒ&L���ʍ�����9GƮ�<��̼P��^ixuFw^��r�T�����%���N�    %l�d�.KE�2�Q�Qdi���l�f4�$�.��]擑�
k��FL�����^*2t��$���S�Y;�$�9{��WQ&!(�P1�w��}����}��              �E��v�
w_�7LNYnMz�6��2��  W74:#a%��>����Eڎ��	5CHP�Qf�M5�\��h{�z��ѡ�(�4�v���1X�u�����w�]����    &�YG�J��~io�fMq���m�n^���D8��CH�|
e��Qt���ӏ	L�D�3����T�mcJ��5���?7�t   x���-�\�|￻�{lf��Imv��������#~���G��&�ݔ�W�;��L]ьT��|��U�
�3J��7��6��j���׽4��n`    �-)]Xr�v�&�ر�ި�e��)���%d�7Tz��ˡ�	��3��4-/�9H冱q���D��~v=��*�ر�����L     i�Y%r���UfMq�y���&o���t4�6���-;y��m܅ڎ�0��kAL�Zn�ȓ� n�ӏIM'�}h;��4?��x7c�w2��##è��F��1��Q��P����T%icH�	BB�P�C
��!K(#Eboj�.��]����J&���I  8  6�                                                                          p vL�g]5V��t�1�7D�<5�i/l�:�rK5���ݶ�mlh�2�.�6�my�Kݢ��d�:�*�]�X��,���ƵnY�:SY��]���|m�K�l�i�F�j[��^V�U�5���˻���k���m��5bn�I�9z4�mΒ�w��5W�ל���R!�x����z%�k�$����             6�r��c�jk����e�ԝ�jM�Bty7KI鶞ɵ�w�/���նo�    ��d�J��wk�|�9<��0�!T��r��](�C	�������1"��P����-k@�B�C9��6����"̕��/>NL    4QB��-�m�Ȼ�~cH�|
mP�A `�  ��CH�?zJi?{��r�Q�nh)��Yi��tDU5��B@w!t��A��ϟ90    �
F��KiJbX43Tf!�bOP��D���c��笲�i�}�(
 �n���C����� ����:/��o�M��
� f!�1i�33-� ���Q�*��K�ȶ��C1GNނ�t4� k����R^j[��<���z�9�C���b'L� �26��Ʀ�sP��@w!��~�~�o��@ ����L��K�YV4�w���;�꿛���\sw!�|C[\
mP�P��b�zJi8�TI�;�z�=}�
e�◸�W�5���ӭ�m� m               m�-����RiN�����/k��v�4�ĭ�p����w��{�� ��Һl�e���)Y�2�oN�ՃX.��Dd�Z�Ƽ�X�џ����O���^��t>�b�7Pʯ���uW����t���~�@ )#2��Ī�Sk0�J/`�Hwk�S)��'�Ob'
R�J����aT�R$T��
e�ER� ��-p�r� �|5�v7V��y��{�տ��  r�6����3�F�j&��T#n��Q��Uks&L�*�J� BP#��Bl�)�C�;�f��$(Gy�u�u܉6�"�&���:     �B� NWv�������kIkq{�U���$�͘�@U�寅0hf!�uiI��94dI��`Q�c���0U+5�ˡ�ln��C�(빐 ?�׽*k���V�ӻ���ڎ�p	>ʠSj��?�'Tú����*e9��#u�N^�t0�T��(�J�yz�K2(Y�j�}S}�$ J             ������
���$�G]��z�mwL�t��ŷ��������_@ -̺Y\�-H�����Q[�SFc5�B�"&��ˡH^*"�U��d�&�n���0ՌҢ�@&�
�5�  X����K�������$WVd��TТl��r)؇Ʃ.�܃�	�QZ����Eڊ��3��ٹ�]7�� �;mu�K6ktt"���Fb�~n�#�=�+w = D���SaP�B��] E�/�u�R�;&.������6ٳqыB�$��/S�f�biL�[��Q�>���\;��.�L�%��#J�����@�z�)F���&S͓�xJe8�@q��F�;z
e�	6��_>|���gϟ� ��]!əjD� w �܄k�6S��� � O�d᭔f7P�wP�Q5׍&].��C^4u��ߛ��܇�*����{t��~/��  r�a�Xrٵ�5�ů��_��ܮ]fO��3zv�ˡ(f(�A�^r~ w!���9!Z��%P�QX�3v����<��������ɷ�[@             v��n5�-�J��J���å��'MM-���9w����z��  	6kn���6�h������3Mz�ˡ$
Hf(�C�^nC n�6�ux�^��Sj��x�_"��q�\�̋Y�����_o�  -�Н �
+9]�m �����Bi/3�d�~� 	`k������X&�=�7V�W�MD@��q�x����_^4�t��ްuG���߳���  Ng6�g2܆a��*�n�" ��%m�)�C�p������@�[��)��@�$@tp�Sb�G�W��X�� �T��s�����H�=冒�����33  I�-��&֮�����_H4A�/�&��r��3 E_�ZNT�3h=Qv���܆b���Qԃ�$�� ["a��/AneP�Pr؏�/{'���  e�Sv�IL��;��b����	�4t�r��$φ������	Z�J��i@� F,J��xrh�W!���}�����O�h             n��淴�2q��٪��޻�X���JttԻ�g���  r�#K	��kt���=��ܢ����2�j7P��������A�=�>%2�����C1|A��S�ݡ�I�r*���    ���N���Q+"Y�Rk2-K�9J�b���T� ��#5k<54f6�.�b��j�ˠHf(&�/���ifDrk2%�p}~�    @l�%�meݪmfO�w"]�
�>��ĦS�x�(�j����4����w*H�DC�掅������S�jTn�(�[\1�T3���D��V�_� �L�^$;T�NZCI�#u���˨5hn��C�^nC n�6��r<��tˡ����� ���=ʚ�<%2�n���|���>|�@ ̵��!���T����#c<�*Y�R7P��py)*������/��3�#vX�1�>�i2�D���ġ�H;��d�,���E8���b�Ȑd!�HՌl�DH�ABF0  �]J��U 2ڐ��	�������|�[&`��8  6�                                                  ��                      p ]��-i��s�k�,��۷nI�γ��r�WI)'d�U���6��RK��k��6����y{r�Ӻ4�[ź��T��Clp��h� �vM�kN�վ[dη^ܒNx�:�e�k�[*�!Xݶf�j�X�"Ź���-��]wE^7V�I��q��9z\A�����O��8�VpXe �=*#TL�s��!��%���m�             �:[Ֆ��ʦ�v�����fܫ�N�T+�]��=�zֶ��=�@ ��^�������;���Q�B�pˡ����L�k�T̹@m����y�
e�4��2�~k��}(���ݨ[����K��7�  -�颸�\�}￻�W��f(��rh�w!m�R�� ��f��t"i�huW���w3*�Gr}�'+�]�K��\�_s��     ��"+���K��������QUw��]Dzi���������!�PiV�H����U�X��r�UB�	5�C��������f(ʟ��}  u�k���Ɠ!Љ�c1Fb��r�t�uz�(w]��N��mK� ����h�����.�me�	����)�B�'���>^��ߟ� �	��,Ȃk3�W[z�'�)&�5�MsP��ȿ��Fcm@�����i2�D��n���rue��_|{�� h              %�nn���puFV���-&�wW����v ]U@  ��(��'+�^��;�I�����SI�r�5Yį�Q��2�r�ꋴ�NH�L��C��|��mfMb\�V�ع�>�     n��,�Q��Q*��"�d\�ez�ˡ�8�hh�kA�=5��dՇ-���/gAM'Cu�������q���� ��f(�s���  x�]Mڙڝ..�9Cuq�U���܄ʍ� �^�*�+� 	� t����L)�Ҵ�:�ڇ^�i2�G�ln��lb�i�� әͦ��Sgiù���5�2�j�3/vzrAL5�Wuߧ+L�@���c���99=�?��ϯ��_�  �mon�6�S�-ٱ�j�ᩅ����U�Ɠ/��M�9�zݺ����'��L�꼻c�r}{��y��O��h             nܺ��^I�e�;j�Q��v��0lӭ�N����[�O$���q׻� �RJb��jt�]��g�+L�sx>�N������<:ʥ���ɼ
��p���9����R限 �+K3�F�M�����s��gw@y{S�*AS*o.�]�m�)��g�{�����AL��5��'�*��  u��&��r��.wl�\1�Y��r�_p�ԭ��G�_Tm�=*���P+F`�4 �I��M��R!!�D�b�X`��8@(�`D�#d*m���d҉z��dN�Þ�
��$d��Jݬi>S�{��3�\�{������>O��  �sfeZe��_wfٝ�2�~���{�J��9��ۦv�|��ܧ7f���+�X��".g%|9�U���;6���y��� �"�x��N]g�����w�֓/D�e��U���^uY�N�2�.����ݭ۹Єw�����             m^�3Nyrtn�u,�n�f�%�i,�%q+n[i.���_K�  ��aP:��,�	��/J=Ԫktv �H�){wlj�U�M�ݾv��e��V}�{�흏���   1�*h%)��2܄��޶���S+/��`@�D@Z�=כZ
e���Y��X����y͜ߗ��od��+�0    %WY �	�m�ܙ�{�W]�SGn������ZL��������[�|]�y�� ����ħ)�;�w^�` V��C����C��Þ�Zm������?T�	NN��t�^ĥ��a�>�b+�Q!�zg����ϻ�w��/    0$-�IGZY+�7W{́�)e�N�׹��i)��V]�mX)���������m��s���${�� $               m�HC�j��\�x3_6פ�f��s�5���4���y�OzǾ� $$]�8����=�U/r�d�X�����I�Y��S���+��^.�����Mn���u}y7��  :qt�F�J�ݫ:�3�ـ�^�������_سm�W���~��'�Dw����*��\ə䴓�w�ퟙ�`    ��$�NL�-�M�{��z�����v��Кݫ�$l@s�W4JefU���{�s�ʤ��fs��]}�    +�U�F��{���s|r�2��Ϡ9���)wm`�o��ɣ�c��!� |@Q $����i�rk2���}�� �gi���HA�ݼ��=���W��y�>���L�]�~���[{�Kw�����✚�tU���~�?(~5L>T�*I$�H�F�@.Q���
���RϹ��_�9v���ʊ1���Wl�Y��L�VnQ �#,V��4�E*c�4�@�(�`�0@C�@Z��j*!�H-��E����%�FI	Xm!pj
(� �(I�J�n�$d[�m±L �(LE% ݸX�#�B�����j����M���{3�Zu@U���kQE$$����n�<t�~l/�o�B�2兒�������5��\UФ��*�)9���'�ߨla�c�6g��h��L�b�g����?i��>mDS�'����po��{��rj ��PE>r ?�PB"P�l}?�1����XC�?�b~d��J�{_��DY�_���S���=���@?W�쯉��?��������g~� �C�(����[�7O�Uy��i��O��(l�u��w]I��� �}g������}�̩̑>�P�DEEo!+Cy�}���$�dI"H1��$!�.��b��R���� $���������!"�0���H�"�� 	"�"H�F"�����"0�0�ȉȂ�H
H#�$`��"���"�(��a)$b $ �\V�	(�!��CdI$FE�FDD��DY�P�	�F",B� (��
� ����F����6ШQBT!BAP�T$ET!BDXAP�EBAaBBEdQAaP�Q1A`H�"2@�>�űB����dX��v��}�O��
 ��b�A�U�����@ a d��|�C����?S���>G��h4 ����Tb������T������t'ƽ�u�O�nK�>��?���*�AQTL�|�����{0��#��c�oiS՟�Q�J��,�b�.6���/�m?G�g��=��=̓�~D�~����{������J����@�����>�������S�ß�!�� O��
��� T�/���`)��C�ʔ�,x�uUpxǆ����2��" ����x�	-�����y��
����
Ću	���@Ѡ-�����5 �6��iCKԴ�����1Ay0�=�F9ҝ�C��&T@(�8�����[���*~o���������~{�H�y��K�j�y�i�ޅU���}o���[6C�G�>����/��O�~�}8?tA T�}'���(�c��" 
�H��(�~IG������߿���{�O̾��~	���#�`}�S,(��!l����?�]����Bx~�7cV�n���M���=ǭd�UA�k����Bc�(>.���O���������@��@(�7�>[��M�����������U@�؟�g��Bp��(�Oٗ/t��)��� �O�C���o~���c��?w�8_�C�j��������8���.�p� �?�