BZh91AY&SY�_r��b߀pp���f� ����an? ��A���Ҁ  ��fm�
�N^�P  P@�R� *
                     �                  0   ��*co�O����z�}�J�k���[Mz���3�m������ׯ}����ek��r�W�^��}��  �� �H�5�ΝR�$n�w5B���0���iT��hҶ�P��.�m�
q\L�M�h�6ƀ��:h.R�6tt@�@иJ
�53��t��R����m�zN�۶�U��t��mJv�6�n����M�{��*��7R�;��������;�
D H�����l����^ʮ�ǎ�+�v�isz�W7]u�f�Uvʍ��m�n�Z�i]�U\����wp�A &;�Gj�Gj�ֹ[J�$��*;\=�*;z�WN�x��m]]�U�z����Y�v몍���= ���
@����<u�f�[ۼ��ͻ��T{{��j����sR���{ʮ�uIۮ���z�wHe��� �
,�yI�oZ�osJmZ�:���y�ۀg��*ۮ񴼭�-{V��(��u+�;r��޴v�\��V;ק��pW)�����]���F��{z�y�E��N��Υ��+�/Z��)燥�oeWo ����Qޕv�F���C���YU۴7*�w5Gn��jҸ��U۲7J��Բ�o  �@ @q��Vz��uҮ��U�s�GV���ʹ����W�r�n��ӻ=i��\������@      DS�@���@  �d4 U?*�       ?&�RT�G�  4     ��*HjT�  �  &F?B)���P 4   h �	J0S��444h�<��?�*����O������u�>���{���u��PU~�7��Uv�**��TU��P�������?�������"��_���Uw���Ѐ��������?��s��?����1���֎����x\á�������/pJLL������m���(J��}]�1�DjB�:�pHw	���)��!BrR��(|����Dfm�<��^b�s.M7,��3�����'�ˤ3_w��od��ɪ2q=5mf@nRj��MH\��[�)�&�)JB��7!JR�Hd&JrB��MHP�]�|���Q��Ҡ�Y5ˊ���*>���wǦ���fw��2��2w�A���odLa�83c<;�-O��3�uw�x�L�dbД%)HP���Do/v[�Ƭ�����f�n��᣷s�6�k��qsK���d���P��6jN��*(ѷ�wݝ�R��7!��:z�&z�C#K��#!�ޤ+��������)HR�M&X�Bj��:�"L�����M��f��Q��=��i/MJP��$9	�og��ߜ׾w�~�{燧�=ώ��K�[֤��l��a�Y3�v��rR��D9Np�u�Uw뻼Z�$پ��8w������÷<Lt1��w�!�NJr�[뷐h#"4=C�Ec�I��H�M�8�\r5D���' �"���f�<5	BrS$.i�j:��zk�{�}�콉'�.�h�y�x�В��e���HP��)Bd�!�%O<��1���A�ձ�w�JR�nw�;�ɣ>6}�7ߖW[��;�dH�6�)�6��b|�vw=>��lɾaZMh�M�����%	C������y����q"��	JR%!������n�SQ�1ș�I&:H�~��9���w�Cz4�^N�Pb���Q�<l5�3}�������P4�	�{5�a���*��N��9�1������]�F�A=F�����p�'!2��M�n��)���nȽ�c3/ӿ5��M-`�!2R��;�}³��������N�ϓ�WN���<;�C�L���aK��s��9&C�2\��hrR��Ί��f�Ѹ�[L4hgZd���Y�9�#s%�Z�E8�لl<����v^�|:���v�-�V�����N�_9w��{�w���K����i�:b��l�ቖ�ւ1�k� �� �typzy�/8��o9Y�K&�|�g�t8�y�>C��l����1�o0�]BP�%	BS�E�f>�f�a8Z�̶Z54�X�ۗTε�C!(J��)�c�Ns\;���p�V/Z�*B2L��B͆�Q���a��6�6`p#Zم��-�`��F�q��.F��38g#���q2^&&O`dj��)JR�<u8��h���Z�yᾝo�t�y�p=��Խ�:v�#�Gdj\;�{J,�a��y��~<�Σ������M�K��xjpٮ�s�z�=�4�X��	�oy�PY���pmkf�o��sI�Rj,�G��9'O��N��k�2R��(B��)
:���ԛ#�����]�R��r	��%	��%f���'��G�|-���9цk%�F���t�	2�����(JR�(s^Ju.��"!:(`�.�29Q�����S���eF�t�������Äe��kÁĴZ<#I���:�Y�����{�|Ӑ����̸K�ד��M�2L���hʃP���:��$<�th����s}�vw�3�6��CFl���#�8�o�
+VhGs;�����u�yU���)�ۣ(�b�1�wt��]��da��.X�Ԝ��c9����:������=�{9�JR'r�&�)I�\�'�y��Ӻ=�mì7�x�GAj��ᮦ<Os}<�n�t�
QQ�j����j}olu)��{�Z�%����F�cZ7;"��s����:���e|��T�멜=2�/��ʤ|s�[�d[��ĵ��G7s^u.�=��)JC�:0���L�]G����7��Q-�}W�3�5=�A]4E�f�X˷K�0��u�Ns�>U'�]v���W�"�W�@�P��3��,���ӷ��Ru�2�Z��X�ĘNg����rC2CaPbV�=il��j��������z�����lg��&�|��W��}*Qj}��O
�^��[Ka�N�F�5>��MHP�JRI�sSC&	���r��dړ�!�Bw!���(JR��)J���ɉë���
�+%wٟJ��;�q�ʅS痢9��X�p׎��L�Ðm�睜߄�D�k����ӧ
#W9ã�|��駷s=�7���i�j1�ߦ�A�J�k��7�-Be�PW��_G�:*��+��}�c�� ��8��f��Ǯ����`�[xt���>�[�Eg��9g�"�����~k��:4��8&&^K�V�deL�&�,5��sY�o��;3���֜���8w���F����uгp�c�թ �(�:ߞy����S����ц��\5�nμ�}�f�O7�r��'�f�m�	�hi���ޗ�a���ggh��++3;]�$j{�~j�g��h���#��NBjM&��C"8�cޅ�Y�5�sb�OO~���y��|�'/1<H��c�ϏI?x=��������	JR%)H^o��fn����<c+A�2Y�0���ԥ8A��`�Y���a��M����B�.���J%�X����NS��4NXF�:Xk ւ�Y&f`Tcf��RZ�̲[��F����ڭ�g���:�8͘�%By�cBR��I�d��� �(�{� �8��D�PgZ�R%)HP��!]���U�R�-�/��r���d�!�����ǏV!����!)u`f�5��=�~HrM�)}7tv�j�*cN�-F��$�<����˧7�h#S��7�&�K��[�y�rqr4��C�z��o`hy���%i˺�k$������$�İ�Y4P��X%%���U���j
�vN*j��d%@E,�T�C9b���ְ��	�ZҔF2jR���1��Ʒ���j��� ��k<�l�;�b��e�c�|��>|Г�ڜ��o6�����^��百��A݋EFDWR���5������1��e9����ӎtA�&��������=�WwXgN���(4V�;�fa�ٝ$���z��G�î�B��h�g��C4;Jh�w���!Z���3u�ԘF�A�	[gM��h�o`gz�A�J�AQk�,�05[,���i�Ih��DG��h2w�\r0:�X�'޸���M�>���y�w��g�e���|��#�n�yA���<a9e�~�')������ɖ������=ֶec��oso����s2��[�!��YQX�NC��e�E�dFO	3[�m��1��E&I�d99	�56X0j\�y���t�F�,"Й!BrR��v��^�s��&c�n���.�r���rL�2#3��{!O
���������7��#�wo���W��y��=�6���!�2C �豔���Z��r(���9QE4�	Mq<Ԟn�g[0��{�䑒�'P��{��܌5f�1�S�*��s��⢯eY�t>�@�
$��=w���ơ��������du���$�$��f�.�ALn�Br��g"��a��O���=�
+Ռ �L5hz�	�5��y�u���`i�G:�j�<"ٮe.^���]tp,��Σ�p̀�Y�%@z9=.X�q���;�k�/yoA�\�;h��͋��W��U�ٔ'�1վuto�s�r�Έ�]p�r��s������A�Ѡ�Fu�͝��o~gY]�%uT�\����Q�TGM���p=!�F��u�ZX�6f�!ø_J~����T���T�b��)�QX>$�G�Yk$�TK��Φ�'IJPPw�:�2\##
��F:��㬫17Ԛ'0i	���
)(jwӅLY{)@D�g0no��d�99�l`�d�l�>�Z��莞oBu��;�ݽ�ǝ	BP�%XCd'Z�By!I�������C��:�o$�.I��l|���֞�O[��D�I�L��(fщ�J�(JR��)Jy	a����r�jR� �� ӬB��a�3���	JYO�Z79�ٱ_B��4a������O	�\�h�P��6s7��c��V0NN�xh�E��+��St�1xÓ�J���B8�$�6f�5��I��T%:K%ӓ�e�!������07���Y�0#%��B�A98a�q��5I�q�MM��\�M�Zu�L�I�� �14XFKo5�H[)_�V��5����ߤ�e�[����d�4�Nu����	���n���h�[���Y^}M�aw$��7�Nܔ�,r�'���:
K�çf��NM���^N���C��LL3Z�.F�'y����]Hu�d>�=dޣ�:�✄�r1��|�	Z�,�
9����G��ӿ&l�(�Inh�k���&5�Q�9+5��FZ�5�Nh����͘oQT��CFb��c�"�l78��Ĳ��<�D�Xj�х�p���h���2}��խf����ފ$��zL��n	&t8���<����������?y{�7�����#\M���tx?�ɸcd�}��U�
`�w@ǯ��2i���K�Ʌ��E�����a-I"��������Ǖ��}�w�,���$G��uZ�f�������\Zu�K�-��E��N��V;vڨ�OWS����L��,(�`G=�����5�כ�`��~]����`�6����K�b����H���qd�����N:P<���  �C���s�%�վD���ѡDj˯;��jI�k	Fdof����A����Ӻ){��`����ofC��������|���)�=ݢpA�;�%6�I"��bC�w���V��똟w��l�@��䶉*s��ky�o �:��5x���[H��GC���t:pˠCĀ����(�M��G|wfrc�k�\���)U�` y�Y٫|A�C�s�Q�G�+%"��$DO%�*.��Q�,�p^\�+�r�x�P=v��4֧�jꑺ�E�q*� +�;ϔjHa�$�� I�<�S�آ��j�C���t:t:� �C���t:�d��$����C���t?����t?����t:�C��輭t:�C���t:�C���t:�C���w���t:�C��-�I-�@�t:�C���t:�C���w0:�C��r�C���t:-��C�[D��-�@�t:�C��&��4H�E��C��$�4H��(�Kh�Kh�:�C�����t:�C���t:�l9�	�[D�[D���t:<dP$�C���t:�hv	���-�H�C���t:���C��ΗA���C���t:�C���t:�ht:�C���t:�C���`c%U-��LA��t:��/���|�C���t:�w]�C���t:�C���t:�C��� (�:�C�ѽ�2C���t:�N�$$���:g(t:�mImC���ܐ� p:�C���t:��$��$�C�F�Fղ����t:�C���C��2�uTZ�C���t:�C�Q�d2�>���C���t:���t:�:�C���t:�C��-�I-�@�t:�C���w���Iv[D�[GH]�C����u%��A��t:�C���t:�x:]�����<�z����t:�C���t:�C |�C���t:�C���t;%�H�U�vKh�Kh�:�C���t:�C���t;�?Q TZ[��-� �w���u�����j���t:�C���t:�C���� vB.|-��C��`�H��tJ��t:�C���K�P�v�C��$��:S�?�:5�t:$��R�4:�t:�QyC���.��C!�@�bI��	q�z�����(o�\�w!X�<�*')��¸��'�kQht:+ �J�C��o�:�����|�u�bD�J`�<Cց�@�t3�F]�p��,s�m��kRH-�a�@���9� U�C�U��C�g.��\�I�[�f��_=��1.$�=�7���` n�!���8�9m��a��t:�md�� F��{���a�[zL$� ]���m�.�d�HaDX�H�C�l0�ē�,>b�ƶpK����kw�ͅG��������<�l�q����
q��W��X���H�c���z�&��� t<S5�[�q���>�]ݲx�gx^�[#\s	$;�	5�tFĭ�a��v���/��(�h8~ߴj|Pt8��0H<�t�J�W$�̈G�zz�I�a�'h��(Y��I�BT��%PHH�C��wP�I$�����=�qSL�΅E���t:�C���C�� ���(L�`�FM>0�aA����T�}�l�J�^�D���tk��t:5�$�Psw�V���y��9��I/74�[�D�3�
�V��a��{����C��o�`.ݾ>�zw'�bR-kΛᧁ&{��0V��DZq�v㫍{xV���NIT����HT8��o�nZ$�^��q�$�թ,�N*�n�^G��s�3J�P)`�%�G���ʸ�m��I�ww.گ�MS���o�h  ��k���t:� ���TZ�"��m��C6�m��n���n���(l:��r�rj�I����#՜�cz�)9Qh��;[h&�C���N�F��C��怍g�͹ĺ�HEu~�7|�Y }휈���i�$�C���m�m�C���t:I$�C��� P�t:�C���t:K|�Fl0�Aa��t:�C�wdJ
�pz��}M�-&��(�J�0�y�nhH��Ba��s7���=�:�]6$����06:��O��[�q!Z�d�HR�/#�������v۶����	��rtʴ����Fb?��Oz�����i�ّk���װ��i�$�*7^�]GD�mnH��s�ZJ�o^�'ۑTM��6ǃ)��pV*;�L��R��@��
̺����A�-�
ʨ;�N��RH�Z+0�m��0�d	�`;�r෺n��w�K�	���n�k����yP���i�G���tgA�Z2�cZ���A.|к��I��s;˹	���J����\�v�|�}�*�Sj���F�f3�LKo6I-�9�K-xq0�+ز^O�C�u�������l1����<��$ݭ�	v�NuWy.�@%
c�͆	}9%9$��
�I�� �"�K�$-���po�Q��'�� ��$�C�s[pR]	��\M���l(������LI:,��7bw�0�û8�F�is(�J�̼�(��Q��@`�G3�.�ԻF��P�rL�4٢쪩�m�^���^��,Kg����ָ=o�����b6bbvE��o��e��'��uL��o5�����
������[�K˹�&N/zU�͇�i@��ZI$V�̪79�J�m�FѪ	��b�kcvk�"���d08�I���{�p[l�����嫴"9� ����C�L�t:��7�@�����}�<�-�{{��m#ªUv���ow3;�#1n�ԖRF�&�ԉ������ow!7A;�q;;�a�-���� ��3�I�nf��F���k�N.�=Pڨ2��I���O��u���wwY���t:��0���-�$�I ���$�.g6�8� #� ZKdHx V�D���
i�J7�_.��V\[��@d�J�t͑J�H�	{�Y�5����(No˪N$�2r 2�3;E�O���A�E3�j�UI �+�qo��D���RK�	� ,$n��T� ��w9�h��P��S�v&���3�]Ԓ\��=��<�+-�}��O��7$��� l877r���Z�g��u+�jH  �8�\�����TZI#�X�H�C���t:vK˸�-�C���t:�+����{��b�wwA!������G~W �
�Vۙ��� �ݺ=�d̰Á�]�KA�3��ɐ����p#����Ğo���u��71a������{�F+i{���m9�y�%��t��Ĩ�'1 i'��3�w=�`��&�ѻd:���Q��mc������F����һ܏�X\��
�������w�,Z�b] lZ��Ȣw�c@ē�Ul��c7�v��X*� �`�r����j������'#�#����d��ۍ�l%�$s|c��\_y����~Xd�K�wB�7��[L �޹�4J6�{82>��~����[�nwj��˒�����oqnqO[hw��ǫ�@��.�����ηE��z>�[n6�܀�퀡��⹚/a*�e���π b2si!���ٝ����P�nv�5K(`<��}���K/!�^�t�{��ט�
��tR-��'�H�<�\O�<I�ք;��	nu���O��4�M�m���!S��s}�R`S%�	���F�,z �]k��I@]�PB����]CkH,��<�2�.����O����u�?b����RL��N�'L�  ��i�h��
C�����>��Q�Âͳ`����n�>�|�t����@̭�d�G����:��܂x�{1��-ݶ��C���wRH�x���U��͈��9(�l� �:8M	f޴T��}U��z�;��i)���
f6�E�����0n�b�á��m����׬��c��:^�˄��g<4Mo�\To?X����k����;��3�K��^�ͺ�m�_)�5b� 7̤u���;�z�x��.��/i���h�l$����B�Ɇ}���'@��8�`�[��0g�Gܞ9`�8���s�H�*8R�Ss����"�����\�G���4'::�f��q#��#�ޗ�	=Y!J����I� sjE�/d��A�+��M뇉$b�$�H'�U�t�D�C!�@�t�k�NGB!�:w|�۰j��>�����=C��@LU����$p~�Mԕ�dV�Ƀ�IdK��A�M�Vl,:ō�f9�T�!�Kƒ���L���輆�1�����htX��a��t:�EV�$����t:<���	$S�ڗn܎��]�ͻ͏0��`�>|�a����_>)i`Rh���� N����A�����t: @
��丝�$�΅E���$�d0O��L�w�HZ3s]��{�HQvC
�s��w �@
�'��F��
�^��17@R���0�NKoN�E8��L\$�yBm=N�ز�r�C�U���� � �I�t*-�·C�w_)�|�)��/=Ь\������diA��_$�H��6�tn�@� �M���9&���Ӥ
�<��y�*k�F{�ȟ>G��n�b����ܯ��?�|���w��x����%9��i��1��Z|nD��՜伺��j�� t:.]Y�����)6:� y���ݩRF۠$/��MP ٰ�����$��$,0ݛ�-�I�c��\���;�����<�L��&����t;;{�7(M�g��p&,�X��|n"Gh�1�V�@�6�拻�D^��zVJy+�S�y�x��y�p$w���8�5�7t�6g�@�����	�����T�]��h�{Km��u>�X��5���8� �:�w��w��ڦ�j��iP�t�݈����� D���˙SAt�om���	�C�2���_g��F�I���w�k�v��W�2m�^Vyy{�g��ݿ��-Q���:���t� TY �M��A�j l1�����d7t�(  p�p�$�[�*@#�0r�ʘ���$К5$-��bd�s:��V�����$d���Ix��S�
�I!�%w�?7Ķ)�>qP��W7!'�	���hkI<hT:�s�(�9�C�y �V��٘��@�t:��l�� t:/Z�t:j�^��z����=R;�g��,�\�!$���qB�A�ãKn�'���k����
��}	'0����?G�+�΅E��%[��w��,*/+]�΅E��輋I�U��I$�M�ɰ��T
���t:��O9��$�eI�3p@��#����q�y
ZX�*� >E�`�=�̐��[��OI�I$��ݽΧ_6�N0���q����f�Mj(�U��1k�q|�K��A9o�ZM[�7�N{x���$�#�󣌝ݩ)B���}�ќ�&�`�T��	�x�h�̶h�M��7��D�	{����RU��ׄ��t,L���Y#:{�[��($o�R�	��vk¼?wu��;*���z�-�H>�;t�hj���Ԙ��[\|�({�9�YF)���Y�Q�AݯU�kRJ�gA���6Pbʒ
2@�.]�}������L���`�·C���u�m�<�����vz!&�A�I�I"QP`�$d黲�N)y!`a^�a!!������ھ�v��C���t;�C����Hks<kӮ�O{K�P�t:*Ԓ�7$�jKwE �Di��쑾PZ-�<`�$���=��Ot���\�I29i(�=4�22NCx0�K~�5�]�1��	N��ݏk�\�� �	�J��B~�d����:кNP(r��2N+��A�E�4��s7������I�������Zwqۨ��:s1�5�0 	�A�I�C���t:�C��'Y���Au�š�:H<�|~K�椐�	�|�" ���w]�]�IE��n�U��5IT%�1���t:��E�Հ5>}�H�0�t>��,%��H�jIuuZ�̜�t:�r���t:�a�þ�����t:�ڭ7I')_)�����>\9�t:�C���$����H6.���n�ݼ��r6���m���;��<构ܭ$��-X���᫻��i#	��0� \�b�l8��v�+����Ĉġ��^�R6$��]3�.�9�3�x��xJ���wك���4
w��%�P�f�Z���/{ٵ��:z&�����X�]c�o����I��$=�^�IȤ�s�^%ý�M�}Ǡ��6�ښµ��VFR��3 t:l0��"�aI=�L  ��ۗqy�F�tzH&��:i�8�ն�:�wC����	?5�?����t3�K��Gfs�C���t:�_6ݞ���A�Kq���t^V��C���u�m��w��h�53�\�t�'@H:�I\����ٖ׻�:���C�ĳJ���I���
����i��j��}�%� ��]ʏ�h82HJnY�Sׂk��\����QQ?����AP���_��Q�������߯��lMUd�?�?�0?�8�������h*(����Ң!�?���S�EM/jt ����L�R%T1"P�4l6����O���h �"���fP;�TR =�)ڀ����T�08vw��1.	3;�Ј>� ��E48���A+j h
.��D�;PG���P�$	M�.�=@;D=T �6��Ю�$��x
�U�/�EdE<�$±R�)4�$�RJ�JB�$K1��N�v��!��DBX9�2��� �4��@�A�`8U��*&@e�:PN�|�JJ���	B�g3(&���>�QB�d�dI�I!�$%TzM,�R�H�K�b�����X_ 8v ��@p�Y@��8�&�C�C�5�!�_����i�6��(XT;�@l�pI ��=b��0+��F ��TWK����������?���������x*��a
�b@��%J�����*��������3��t�j6S����U'Q`M�h�.�eB�5PU�t
�κ˖�WJ� T�u��Uq@�kUFl���n֓.������R�V��f���-y ɢ&.�lq,�We 6�\EjF恜�#R)b�t�a��FQ�z��r�mg�i����]��f���t5�V�r��6x�j�m��Ar�e���^T�V�׫�:�Y4W]��ڸ�ݸ��Ҽ��}Ps�xa�Ì�F���%�um,k(��%���+��,�빂5�ݣۜ#�vV͚+!����@l�<��T��#UG�! #��o �]��-�S+�L����#Q�Zs ��ڨ\�
��4�3f.ڂ�67o{7Yf��o?�"iC�+��� q?�U1�� W�A�x+&�N2������Rl�5��.
�q@M#4���é��HD�N�3h 8��д���0v���t�J�j:�ؓY�7k5՗��
�<�i!�B2���.$>a�>��փ��؃>�n��.��Y�RG�ʎ�KI][/{��o��@ϽP�<P7��7�)8�[J7B��yw��>��`g�OZ�y��߻C^��n�H�8�{&ӹ���=��f-y)��:�*F����N��g{<Xr�MH���T�Z�q4T֢��F:P�F��/{�|��a�vx����K�(���,��p�r�iG�M+�b�I�1QM������u�������~��m�u��%���h}�[Ѽ�ܫ����b���
���{�G���`{�^����2�Ե�㌗����‷ú��}�|�ڥ�8v�MA����v�T7tӒ�g]w��=)��ů%=��짱zNݣ�;۠�$�"����V��btt��r%��� t�n7]��xْ���]�Wf7��ů%=�˻�h��{�QQqLD��Ld�1����]�~����論�~=h3�Ow��	�,�Tv(:�g��@^ƝN������w3�<G4�-;�TN�b��v���Z��s�U*��gg���>�},3���dr�v1D�T&���U"�O�E _>�@^�W��?��u!wvGc������&���C6MR1�(��iCgf���g���߳���۾�;�����5��M�%�wt�F�,�c�e@�9kZ��v�^�M�u8^t�@c��P7w���DI��+�FԒ�3���Aߟ���.��gݕ�Ew�]� ݷ-�ht�8��m��7��gr�:���^8z��[n��2B��}�; �/z�g{+֎�U]b%R)A8(7!��*�S],�nh�q���i\���۱�nz�Э�X���3��t��/tU��дY�46b✺T����mWK��Ʈ�i��6(��V;#m'mL��v�c[�֋���+�Dt����0:Se�+�L^|��{ﯻ���y��JD�.夔��.}�^�E!.%�>K�����Wh&��%NJ��w��wν�a���aT��v+�-��94ڶ��F�P��~~>�����O����{���ד=N6�lw{x��;�\�s2M��cpz��Z�vt]o̕�\M
�偞��`�NѼ��O��},�IS210�L%@��@_l�S�f�u8��a^��%)Y%�ƭDp��;�a�9%���6��bVK.b��m@LHR�T�H菑O����{�ŀg��h��$��r:�r_%���M��Ŷ)�+�˷lj���v�L�j��0�:��i�6��Bq��Tp`15��$���0�9�����@^����.�ݝtB7U�J �K ��4�:�;�`g��`g{+֊���ߜ�d�w*�tD�!���^���ޖTᏧ*����Ϻн9+i���r����Z{�ә��p�cג��Wws�n��$ ���{��N�-��y�@fl�Z+�Q��%*�Yt��Ɲ�ξ�X�KBmԚ��3���$fPD�	�#cp�QJrg{�=�^�y��ý^�U����@Q��Ri��\9G'm�7��� �ޚ�e�|�\ޖT�О\$*=:w�;v����~�'%��$�����3`�����g�]sV7����`�;��������|4hi���z�z��/z��ި-�a/GQ�.��bV�(Z}�^�}�K ���X�;�gOt)?(��w%�u%+��vx�.��LIS��RA�F�	bA��2�)�RKlF�z��{2�ى�|s-��w0��h���派SY�mƈ�%��/�z�/vx�;6[�����r��i�T�wb⒣v/���g�w��=����vW�����R��wn�9sdk����������k��I�uUUL�W��f�ia�����n� �H�x�c�v����3̔�b�����5�#Hc�[R�FX����B���B{t&gN��Z���ԉ�LkD�����ϗ��{�V�^�����F8ӱک�qq�j��b8�-%W0����?}�(͖�p��~L�7�p�)�nʒDwrX�6�NT��]����x�3ݕ�A���[3�S���
�v��&���9���g��e���: ~R�)Kwq6���ٵIw��`w�������d�r�D�m��l� B:v�b��9�/V�<�Ѷ��6ys����
�DI�T[P+k�2�Y�Sj"�[�Ѓ���������K�N��\h��*iCE���L�m؃K�vI���c�j=�Vv)gلP�4�9d���_9ʪ;������/�V[�6;�`y|w���ټ���h��roDt�H��P#T�:<����{����ߺY����� v�:Ж����%��"��䎑`{�������w3�N�G���s6w^�� #{�PTK�P^��S���>�}�A�3܍�U���M���^���A�w2�O�f=wi�����f������5j"�F�s�K���`}핶�;�^�o+��_o�K
��=�������M���?�n�wRt�.12jЩ����/Z���!�
��߽:�W}l3ݕ�Ew��~s��v���s�a�eE���D��Q+����9m�Y�df���#�rn��#���l��I�]=��wx�u�=����,e�C�ƴl��r3��=��v3��\� tux�:�L���?� ���p���/v[���w�v��+i���r�=���s��8���v�}��m�����}���҅9N�E)�E4���u8voSP�oT����n�k�(Jv��І�mXo*������(��s���˯%='[��7����9{�>���f1�w)�D4�@�E�)�z�mk^�E�;m���s�9O�yμ7û437���`��5��˞�F�N�[��=��>R��;Jvp��&��y�|z�<��U�X@� N ��Q���v���{6���`{�n٣3�9O�9{�n���e�m��P7��I'7��|�){�<c��VQ��i��v��Qf�Xϟ?~���a��nn�i i�[a��cF�q��������w9'�y�i��/x��~�N�G��9q�ֈEyLjу�o���>Of\�N��/z獲�_=�7�xp��0g�~5�+:盷�_{����9K=���A���6;�]yy��y�~��8�u�h�}<ޠ(&�4a!�Q2b��DI�G��M��G���D�K�z07�pA2
C' ���X���N�I-��kN��5�pI�y��9�٦�Z���4oy�r�q�h'I��0�,Vb�1-Jb�D0!�1������W��zq�
J"%�	Ie���1 �$�y�3F�Gl�(Q�b+��b6h��!���:M��`�д���A���Zh����$'
�����l��n6�¡�
��5�K=C�u(,��K�X���޽3؞|���)����ח:�
�f��á���P�m�:�bVڽi�ֻb� ��M�ffm�ffeY�4��g�%˚e�ʳ������t�33m�3#���Bf�f�f6s!1�q������˥��^��2�Y�.���i����v��\���O���2�����ݺ)�+t	]*L�b�eQa��ʮ�*ܦ�Y�嵡�>�uc%�n'q�(^��!h��ݼ�D\�V���Z�wf�lݵ�k�ؠ�Z3mnI�\fnۗl���K��^���Y]!�z�E�0��i�����x�����8�&�y�H�ضWK`��ؙ��&*��v����w1��rj��q�ӭ�I�Jjs�$��u���9�,���u��.�.��n����>9�x����/%�ˇ�,N8�)�t���mv��fj�!�;Z-��4F2�![Ce
�d��\���p�f�[��fw)���X��9sl�6�$����������k��\a�v�c�іֵ��I���e�"��Rn:v�82�]g���'4:t:��$Zx��9��i��4"騅��˕�7@I�m��e!�Hj�V��k��4��敦���),�*�I��Z�X:VI2��r�G���4��o
V�P�������e̫1����6��;�-U6u����s�}�X�q�����>Gj?�'J��]*�z~��(���
��^B����'c��S��wo�&JR~�翸=JS�y��)���Iz+���;95�%��{�?{��JR�Ͼ��):��}�P�����9�EUw{�Z�iƝ��3'�l��XUp+�����r�U���V�/c9�-q��W^�L��Fo,��Yǿ|���JR�����JR��<��؝BSw�gƾ,�|������P�-��6�+�R�k[�9	I�{�����߷�� i<��}�����/?k��Д�~߳y������ʘ�r;�Ü��(�}��	��=y�pz��<�����@�wz�uUa�Ps�%�i���v����U�R����4{�P��~{��b�	I�~������߶}�2C�*�{h��K��qբA�.�r����~��	JRu�=��JR��u��%�ry��Y7��;/�D�+�R����k��P�*q�T���s�vk���n;\q���LUDr�0��6��bf\ۦ��]@-ғ9�m�ey�����Z-�V��z^�l��t���8�v�m�]i*�3$N�����ۈcDo
����Q�����eͨ��;G�+���?�*�n�
��$�ꨍ�^��e�(>�^���%!�����=�6<F	����@n�IN3�:��=���W/�;�\�g�~9ʬ��{�Ԥ��˸!A�F��;�a]!����-�����r[�O�����JR��}��؝BR���~�w)I��~���R���n��Z�g ַ�B]���u�g9A\���NV�9]�mڔ�'^}�߰:��<�-{�)�����Xr��Q�]��«�\;����2������JR������R�=�����Jo�r��5��p���[��\P��w�����u��2��<�Iԥ)����`���y�7�q8���^GY$2���V�r��k߰MJQ�C8t��ozް�٭�7<��.ۤ
���79�co7�ٮ�|�_~��R��﷿�2R����uUa�Ps��G��F��Tm]s���R$ 	�޷�TKc\��ӭ�m��g39Bm-6�]�h���#�+�v��x��j�ɠ�O����6�6��:��%�:a�NNN}���^�-�2ܻb�"Sg��[~��r[9��h���)K�s_}�j���׿buB]���!�~�k�Y�5�Yǩ5���f����u)Jy�{����'%);���~����=���u	I�~h��N�9l�g���̬;$���;��g&�h:��}�'R��~��4%)C߿h�UXs��j{��L�W}��'*�$�[�k�쵭�z��.��[�%(z�϶}R�����k�R��y���N�9-��>�=�{$��:�;w�������؝@��Q�:��2�޷��5��ͤż�K��=h˵eY�ٮ�=����d�{�߰:��r���S�Pr���#���+�����}����^�uΛ6o��%)w�}��%'���~�����u�����=���	O��Vf�J��)q�whU/���Pr���ZQ�~!��lAv&�>�Z��	�����`�)Jw���	��C߿}�H��u�+2�c����V�r����pBP��}��R���5��&���u�W+r��݋P�t��SNҶַl��) ���{y��?Aԥ)�}�o�&JRu���:��<�}ϸ�^I����u;�,���<{E��O%)N��[��)J-s3z�ff<��Ya��lК*���
]@�7����]��������j��)�J����XUp+��(�R�q���Zwup	�zg1fIrsFkQ�C�r���׿bu)Jw����	JRyw�>��JS�����d����5}����S��&<��0�(9����ҹHR������JR������)I�j{���Ky���=\��{$���θ&JP��{��N�hK�s︦����ZV!D�J�@�Ep��G�;���G�`u)�n�ۥ\��W}�V�V�q�u�)j�s�[�pz��ʈ�'�����r��~������{o�L��FA��:�˕�9Aþ��BwUW#v�u��R��w�������9�Voy�6�fV�4� �M���P��$��}����g9A\�ۻu̔�/>�}�	����_�n�I�掉�wU�J�˙Y���s6�Mo5�����R���~��)JO.���:��<�}��)������N�h���~=��=��:ڲ���,��O>�ݿAԥ)ߞ�X%)I�k�z��;ϯ~⟁-�}�_�߭�o[���g9�ٮ��'P4%�����&�h=��{�P���{��b�%'�~a�؞^r[/����QW�K޹=M�ɠh;��~��)J{����)JN��מ�O,�E������"�,˔@�f6�TL�b�pF�	i���յJ�WC�ue{����T0ф0J�6�&I�u&���8jn����]�n�ÒK�u���	͖�r<j�N3��m<e�:�c��s�\�4C��������p,��	R��#��9�������j���m5�r�Uݺk<e�a�U������t�/9-�F6���Y� ��q<m�Z6�YukCK��F����5�؞�R������)I�����O/9-����gd�ޣ	�f7�#Ν�N���mS��~�)<���=JR�g��qM@�w���N�)O|׻�X%!מ����3yK�9JL�YRe�\¹A�W��W%'���~����>���&�i;��{�'R �ɿ~������g �s\9��sz�	JR~��~�����w��h���d��{��bu)J{����	��[�}M�'��ɒ�!��wU�9T��k߳�R��w��~��JS�=��L��
NI����?}[��k{�vH,�Sfn�N[�������Kd�y��.�U.�k�\(\��ձU	���:�uk�sϾ���%)I�k�z��>�����(����;<���rC�;o�hMs/9]�l���tV�;xɤ%�gx����eJ^����[�j�r1`�p�n�����&F�]41�ld���9ʷ�n�d�y�K-��7����ӆ���O hO3�^��j�����bu)J{������� �5�����V������uT��t�{���9	I�{��ҙ)��5��R���{�߰:��/<���S��5_o�~Q�Rr���'���.r��(������`��'�~g�bu!�TT�L���߿qM@�}�>��ԥ>����9��M׮N���9-���^rsI߾���=BR�}�{�b�	I�k߱:����k�MHw��sY��oyǨ:��u�o:͙��R��<�o�#��ù���m�vm�`��W����Y�U�"����s�������	�߷���~{�ǩJ~�}�c���H���A�,4Z��5�7�ٮ�9uβ3\����t}��JS������%'^y�ߡL���	��ow�$<���S�u#�Õ�o#�����9A�W��s�z��Y �De��'��JO��ï�R���������JO<�߸=@���!XW'�O�D�LӨc����N['��}��JS��^��	H�����Ta�>��}��JR���߱MEV}�M����7w1�9-�*�H����%	�(T|����)�4y�_~��R���kﵡ)T�2��- 44r�7ʷ��a\��V��
S�5uTԵZ�7����y���N�iw���+4�&�KDm(*`[���r�[ՙ�f���qP� D�$�,By�����%)I���?~��P9����|�*��щ�E��q���<�ˋ{.�ͳ����䟂�a� ��宷��;��/}�}�ԥ'_y����JS����?L�������>��ԥ?{���Ʒ�J���mIE�K�Ps��=��U�?���J}�~��%2�Ͼ�o�'P4'}�����$=��ۏ۹��oY�=A�9�k����q:��?g���z����4{�'P=A�	�w){�s��JN��ݟIԥ7g�}�,��9�o|�p�+| C�{��~��R����~�)JRu{���ԥ)�����?�G*����~�+�9Yy`��i�8=JR�y��8�_ǭ��3y�f�c9�ګ��ڝc�p�U�Xl޷��_�o�?��R�g�~��	JR{ߚ���)���|e�7��3w]�Ժ�!bm����Uֺ3z���);��}~���~��L������؝JR���}���PUW��׶���Ô��Fe؜򺔡<�>ϸ��5)A߾���u)J{����	JRyw����?�a���{��ˆ/d�*\u�p���O|�G߰:��/<�}�	�T��w��o�=JR�~����:>�=�����޷é9�h�u[�F�JW�)��5��	�JN����Cԥ)�y�o�L���Д d�L�F ��JR�I�#C��[Z%�h�� [)�����;�y�2Tj�m�#�<���9�H����AQ�&miRd�2i�Lc�����l�gl��'���V�)ݳ�p:8�й����X\�W5M��' ��['l���>������[�y����y'�}�g�:�o�a���uT\�n��I�u�r����^�\¹AUS3���A2Hv̜���u�b��z��z�pTP�~���)�JO���߱:��/<�~⚐��,��Y��7Ǩ3}k� ���f��Ì��E[��y8BH�*����r�rN�)O?f�~�	JR{ߺ>��JS��}��#L�(@�);��}~����䑿�T�WUI�R��ҹu�G9@�y��>���,�DHP!E00@2�9)��߸qJR��s��~��JS����`?��F !(()��$��dYI%�H��P܇�?|k_��L�Xr���ʒIu�9�r�y=����JN��G��u)Jw�k�BR���^�a\��������U9)�uv�o.)�$������H��S���DA 	 �I������@О翳������'R�?� BJjd�@"h}��}���}���5�kz�k�Ruu�4h�o�38�BR����pG%��NI$$皬͖�%m�s)�L����q��|�8T������O`hK�s_�`����}�[��r���\R�d��Sk�J�:��s��F)�z03������]yæ:٢J79��Jf*��ld`��H p�پzh6`�q,�H�3(0��`�Yl �ɱ8hݮm��p�.0�ֈ,�06�Ύh����4��IxF|�˘�çyee%ނL;n��:�WV��ZUd�G�I�E�$E�����twӧ�C�vp��< �ѡX�	�JlcRP��9�+:���n�JPL]Z
@��;F6)Ckm>pPU�uPJĊ�ڳ�[f%���E�5uIZ:���C�u�@��n��c���(du�R��1�Y⎉^��v�jΞ�7ՎRNs��.�.B�um���!�GVd�nu���
�.�jy9,�n�oF�����کV�nr㚭t
ؑbh��v��i�L���97M��I�lI��@���5�D��3��պ�r���n�mٚc	�S��ُ��%n�Mfn*��<n4`J�6��7���Lc��C��Lm�=�2���
���y�j��R0�lV�M���t�yt3lu�E��(mX�M�CW Ͷ� ��4��6�fݺ�mQ����^����s���������	A�GH|�:��A6���n���B�
�=�^���ma�l����cd�a����N����J���B���X��1��T��Ÿ�.AlZ2�2���%S_���o��;��#9���46pl1u᙭Lo�?�NId��g���7oy�)JO���?��:��;�F��ԥ'~��~�?#+ܥ)�{k��#9U�����B��R���K�]VJS�>�|%?!
d�'�����z��>�ֿ~�5	I��k߱:���<�_A�\��u��:1�y�Y9o'�>���u)Jw�k�BR�W$���>��ԥ	���p@u��sY��oyǨ:��Z�u��N�hD�<׿oBR��y��>��JS�}���G�}y��Y<�r����&m��sZ=�������=��ԥ��g5�Zִk�Z��ck�sn��\e� �a��7�S�H�y�ߵ�)J~�G��JR���_}�5!���F�޷�dwXr�-%B�2���H�B�q0{3�'����Eo�ܥ)������`f��nW������J���@�n]�.$����/��3y⍪
>L3�٭��-�:	�J��DF.���8�
��S0S�c�]#�����
x��G۬�y��^~��u���߷�蒫��r���S;��ɷ�R'�.٘)q�#Ϋ����ey߾��R+�IB�����a������|��Jqƭ�Z��tK ����&w����W�}��*�;���@���c�{�?s/��������n�b���f���`T��aV���֌���pA���9wc����#W��JYS�b�v��	��{_��=�(���U$/ImJ�r�_��
�*���o�a��E{�������o�}��w�~��^��W�-Zq��.]%��/ �s�_���J��k��̈́���4�M[�`����o�0Zn�����9�Љ����V!��ER
Z� `��E��BeAJ���οt�V���;�E{�(�˗�\�(�a�UBb)��~�W���߷�^g�g���T?��~��Ѻ�j�H���r�7)F; ϗ��-{�7�q
�Wh�k�-�s1��r:�p��h9{��|������W`k���x�2hi"ʫ��r�88�(���ƍ �7+כ��ӕ@_l�p�YS|�xo������]�_�?J�%���9,�g��W~��sUuߟ}Ϊ��v}�G�#������Țx��E*7��_�~v�ey\~��o���^������_LC�EI��7��Y̿ ʿ�D�]{�}���[����g�|���e5
C������y��#�m��0g;iz�g���5nt,�3)�wd=M�j�Q�0�H��[��ШluFef�uc��l�S��B=:'/s�wdф]6��4�+m�&jRE�ve��1��ě�r��	Xrrs�������I�>���w�]�����ff��]d�VB�R��Ҷ��s���0�����1��R��ӻOZ�oVkfk[��
 �O�}�����~v��^�ei�7ST�V�%7E+����
�f��*�Gaz[�}�]U�����]�g�b�`FP'�<������_���"�<�w$��s߸�$��]�����?}��0=���*�9��\9\^�j�܄nۗH*%܊������R�K*s�w�q�9��%K&Sly��+�T��W�f�e+���?�\���f���V�n����p�Ij�tℴ�z���.�1�v���e�!s�^h�KY�V�����翽;i��[�����l�wvF
�m����/���l�!&]۬s֭bq�9杸��:K��m%幫�k\8�C���g�K�N�\7�WQ87�Sl��<��Nͱh����3^q*S�\q�C$�L�>�J�A���� ��|�7�����O�p!����Iw-+v�Jv�ϻ�xUU������׸��}��6�k��I\�㻼��o/V>���r�=�|��������P�uc;Z�Z��N��-;C.��}�Η{�`���5Ҹ<��o�x�������Tym�e�K�fV�m�v�(Kn,2-�&i���V�H�'J�#M�N���{۵�<������g��ҭc����W�%D��m�0�X���{\7��w߹+�3�*��ԯ��P^rx�M$��-���9`}��^�mUr��R
R��uΩû�[_�����g�'#Υ8�v�V�)I�v~���}�M,��U/ꢟ��_�������l�驥��ȱ*)��]���P�Ε�b�E�>��R��~�؍կ�F%NX�LN���}�{r�d��c�J��4�l�I�s�,�������}�����wx�8j���9J(7�Hțj�BǓ�eEEfB��(�b��㑩`j���۹�j��� @H�n��>�ߺ�x_�?~7����m�r��}���%*�|�0�~�����[X�§3��U������R7�{f���{qڪ	���_�&�P! ���	�{�:��W�������"�>2ٜ�s|�ַ�ծW��(0�J�"����@�^�3���U�������?3}��y?��B<�i��"���۔��+ �_�XZ��L�I)6�OVR�j��Ʈ��Ob�{pֶ_��D`D A�X�>��jU�8$��N�ܦ��2xS*�z���-�7WT7%%����zQ HQ R�����i�z��&�1{޻�䦘|O��>�J�F{�ڨr	��KV�tf�}�}���)�X!F��To�\�߽_�ν�(�T��33~io��b�Uߏ���m)V;��wh?/{ߦ�1?*���������(w��{�r�枝�����Tާ���uW����������CR��{9�Ͽg�Q#�ڀ4[riPhb��$,Ɔ��Z�0I�\g�xY���:��K�j$�mP9�2��׶�������^2�Y��u���JY�t*rZ�����=��cp��rm�4e��V�5�5�oUk3v�{�%�T?���_��w��u��6�ĮI6�&�ﻷ���{�Zc.�f\�F��J�)��R�T�G%�'��V������{m���a��Jy��X�mJLı�erGd�vw��ym��ht�+���ʙ��n�G9
b$"e�`�"�g���?�W9I^�������g)e^��f����<�zf%�&˺h��"� �:�@^��S@|��w^�V��NZ�Z��9%��[���O�U}�H�>l~���	X;����Q+0>���A8�Ƙ�dNT�%y�t�5�N��m�#@'ss�ݚ�[��=ٻ��[턊&).���^\��T���Ury����[Aբ��e�U;����\r�Mlr�/}`��f�T�nϗ�x)s�4=bz6�+�c���-( \t�Z�a���qQ�J�9I�8%�Tn�Ԣ���W�wt�����}����w"�^�<�0��|����\�W?U*�@^���{�ާ|�S~gf~o?��-=;S�9��}����1�%6.��Gk�Эi��Z�ɕ.��ԫ����(]>=n�Ω�7�7�7�����j�ү�(�w���'-��^�`���e^ߚԍ��FJ7^��F���'�{vh��n0�wV�;�דZ�o&K���b|�H��J������ع�"����������)\���e
��D�DÔ�R�����w����J����p���Mk4�f6bkLDLDQ32o��f�.����t� ��k�5�R?{��4�G8`�d2ˊfW�/S�?o)��|����[���R�pwtB�}�Vf����f˛��W�@�D_O�[��Kz�7u+�3T��1%#"[V�<�����Y�}��`+J+��7����0�
rn���[Uf�ݬ�������{�$P���߶?'�8c�6�!&�aɚx��˷nK�B!s�K9��0@��<�>��e�3���̀j�_��E~�ĥ������vV���3�|O��\����J�I��wL�IZ�նĭ�˽ݘ��K}�������F�$���@2&&M�1TQ����!BYLRD�TR�	���kC�R�e@P�0Hđb�֫Xi�¸@b�9��Nb,��,Ѩ����c�w�0�����G�a�hxg�hW �|����<��{�&���i�g�vZFcQ���,���8��g��9马ţZ��4j��@ f�l�uV����l�Y������f`fd&�ne\lƖHLl��S�J�ffybn6V'+a��V�feY50�38�fH�79\ͬʳ3˭5�,�ˣ,(TU��i�m�o<�dѰ�x�Zs�z\j���R�:,�lgU�m�� Ґ���#*��9ͻ�e�F���B� ˚ՙa644RdJ�"R̻#���a�^c66v���l-GZ�녫�ӗ�Qʜ����\���E�Ղ�us=����g�#��oc����\�������6Wg��k-�SÖ=��rr7J�����5�.�t	��Ż[,=�H�]��O2v�R�ݰ4YvG���y�Y{����l���$s��Bev��Y�<�3UM�d�%�)�	6U)��uͲ��r*ĥ
�Mp�z����շ2�w;��R�O<Qf�-<sY�����ٛ��]�I��t���,�;H#�F��0&�m�+�vVj�j�v�j�%�ZU��������&�\70�H+3FY�\W�0�kh� ���L�P2#n��1�ӰEZ��˕h8D�m�!�;��6s�ͷ<�c;�� �5l�R$3�1���3WJ6t���	��sь�9R�f��g�d��w�����DCh;D^�M��>W;}@C����^hN�zXU?
��[���_g��sW�ޛ[R�x���ZR;����8��u��w��vj�P}�|'��\��𤘗�����$MKa���`�B��JA�����P�Kb�غ���H��b'3S��n��n�Po���p��	���)s2+�kQ�ʺ�Qn$�0:�{m�o}z`�,��3[7������A�"Z��w��G(�+�1?*��Ԯ���[|�8��җ�ZP&,y���KV�`y�(�7�p�r��T�@ڔCӉ�I�Bv��h�UQ��7q��٥��}�}�Z�Ns��°�SA��8c�`���P�Mw$�9�O��>���!i��tGe��3�k2l杺*�!���Phjo2Kx;4�%��ח=Z瞂�[�W���YEJZ.�A�둧d�y��XY\v0����^1][�ۡ�lգbKK����i.�l�B,�s��#5�$�I�>���}�~|��M��X���ܑ������0y���Xc:X�E.W"j5	$d�i��+��{�/n�~��q��{���ݟ�U�;R��U)���J�F>Ns��{u�n.�x�1t��[)\.�P^�(i���u0ɉ7x��`jݺ�S��n`.��A����"��Z�I9iIe$�ɇ��wR��%P33کwK+Fo��
���YR���K:�J�N�@�7�n�v2�30��C���n9(����Aw9�N�P���s�rR�GY2�.��8։�e�ZY�;�'��Vᯧ*�?2>嬵��:�7� �L�0&H��߭�NWq�GLK�]�5�gϱ��Z��nykPخP�nzWncFV?���uL:��d��ZLfkh6��,F�g'%�$���
t��uչ�Sk�$�����W]W��P�<�p����� ���V_���%)Ӂb��D]a��=��\�~a��z����(��s�uL��cv�e	��Z��t�0���A�٦��饁��n�=�M*�m��"�dT�8�0n���3�*����p�SPj�ݡ�Ry2f5���93�|��2���>�Mڷji��E)Hn�4��F����n��=6�g�4�GwQ���E�eQ(�4�n&i����"��׶ߞ�}W��*�7RU�5�bt��èx��y�˴����wn�qs�ʫ��U��SM*1CA#TU $@bꪻ<��N��'�uNW+��7����3;$����˻v1];��}?�۳K=���޸�bR2&��!ǻ����yiz�M����8��}ҽp�- [���c+�x��j�Ii8�t��V�{�o�[��|��7ͦ�J�R6��#�������M��e�r{���p��L��7�ھL�g��n�-Ǿ�x�"���q\�u��B�{��G*�;RU`��f;g����<��%%i]��J�>޽�a���@-�W`v�'��}��!�.L��KR[����h=���
������US-=�����q��ד؅N��"Iz7���T�pޟ�R�˧����l�&�9s"˰��ݶó�ޥKh�e���^a�%
�c.%�qe�3�Nyy������9z[����v�t&�%�z*�ح�ۣ�{�0u�O n�%p$���������f�|���?���攢fG�㬖�'v>���u+p�O@,]L����'%��r��l���h8;������z�t%P��W bJh5���6R�\�,��G�~\���+���w߯�`���x�Om�UUU�X�
�o���qډ������쥪���6��QG!�\Q��nWv�r\&�0)�b��d�k��>�O�.�z�����]�E�3��Кí��-��-���ʑ#qn���#�ӽ��1H�����V�͙
�u+�ƨ�)a�g9�\���������'���m;������O9������rMGy{u���]�K���\��}�_��|7��&��gr����P^�;F�'S2�����T��J�T�ТnG#y�}��`}�On0��i��������ׁ]���6:I�I��CD�<�Hf���������3zY_��+����.��!2#�m����?�~� ���pj�N�<�%1#�����v�(��T��{���5{��`}��n0�_��w���m��X��t�&Y�}�J�Ap�%i$��A.6��
���x�ۭv�xK1ۻ��9�(�ݎW2t��塢C�=������
S#�9��-e�˅ܵ8_k\̗e�U޵�]F���^�wag:�]>^����l95m�j�N���tu�tT�S�8'��J�wws �R� 尗�A?/E7�ûy�!��ȋ*�i����ӕ@^r�X�YS���w?E���U�En�iX스�wB���
�/;���QA��Ɉ����y��%ƛy���k�>��n0�t��?���r����������h��U�8'���n����5̀:qD�h�r�G��Aӷ�������yz< �G�pj�N^!@��d����zЈˌ�f��X�si��;�݁ڥ����s�(�3vy[+�^�R�%�di�S���ug��<�q�

i�*$���>�������-d�ӂޔ�r����{��?-�m1�<y-��;�����\��7�����{�޸X�gt���4�?;KT��@f��}�͔���R�m��]���,�!�˰�G/�E|f����{\T<��\�7�W�©.���ϿO}����^��}�����A)+m�m�n�M�GL���n7PZN���V�W ���7y]���*���������2ԗs}�_�?o���_��l>�g�`W�^Obq:�%��FI̮���}�W�{�[%=T:'][���������gt���Q<��8�X�r�͖J�1BO@r��p6qѼ�r�e]���]�����e]`l����[u��6�f�I�6�F8_9�����������w}�V�J^�iJ&b�"�Y)� ����R��T�@�*�.B[�� �ۀ�]���*f��!�����ܽ�R&�2���������-7m����� �W���W�T^�~�A���Iw�KL\�a�^��]ҭ���T��o�ObrB�`������U��@�j�ߵ��u�������^�����^���䗓�</Ʊ���a��	Y��B%V���t=Y3l���J��.|=�x��@��@�-��J� �	l�b�[Xg�a*�ӎs�o�-`l���\���D��gn��+F�'dy����*J�5�f�cDk�82�S�����)��qr�ή��owʞ�'S.�'r��� w��l?��d0y]�P\������ݣ6k0޷Z���y�E;AHU&fff>o��/O�pKަ�K�[��&�d�~�d����xZ�7&.I)!8�9R�w������`�^�0�^��2#��D�@������~a"A	IIbW���]+�`��@Zޥn`�)�:��).�q�B�;�� ����b��� HJ0�#���ߺꮭ��ý��+l;�fG�yd�0��	�~���5_}�ߺ���﹫�$�L�BL�y�>�֯�����3f��f��WI��g�r���g>��N�n�{2�fQ�ٸ�Z�#�&e�a�!�/y���� �P��e�w>�ַY�k]iz�&�eL"V.�c`IK
1s1���c ,�gbM�;bT�F�(�!�
JZJ4��	1G;v] ����HC�2��w}h�]�[ٳvY��lC��\:��U��J�wb��PUAWZ�-��m�keu\
�A�%`���{jꦒ�mUG]e��dz�j�v"bu��6�@2�.˳(	M����u�#s��nʮ�k(��nڢ�q#X����crq��H�e�6�um5/>�����a�%j���v� L	��<�!��[x���lun����3a�j�0���Z����D��s��E��W:r�n�t�1jec�V��Wv�Mm��[�Y��uk��qh�f��n�+�׌�.Dۢ�CƻPݜ'.{"��L5�qg2f{T�q�ڸ7d���d�u5e�nyRN�ccj��Ͷ� *����\��-�-�X�l����Vf�Z�a��(x��)��D��D{@T��Q:x
�Рl|Gb�{ץ��:4n�y��ar\P�2[[s�+�]��� ʄ�eR���7cU�lDK��or�q��	{m+�u�:uj��tLv���ܓD�H�(��	\.�_�f��>f�Go�~����ү�(�w#V슝P^�+�3R��g��gr���7����~��D�cɔ�i�����h-)�p��(�BW�<�D��+���c���\�9_Թ������`����l3��7w�,3��a"rd�3-[j����*8P��j�!(&T�iv�E��4%D-h�I��1�c�w#@;z8^��y�L�����{�u5������5
����>w��%�(�BW��ʜ9w+�5i�l��<T֭�,�yyj[R�w߷͈bK0��/� Fg�TŒ9	J�3!H���ʐ
@�#f�BlD�� D��"��A2'aڇq�:9������W����`{}���G}Ki4����:����3�<�R�<����z�7�[�����,���$��V����X�W��g����#�����mXG��޽0�^(�"RJI���P�vi2���fi����/�����P�+���*��BR<��<\E�6�y�]P�V���5+̼Ձ���8.�n�(�0���ҿ,
�����
AU܈Q[$V�>��g�3|���Kz�=�-�\���&u2�.fL�#�f�Ƕ�gϾׇ���0�@EC|��������M��[h7���b+�<���,wh�"�������Լ��z�/5+���;Ҷ���Ku�(��edRn�`uw};m��g�>n��,��j�eU��va�b���~���[w��l3绯��n�8�������q��V��&��qL�y�X1n�W����hݞN��}`�ʠ�w|�6��K�n���}�J�A��W��E�ҕ������~���=/$�5;Ӏ=P!�	z,�T��z��������X}�j��H�e��y���>�����~Uy�]���ʜ�fff�|��eÝ3h�4�[����WmN/e�Ƿe�kLZ1��ʥ�G9��OPt�Z{�t���P'#t�xbb�-u�xT��4�fҒڴL9ջB.�If��Kt�� �bPǛ=�L[��u\:H۵�0�@�v㫴�&��W&�{[����{Q����+m�#�;���0ʖf"JR*J>8�:���\ZӘ��ga��r&`��N��]�X�QA{��w������+�ʗ�rH�S����4�s�\��ڶ��k�h7����7_�@Z�Wa�%
%�`�i�)�`�Jf�%~fi��yת�{�`jݶ{�t��t�E�d���L��Ҋ�z��k�uN���Ù?8�S�8X���ҺWs�f�{q�����߻+wj��2���V����]ICy�jݶ�LIS���؈�YV�h����f#�aʌO3��-�E�z�����L��<TL����|�Y���N��
@��G[�zy��Z�N<��lvmö��/q�����ۻt�rW��&��m9=�#�����'<�l��z������H�:��5f��y�zբ�H�!�T�IJB*����+ ��%N�y~��o��l{�⃒e�Bbn�m�.na�{�1?*f���W`�*a�^����j�G)ĝ��v8���+pO����߷�5��Ꜿmq�N�[ww��«>��`{�����^�g��s�������<��JN[�����p>��w[��% )��'�(/:h��Yc�ܝv�
H���B�g��k�uNZP2%E;��Pp;�[�+0E+IX�j�	�k���8Z�J�3T��Y��\�=����h�WNSw=������j����T�����],��d��Ym��.Ƥ3�|��}�{r���������#�H���JJ�q��"�t����T�.W bJh/�n�F�4�<�NG�o�m�n�0�3wY3nk�t��g��)r��t�I.����վ[h>�z`i��{�Yr~�9�:���� ��*j�F1�C��m�����k���ʜt����T���$x�Ğ,f]D� ����_�J����+��w�-��;5+�ӝ@��h����u��r���y��]����Z|�"H�YŌ���Ă�
+"T�0�А��O�v	���=��o�ҿZ=�)n���w��0N�K�N�@f)�pԦ�Z���R��LRӻt:w�E������U�(���٦���]�b��r�t�$���UTUr������n������a���s��-����1Vr6�CGK��Q'�[���ʜ������!���\�;ǥ�BGV������n~�r�s�_���|37���w�-��<���`k�A}��
H�h��f9�K�:��v۾��U�?���������_���gT}���"
KW(V��G`w�Sw�=�߶}�Z�R�U��֌��h��ն50`@o*���mQV+[p��P,^8Cd����f����`Lڭ[h�:˷�J���vun����!��Z:k��z�vݺ�2m�.p�:
ZX2��Ԉ�-�8�@ƺwGH�ڣr�X�
���������ў�5Z��#�t�p"��������s�u[v��.�T�-y�ch��\-u;�O����9�}�y�~O�p�ܮ�5C(��y�h��ט`�ffW�u)Z�#0I4�e��7���)~����<���o�����;�fG�u�������|��1��>���r�~����3vY+���KIN��q8���W���0��eN6Y+�1%4ؓ�:���{���i�bK��|�����{�`wt��}ٻ����U�(�w%�JY%��{7V�U�Ug�V?����4���WP�nݗ����l���f_���N�޻K*s{�� ��t��n���+,�����(�UB��Xd���vp@!*:WX�4�MQ��16��h�;��.�갡`�-Ǟt�+ޞ��S\�"6S�f��ʘ��-�=�׶��<� �P��n�Oa����h���"���픯�33O�矗������wޕ���w�V��H��h��0],�ñK%p$�����p7�AJN[rݸȜ�g*���u`�J�A߽7q�Ww]�wY�֝Ȗ1�+�����m����:���
y�5A�mz���Ky+��P�,����p頇��ww��:YB�<"�k�V
����gi���ΞW n�*pX��`%��a�s|3]5K��������I�������[��Z��5)eN6R���G��A���Ұn���zV�03�*���W`�9�㔎��Cŷ/)G�ܙ���r�9_������~��:�n���nV�/6�% ���M[%�~����IVASu)�A4H!�SGJ�j@�qb��f~z��,���*�u�L�$yr"�"��0Lc��О�:*���fe��uB���en	�(�/:R�t<�Z��r�e%-AȮ��ە�j�eN6y\(����$�~A,E�M���͏R�v'J��Wf�6&��j"�$��!aG��њִ�F1�Cd"ѥ\X3f��p��$��Q�ۼ���0�aa���yof�`N��Y;٥L��P�Q6����[�A���:�MI�䅗9q.���F�宁/4�NH��#FD��)FIM	���`Q���Z�+$�CJ�X@���")�)JJb"
&6$,��e�N,R2���x��D�K{DJЙ�jbJ � ��`�XjU���H�H�9	I@b� UJ8�!�ʊZCP-�Ġ���&,�%��0�(��)00���bįP��G T�K	)�������4��WkM�m�3�Q�@[�hJh�2�σ6ٮ���@/RL��cC�e�Ͷʳ3/,�̄̄�*�}*�L�2��V�i��fu1��s6�3��R34�2��*�s)�30�f�̺]��3��h��avKړ\�<�m�ؙy�q�dg��k�̦C
���뫥Ê�մRp<;�[�3HF�s�6c`r* 	�qsi+G��-,���*�s�Wl�5͜�f{6����3�U�Z1�t!k�hBbU�v�M���.na�N�nڃ;[�����X��y
�(VNDNy|u�b[����9�3]�Dݶn��&^'B� b�-��^e �/3*ܞ�[nRlm������e2ӹ؎:<8�/ON�΂�� �u��<敭d�yy;�ܬ�d56xٗv�2�u*�^��Pܛm��*��<�ɀ{9q'���s�[t̚�x
�݀;l�Y��Mӳ��pD��kv���9�$��؛0�00T���ku��cv��
1���������Me骞��oI�vÜΙ����˭��m��[���y�%���+��3�؁f��&z��r�,�n��mN�n�dI�J B8�q56l�v6�0S`v�l:�*��c7[�ą�:[�꒸M�cl�W:�1R�T"�M��e��#� ��|���辊)�l��	=T��C�<����y�9�ߟo��<�=>�L��-��+�>�qޭ�a��ܬ�]��m����6q3-^Z��n�`}�ڬ:����TI	�B������k��aDnَ̥]����Y f�Uۼ�ù;�)x�&a����jx��Ct�AK�l��d&d*C�g�n��(��C}`�v��o�=�ME-;����;�M+��|�;�ޕ��C/T�K%p2�M* NYq	ZN�.��n`��՟˜�[ҏ[����Nn�C���.���܉��5�J�/zy=��Ҋ��37�r[�B����dA�e]n��l�U+2�m������%�.څ���F�Ƹ�`nvp�:�e�[t��P��Pu��\EM��[R�v�V��6���a9������.,�CU�/\�q��!��������Ra��J'+�\��U�w��Ϻ��SL�Ge�J���a���*�U�<�%�)-�����&�l�sF�01#�{�>�5?�P�>��n�MA����;�:��>v��<��˭�SM�N �Ӕ�*u�վ[h3ww0�ym������m-%:���FۺNL�͔�>�|�33����@.�{�`�vٕ��*Z�p�<�*f{�u@,�nW�fw��?�û���5<;��}�Z�5��Z#9����!�`��u���������@Z�J�Oʠ�Mȇ��y��26�W�jݶܪ�X�����#��ol��ycnR��3̸�	w{��Ҋ�e��3������o3\����|aV0 �뗟o�MF8����+0�\b�Vࡂ�`av�n �ԻlV֑7k���^��xv�\om���e���.FFV.u��s�w�bx�4[(�"٭���z?���mr��Vg[��{�`	t*p��~���7����7x���8E�s2#�ڽ���~�yU�����}����%FB)����CT�8�Ը�TL�����߱��y*p��W`k�(��tȔA2�c�\�U`f�������1�ʠ���3}(#��g�����uG���~2���j�ںt�6��f�0�J��LI7Q�kM51�ͥ����q�%�e�^w��R{>���C�CM��|�7�٨\����.�,n�)*!��0<��vn���>�����0��J3.��������@~���[�J����k黟ܮW�������|�`(�M����J(3Oڈ���N�#�RExWOm����V���f��c�O��@f�	���R
�n�ղQh3wۘ�M�a��n��ݖ��Z��M�S<�D�������2���%)8�EM���omz�������$��60�}�Q��<�^���V������i�sm��k��+�D�
8F����wצ�쭴�W����_��@��uq؋z��(xk�.��Ji��)\.�T�e'��j�h6Gd�%lv����f�0;yM���8��H�3zYS��3�)����U������������~7�0>��>�M�g{�'�G �� ��A�vn����%R1T�8���4�s�tnEt�JV������P��S��9��PjI����X�W�:�Y����,҂BY]Mh��u�h"k �RާI+�1�(�-F�c4=��@�����I�-�{���j�Eٳ��}���윁��&��,�����P�����Rʜ-)��}�^Z�d�;�]\q�a�������j�=�_������]W`~Tv�&�SЕ\�2j� �$d�~߸���m����¦����*�Q�96�:�d��bfw:�l���l5���ذ�%�n(�CK���,����z��'���A��1��aB����%�n0�l�jV�61Rږ6�cLdׄ�1m�
b��������s�}ʕU�o���a�/W�E��"ƦRUu���W}���u�?ys���ɵ)bs'lu����4LD��A.�w��7��@fw+k�����,�E�N���w��W&[t��)M7)6�߿O߱�����}7�������h�?n���p���J冻�K*p�ܮ ��4��V��-�Em6����	����=�^����g{JR�|�4ɹ�16E��E��C`f�T�ܮ���ʜ���3�k	�ĝ��v$����n�9����hZ�#)4�F&��A�Ԧ�n*mgz�u�~�+ �vV�;����p�.�_7�*�,�R8R�a���HN[f�䕞x_�5!��L�V�2����I`WX�Dq�3�hhlkgj��5;�Ρ�nMc��`��w�Gy�c���m�b�����)�/�Y�V���,}������NW f�Tዹ]�h�r������u,�en�ۻ,��wu{o�*/u~���1�Ȗ
Վ�U6��O��O+�}��;��^��{�����i��bJ�ӎ��������`��M@-�d� ����C��g�x�,��t� >���	.�*C����"+�:Ul1����A��$�bԟ@��EiO+������r�YxQO���飷F�k���e�BZ%��V��Щ�;����n�3Ǐl���N�V\��3 ���پϛ��Y���WZ� �~U����;G��i��4�.�V۳ې'J��V���S�X\������{��%��y*j{U2�������n�4�
�w�p>��u`�Y�7 �CP�%8��T���t��j�(CEYe����}�{m��J�N�Aܾ~hN8E�ӻU#L���wX�u�N���� 3_�@g.�n�SPWS+q��2a�K��J��l>�ws >������P�י���~m��h����Tݻ]sy�5�Uy�?~櫿|����T%��bĄ� �Z��S�\�Qg�o�a�����u$�#�q�TS�DL8�����]
�3u+�����OdJJ�1,��݃��k����GN�U�����2ۆXA�J[�6�j�{����-�_�@bԭ�Κ&Y�⪫�\�pWv�캎���VvMdׇ��U�pĕ5 �u"�3T*s�y�R1Dd��R�X�Y�}�l���Gz���ÿ�W�A�����yji�H�T��Ș��Ų��jS@f��䩨^�*=%)#ȝ�U�����m�_��[~~���U�T� �	et�6Y�dVI��j�,1n�lK�	qQ�1ia5e�� � �����fA>rhK׭�]�7NQތ��$���c�I�4n&�9��ssiӮ�c��u\ڸ����N�w���m��8�AE�6��	N��}��=�Ϻ�Ť�RQr\�i�r+A����aS�v3�0�cmy'F��2�nIN��*)Ȕ߼n��g�`����M^��*k�(S�Ti4��B�q:G)qԒ���{v����צ f�Tᛲ����d�.��O5P�M$��@fF��;��8Z\���BU�}�U*<Jbc̍0� ���`}���a��+m���07��U��A\R0wx�
���J��Q@fF��;���ݮ�[��,��MSe�`Z{m����=��͹��u�`w1�M�N�M�6�:M8P���h�ݔn�+��ID8��2�D��7�kc~g W�� .�/�Y�Ug��6_�|0,r�M!2H�ִ��fA��P�`X��ܰ�b��%�&�r7�\G�LI`�u���C7�ʋ0��4h�(W0��X�	��bF ca����G�ј�K��c��a��@%	A�w�6��`��
�IÂJX4Ң���e��8� �!&Ld2��!~ܴ��%IJ��N\;C�P�JJ�"����ZJ:���)�
���
t'A� v2�v��j�)h��8`�!�;�0��o3-��.�0
�@m�<W6ȅNx�E�T*��$���W�@h%�v�ĵR���'U�PG&5����F`ۦ�joF�FjN����n^΅�B�Aڭ��fz�-0F�C٭��- 
V	8έ��2ְΛ͖QJN^k�4��]ۘ�	U�0�妲��j��1�ڷ3	-�+��m��x���T���q��;�v���k��m�2�F����I�\C���NK��	��ݪ;fc0�1�V�P�R���j�-ֆk�d�j�j^h��u��Ks�y��(T�l^�tm��[���7V�:Ӎŵ�^�t����N��g�L�dm�L��؝�C=L��J�.�����[kp��e�X��Z��Y�ލYv��� ���x���j��
hOD�z�]jܫ��ۈ5�v�&�v��J�b�ݦCAƤk�* Rb��#�Ki�m-i�r+V��#��{�;O�ֶ�s�?I��I�O���|�xtl��s%6�T��G*ӹV�Z�wv`jS@f�p�r�7!�CT˽�vE�t97a��ʜ-o+��M�ٺ��U%[�k�� C�8��9%��r���Q@.ަV��ܢ��gBq�w���xg�����*�̄�X�+mov���=����X;�&�����Xxee' �c'���T�Ň��-u`�V$�*y����W`wt��0�R;ÌDM�E���9�#�_<HV�����ue��^f^e��N���ճ��5�K�7���p;����=G�_��Re�%�dV�����u�����*8!��7���_y��X�[���֦k��oeی�]��Ҋf�%p��(�W}�Ɯ�!B���]��>�^��V�Z�[�����g�����<qU`���%�ջl-�$n7IA��瓳���&���j�<�优���;�Q@nl�Wn�M,^��gRa���Pri��f�R�D��M}���]=���}� �}+m���Od)V�dh�QL��IE��H���@-�Wa���q�;.�H�U`w��������s�ڮqW)�ݗ�j��������IR�;���XU��f��g�U��w��Ꮅm��9Kw����4���������V��	+a����r�kD�Ni�4b[�H6͉^.��E˹&@n�W v�*�v�I��5��^e��^,�e��bb�D�`s�@fG�w��T�����dr;�ڤ�\q�{}�Y���>f��������^��T�	?q-0�RG�����<�������o�0�UIj�����^��c>����RQwwʉ�P�R�uΩùr��ߚ����"f�a͌*`�[V�d�j�X�д#��T�L`�u�����if�ZcZ�b���*���M �G�HD��p-nq��v��D��v`U ���/�Q�
[�����
�EC��#��n�\����VX�"��"�����s�twy��i�k�k2�3�ݺ�?�ʮS���P��XdZ6:�D+��h��FƩPܦ���"~�_�u��^�a����i�.ݐN�ģ9����a��k��~|?_}��J(Z�[�:N�����\�H�ԓ��j�Tᛲ��n�M@nvV�3��*�Ԩ)c�	)tQl=���`'�*�̎�ޔPjmC)��yy{��"఻t�S�r�m`�M��޽������"�I\N&�ZiX���q��3��r�1R��u"&1�0-ֹn�f��R%m�w���W`s�QA�����S.�=�l��{p\
X��Bfb	%�a� �`"�&)�`��")Yi
e��F+' f�&Yd���C%��" ��R@��h� ����f��I� BT%�!a�Rb$&Bi���i
���/~x|�)����3�5"PqR��si,2]�*4�e�ň�=�|;U�6̝�n��8v�6N�+�e��Jj��䓜�󜜚=����\��+��n�~[�zYS��v:N���E�os���M�')ܦ�V�}{�=ݚX}ؓ�k�3334�o�g�y�,��ˈ��O��P��W��ʜ/9+��DymJmݻ"hwP�+a��L ��h�ԭ�}�H��M.C8DM�<�rӁx�m���Y�$Ȕ��{�2�`b�V��f,x��ŭ�J?%��+���	�s���`�����<����!��"`��ĕ��r�K���e�wkS5�JM�Wx�Eu&`w�o�z�U�LL?Q(� ��\
�,G0�����t��@rx1���3���|ͤ�Ϲ�s�Tv�+�W����r���b�I`f��ý�eO���fw���v���/�A#�EU��K�\�`�M��J�7T��ϻ7Vw����-��Q�����w]�d�ء�Я!�J+��������J~���Om�>�M�a��V�;���OeAV$�WD2��pITFju|���.Q@f����S���V�\��&�Kd�"QX}ٺ�����v{q��|����S���1,���
�]��Ϲ��~o��I��F ~r�B��fP8DP�*�F"��HU.*ˊ�� 9�u���]y���:�߭l�r*N�]�lr	Z?q~�o�����36Y+�;yM�N)�g�-�.�4�`yw�m������H�E��c���6v�zY�mbJ�,��1JW�d�&c�c���d<s�\��];;�4�L<P�xV�b�T�y_��fj��}�~,?Q�?G����&��e+��M�;�ި����}�A���^JT�(����TN+A��7q����y���(��jRާ5��3�x���i�����3T��Y%p�SA���<|�h�e͑*�@�m;��3 dD�\M�VS0\*�o��.��l�ZDM���иz�=�D��\т��M�¡,��		|hu�k��m�G'El�G�c�on�Ft��p2�Zw$l<���lC{$�$cjJ�*�\�Z^�}���L��ڸ�*B"�3_}� �Li�*x���n�k-�c�ù3���#�gw2N�<�lrz�J�g'��{�B�:�8-f�7�h4�g$�h����P����(�>����7�MV��AKj	
]+;g��'�uN�y=��Ҋ��B���b��u������>���zi`{��s�7��S�"�#J:��V�q���@_o+�9��S��9�P�R�yh&X��>]���T���篅]�f�ιfqlM�Н:q�)9���~��7]n��}z`W��҉��ӓ���V�)I3Q�g��g}Mh,��x�c�m�Q���ڶ��{�Ꝣ�F{W)����Q���$��N��7V��������I^w��^��0�#de��R)MȺ��?n0�۷V�q���ʠ�N2�$\��=�A`s�:�]<+p��Q@^)�pf��mJ�ܷQ�;�F��Ϸצ��Q@vl�ԩ�9��'�����..^�d.�>�����y�8^��b+��5�D��i8;�0�}�ی�'�<35���3k�5H��2�AHƛH2�6���׷Xw���`{Ҷ��ޯ&k����w�\�����3*�J�mx0-s��ߞ��h��+�5:U}��Ã_�C�C�K�-P���gvx��W>��*��B�R��І�O��W�}�|���~��;�^�g��odE�e�� ��,��se+�ĥ�Kr���4�J��������s �}�Vw}u����^��,7���ҥ�Tb�c�wM�޺���*�W�+�#Jr�1BG2��
V�AP��9�����(�l�p%����i"b���8v�Y�b����kZ�E�`x���-ùO���Ҩ��v��ý���%%I��byv�0�Щ��R�v8T�iO'�}�����<͕�D���H�?w���a�_���mW�6x&� s�w��6:f,���P0�a��`A��c�i6��N�%���#&��y��l�f���h,C����@��0C��-�ZM� D�4��ew�'�N,c���⋰0I1}����#g�J=,�7�n�'���9y�Ib^��r�Aٛ�nql#�����اWZ�.���Ͷ��̫3 �eY��̩��Қ�g�����9�������6WkfW3�W�Bm�fU�-n��������3��U�;5��{u�����#\N�]68��Ҷ���ڧ+m�0.��Y�m�%Ɍ���[V ڼe˲�Su�C{ h��Қ�@���6��Ւ�gɇ\H���hQ�`�ll�˙�k�L[l��n]ίmي��i����Np�9]vR��t�j�v^��s͵c۷	��Ӻ��N�֜�^�2;�룃bC���ڪ�&n4I�綆tܼ6��+v��A�0�	*��Ga�[��n'���͇Ǩ ����\.�sF�z���j,�5��S�E�b�j.8r��n�� �#G+��]6- ͘&�fb���lJJ�m�PCb��2�h�\��M�PƊ�tm�D��n"f݊�x�-��Fޝ����;�����#c<W�t�ۦhMb��֧ ��nwVm�v3d���&���m�7D��:�V�jC�b� OI!�4�u�1����2����`�+���^�,��4��Ḵ�;#�ͫlJr�T���Z�M��[C��q�[��c{���Tݛg5Y�ݣ7���ovog��
�G�O�.�Ȏ���1E�:<�A8<\E!P���~O_� o����aX���h������[(V�ot*p�ԮþU��t�Q�)ܩ-�n�j�<���]�iuf3Q�-]$��8�����?�}���{q����FѾ=������|<u"t�ɛQ��&s�������-���W ��5ke��7{�q<���L�4T4�A��]����ҞO`}�M,;Zj�KS5��0�`,��Е@f�J,S�P�R�5!���%UMT�}KP�D� ��Tᙫ�<����|�!,C1:�rM�J�T��9Ԕ;��1%A��&poK':��(�;Zۧ-�5�m�{%����"wS�?r�������0�֓g�����k���Qi����E�����K,�<�,<�P�!�Çn��Ԋ ���'9�r��W9U����џo�����y��Zln^��4�?��T??.A��d��g��Z�m���H�
��䐌���߱�˧��}�ۯ}�j�9P����ClM��9����e���=���-�M@Z�d� ��T��r��3.�dD�CT]�����;��W�R�� �l��W���u$Ucb�ն����� Ԕ��R��(��� r��Ĳ y��z�m�����������W�媝F�Ii�)�KA����^@�"JmH�ڪM�>0�������h$�<F]���P�������P�𤁢�b��9e�KM��r��5�~4�#��[1m��'9�lkO�#��6"4mR��erѨ�A�����j�l\n�9�����qKe�J4K
�M�Q�Қ<̓�''9;3,w(^��^bU����ؑ)_C{�K<��xޭ�a��oq�y0ڕ�n탒��`}��H�1t��I+�1Е@�d�B���-��#�0��7ݛ��{饁�}�xVѭ�$��J*��+���J�;�������3�YS�'�8)I���ۄQf��v�\��ثh1�4�f�w^t;Q��9��~���������)�l�phv��4(W���V�����6j�E8
IRD�S����n� ޭ�a��n��s�@�{�X}�����Is�s�Ϊ��v}�A(�$lQ_��J˰5�ʠ1F�_����%ib �*^j���bJ˧޸](�/vR{ �we�i�N�-���sx]6f����J=N������eN�W`�<CF�)�;n[�(�V��n�W9���g�:u�m`{y���Q���AA� Fg{�u�}��n�ia����`�U� �4�H'n�@�pj6�nT��� �we���j�}9y�f��]�����7�i�&]�C��J�g�7s�9�UTGW��;���\��W���f�Խ������r7k5�U~���\�ϵ���k���� �y9\�W!�~�,��߱���ӧ��MKLıP~�����r���ާ��UK������~�g���e�r�,�;�{hS��2	q
Fۉ.Un,ՙ���4H��Uf~�](�7cD��f��L�My��<G��Б�
"9z�Mq�KK��`wt����U}�H�1)eH���mU5Ox�0`|�u��U3|��s�\���8.�Wa��D���-��ȇ�%��_M�`{۲��{=�ë���߷u�!#�wR�q6��0.��g����w��j�Ͼ�\�@�ȁ����421��d�NK��y���V6S"��N95��b��z��cbTЎ,l�j���ؔ�UZ��
̖���]�a��5�2K�@��8��s9ڷ��
������j:�̫q�lˎR�vƠ�:�Q�!�4[�r�3hfevy�y��$����۾�_��5�ʄ�K�C��U��wۘe�!�}��#��i�[��d�!8�>)8�Kwwk@�vV�0>ջlͯh��9�7�j�tى�J����R��9��"Y����l3��m`bJ���S��lP�44̻Q<�5D;�-�m`'�uN��[�I]Xo|?CB����`���n���v��T��'�l�t�0�4�-5-2�@_)�p��P������9T�=����{���A��˘�8*YY���u`&��F��"���+vI�[j�® �`~����p�ӕ@go+�\s�	�Xy�yߌ}��|��g�b8Ŕ�t�\�BԀu����k�P����`��-n�l�4�´�ǧJ�Ov4.	񸹄�D�I93!5
�\��8���N)IH$�H�0����`{�K=�ی:���7�n֪t��%*:������:��ԭ�$��]����kz�);��n1�v{���5�J�/#NW�Ҋ���)��x����i�%���]�7y[X�P���GC��CۖIv6Ҕ���}�|ֽ��[q�1,f��y���K����S�~|��勵~~�����=���q$<Yu��
��0�՚.���ӽ�t�v��P�y\�9~��f��/[X2I��Cd�q�k��F��}{�˪�*����-����SP�S+p3�*r��*[9`�Z�Sf`]��ڷq��).�߭���f�ɺk\�Ii1]�&&j�
��S@nl�ISP.�[�'	1^L�Sq������
&�/*�y��/OV��0R�Ī"H�*}��wuwu�����+�B�V£�;�� �R�)8&� �C'$��R�%
���o�0.9T-�7�@��Ľ��b^ɛ������i�7z,}��8gl�q���Ө�w%ʑ����n:��v}��P���������s �i�w������X��r�,�X���4��+�ĕ5����e/E��U4~R��\N�6��Wa��=���*�5��m����9Z�K�X��%*���:�׾���>[���w��������w�> �u���m��(�S�����|DN��Om��vxV�n��g����<��DAQ31NCD����E��S�p���p��v�v��H�ə��8,s0>�m8no+������.�z���v�M$MN��;�K5A{���3�Q@k�徫<Q?�K+8�@-2H�*]v�+�Ѭֳ-f�����]l�[i�3����[i�#����L��s��W���S�Nu̺h�578����-�J:r�������ˊ�B�cp��̂�Gi�.M���N�M��SGa7�м�b�٠��w-�6�(]�Y�4����Hr{����v����Ȕ���!�if�o�z[��Y�c��5�����^h�f�c6	���y���_�����Aﻷ���֙N��[NQd@#�n˙v�V���_����[�����y]���ʜ�Dt��uxfKq`�`uwu���n0=����`W���N�C$�w:n��;5R�jS@ol���~U��T����햘�;������w�U�k�QA���g�u{�!<1�a投�ʑ�a���f���Q'%&;�"�%v�p�e� G�3���f�2N��[�ڔ�wع�h�Fo����^!�y��=�|{(�%�\>�l$�0�;�И���P�H���C�;xAD��VF.f��BP�SM"b���љf��bYfFFf�dK�L�&�4i2��2���,�,����
�ͫ�R4�����NdVZ<4��<���9�;�!ݱl$H���4894�E�i8�;JZ6=�Dۡ�/Bh2YJZ%�!�E�}Y��[ݻzѻ���5ў�NI�i�@��ֻB� IRV�*DR1�+��WT��A�uAZ:���-d�T+kkF��U�h"s��:,��Uݲ(7-ʜZA����3S��8�9i�m�W��we����G���[�4m�.A��В��9ɸ7'8��KD�]N�2f�qȗ1��A fv�s�;��yݰ���v�g�nh���c�N=�J�X�,����R�%.���� ;��d7ڤ�!hl�B`qh%���9�WHh^�ǲd,V�s;��`QL�[5ٴTl�,L)�M�2@E.f�X�:fPƣ*]i+@B�J:�C0� �6�h]�@��aHmkp*Z|��돯����<ͺ�kyo �x򀆍)�����ҜAC��+� �VG���I��}��l�&+,Ƹp,��[��p�QC)�ڰ;33R�̱�U)��@�N�K��f��;ds;'Ln�H��K�{[��{��{��O��	l�q��]�Z-jg�ぼ�T��;��8�9\	��oQ%'i]�j)������n��o)�3zYS����S//sUWp�T�0]�ڔ�vP���~U{��¾�^�!ܱܢ�JSv�����5)�5l�p�J���К%� �..)�@V��>練'l�UqH� fK10�.�D�fcEd���Ooyz�Ԧ���V�ot&� �z��V��4&`V�%E��%����\���Ҋ Y�����|��{�!��Ĵ��<�=���J��`���\oJ(�T���?���5��DR�v۶8ݠ�o����<�;��:M.��7qwD�D�]���T��v �Ҩ=���>F�\�a�xiv����b���
�U/5��^��̺g�*i�V�r�*0Mt%@RTs=�=��z��u{m������)�JS9*F��`���\l��֘����Ҋ ��J�Oʠ;Wa�jS1Ҝ�5Wr����b��0���X��{�w^��US]�l�k-ݫn�:˪�~�_��׾oߺע�f;@�e  ��	T1T�-@��%-	JR�P�JR%	D�"�0�!P�1X\�B��U��3���`���g�j�ԥG(�Z�n�:Wa�w0�[��|�q����õ��l��L�c�؞`�YP��n�8�bLQ)P�P�%���۬5it�w�}Kƀ%Щ��O+�d�0IDM��t��%=ל�.�2P͎W g:Uؒ�>���Z��92e�N�`}�M,��+��Rʜ/w�ͬ�rihy�%夙�/uR�ޔP��V�Ҷg���:r%19���� ���`b��0������ϫ�>}󤐔i!�M��2 �n�k��30GTU�]��.�r�O�َ�*E8`�)�@ґ�h�̹'�GQ;W_�܌Jn�V&�keblL��N��v��q�=3,���� %Z%���ͭ��3���u��q�3-�����������;�ԊT��ܫ$�V�;�]n O���G�*l��(�Q���CR���`��~����	oR�](��Dt��z���j��uef妔���c��l�P��\�}J(}N��ټ�S�d���'M�Z}�n`�[��;�]n ;�l���Z���)�ܘ���5a����U��gs|��@b���i���r�.Ԍj�HҰ:��w}�,�óy]���A}��8�3��L⒲���X
r0W�!"��꓎�g<GƣQ�I�a�^o5r�ޔP��V�a�Lq���Kպ9T9�iaM��4��V�2]��h\lh[P�Z�xU�[B�m
� ѻ`�ۘJ�M�
���-+�D��.ʼ�)��0�2�]�9�Zj�{o����'Ԣ����{�l��Rާ����Ey.�M�(ǘ��v�r#��ۯ؀���`g{������5Pm�.N+mH(�r� �t���W ��E�immE&�:3*+M击�[h=�|��턞��7�>wS{�rQ搈%���n�	Z����?Us�U�}�WÑ��c�f�`NZ�E5��X���Ď�A2��/ �IU�bJh-.	��-��;���n��T�ThK���D�%6�W���uo�f��V�����ou7F�)�;w��X�,���������}l�t�e8nw+�>�M,=�Rݨ��fd�je��S@_l�q�w������m�6�v'j�7QT���ی=��Vw��q�}�[�*��﷟��ˎ:���~,��9Uy�R��J�	*j��q�PF{�'�C��y�&�}�1r���W$���^�q�nB,�LÆ�47+̳��� j�U`n���ݞW���8z������:�]��;�J�p��W`b�E Z��prL��yiyb�j۫N��3훸���[kܾ�TUs����4-�����[h�oCh[$�S#���v'���V{��q�}�[h>�wswƸ�j�ۑ�%8�gW}l?^b)~��t�1��D��PR�2�aX57�L[�~}�����y���G
�I���^Z.����|��o�pKw�ˍ�<��氒��C� �O���W����k��魴W����PL�\�0r�������;�5 _?u@��P^6�<A//6�UNK̐�v��S�ݰ���ޚog�^���T��ʱ��H���W9�f|�P�YS��O+��nǉ�gi�b�{F)����J�T��fMpa�;�k�Xrv�]�ԋ��L�x�驻i�vqz:4t�g��7ln6LFo!�M�:sεn�GF݋jwn �v�t�g����q�&�mves��lH�\��Jl˵�\oj�_W+���۫�[OkRl�f(�dM<�>��˲�F�N��D�5"8�Y]�D�5n#)s�����X��S��aS������.�Lѻ���,�K�v�g4^H���,wJ��-��P�<P�5�G��i7��s�1�ӫk0>��Հ^��/�z�/9+�I���,<�<ː;�1N-�Nf����[�k�m�;�k5����R�3 �ޕ�ḥ+�ĥ|��a�;<pKKŗj�v�v��s ˻t%Y
NJL�űa �����k���*>y����Γ�����foM���)y�;��O�|�Cx�S�F�M��rs�ی;<��H��+t��lїV���%� g1!�˥��vu��Wk��b9����L�<��s���;sKzk�ᰮ��ƫ��g�"b��^��<P�-�೧ی�wƶ�ۖ[-Hӌ��������y�]���5~o��.oxy�{����{i-�����ԭö�@}���
����6FZMZ��)����1G
�����.���%:�suu�Y����X�C�*$ͳp��7mƃ���Q�/CP��c�/�k�@{�~��{s{�;}FN�[�eO.�����*VEUD�ģ1{�P�ӥ��}���?�w�V�T����#�^ jt�~i��c����/:R��SP}�m�=CG�MGv�eZu��{r��*p��n�ݞ(o%��Z�f�x��]��>Ǐz�1������z~�g�wZN�%�#�$NB�X__������1��ک�v��M��a�P���d�J�Ͽ�����s �_��w�K�h۸�I2�
��:8x8�<��vY���.�~!�Ҋsg��c�*������h~Zf��j�jxg�Δ���5χm�>��֌�t4[$�Q�r�;$`^��o��מ������C��>��bI�`޸�ە�G�(9��K9�.u��z�p
rm�u�HHT��:$�
1A�ن�'&)B��D�oj9Jc�Pf\�yX3�@��Fa�e��8�f�'z���Y���;�\մ�!������3jq4�R�w=#:,���V6 �1��D&	 ����`����{B6솝���&yl���]
p�;��޴eV�*:�)l��1�)�6$� �Ǒh���4Zx�Z��i���q���M�;:�Е�F��OUh��#�5�+����1i`kh�<�R�)UV�<sY�`ٶ���VffU����'9�mfgas2��KN�7k9����fb:�feY�����̫;�����&e��ݓZ���;Zi7S5�n�s�,�j���g�-m��v�6MY����=�;J���|�9mB	5�a�ݬf�3�v��v��D�JU#��u��̼S�T�ݍ����3�[��g$�M�zN�`$�v��cgk:ùnfNu�oK��e�	��r���%S���n4��	�8���:�筌��.z���N�(8�ݜr*@oI��l���E��z:��a�H�,�c�<(l�b�QJ����{k�Au����{\z�1�g�gn$2��x�\S��F-zT�̶�ù�D�����G&�E�n�Z���O5�\��!�h��9˱C1�C�h�nyJ�8�jZb�P�ˌg���������-ӳX�p��k����Ii��+7���7h�Z2V�ct#��:S���h�r��;U�z¼ud즮;C�T
�Y�����ZoV�[�:[D�;��]/�v͓�� �p�Gd�m����XGl͓u�L,ru�)ݺ���<5�u�G��n�x6��L����1��5�n�DM����C�N")�� �O@8�c��/W+���a���|X������q��e��ht�a�����K>����M,=�V蔊RɌ+2�`��ޖ��wZm���+�f7
T(5bpN�:B�	�۸��V}��h���}PP�\i�,y�J֩-��i\�{������u�����mI��F���^2�	<���i`y}��l3}��Ewƺ�#�ݫ�CwD�+�Ku8_t�S�[��t%PnsDGjIЯ/2շ��k0��=���o�Ϸ����BO<���^8��)gYy� �U�1��Q,����mY仇=��0�a�L�p�j eX�-&!�jW@�`��h(��.z�q��3�?�]��r�ڌԡ��;#ֳ��F�F���*``hE��k��Wj����ёW��9#�$���9�W9I{��V}�*t�nX�X�7t��{׸�ԼF1�$��TAҭh]�E�[q1�`։~}���K��8^��S�R�xt�4M��o��=����� ]�m�l�&3�L>`�eꀷ�uN�t���uO�l���:?T����*I�#,/���3��/vR�ޔP_|��DC<�D�;E��ᜥ�J�Pܪ�u���7^D���v���R���M�`�J(|������ļ<�YW�Ve�<���4�*��Ӷܤ�QƠbV�f1Rʺ�`-�]��D�K���e��<P	o+�m�qA1�{z~��hw��V�3�Mı)v-��,;��q���s�ѳ&�nS;��!���݇۰�8NSY��t���GL[h�[�ח����bێ^slV�VN��-�����1����_5��3:R�|�!�O��W����-R��ML��k�3ݞ�a�vV���,+;���"�wk�L��P	l��I�}��p��~�7��č���#�iUҋ0��K�Uo��@^l�po!�S-$�QP�m+m[��,�k�H�R�)2�t��:��4�Ֆmڮv���ĹݞW�9=o0ɡ<90�_;��Yf��
L19[-+�%E�Ř�嶃����;�M?W9�<�{����ht��v�ʷ*'��v~���Ni 	�9�~h��j����p溜��B�JV71Rf<Q,��G'�-ֺ��3;��uN����N��wM�r8�VW�v�b��v}ٻ�>��fQ�j�ӷ&G�#q���l���|�'J��L@%B�*�,as0<!`�T����߾��;��Vu���ݪK�C$av�I*?��;��+�tԔ�[�f:�7��]�ܕ5���/#y�-�CE��u]�]L%�f�u���Vw޺�7{7q��F�Q�ˍҴ:�s�ך���^g~g�����j�Ԯ��ʚ�Q��w�yg�{a��^�w�}9T�J��nU���=>��7����Y.��G��n��w���	��6Wi�� �g&��)Ԧ���_{����۫ �u�������c�\��m$��(����I�$T��0;��V�7u@[�P���6oC�i�x�*j��)����-BO^o�fgszz��������<�ߞ��)�r%WMe`wB��ԭ�u*j3e�8��3�C��+%�)�J�g����u�l3^���>"�2KI� �IR���Q��bU�	F�I�Y~o�ZI����$m�B�(슈q�T�������L��c啋nq��]�v")5�a�t�=6@:l�`���n.Q�X޸����[��WM6	]��ݮ��-��[�����bv�f̘�ɭ0m��c��vӽ��kfV����
)ਯ�5������-{H0O3%�Ӷ��u�l��MD2�&0Ս5
T�e!"�*j*J�*F,�w���w������7��ѵ )n�ʴ��%������4ʌ2��m�>}g�ԷӺ�/�+�3a�T�.�C�C<�]�5l3݆(I�[)\(d��z���:*n��Q;.*B��a��oq\��͖T�o��N.�O�����"�ڪ^H���>�^z�z�/����ٻ��{�5�'$��-*J���;�]Xb0��p���@��c`�r�M�hԮ�0�ϟ}�������wv�ý�o6�!�<|����h3qFh:����
���p��<md��mp�i.�����q�5wU�s�x�k'>cK���ӹaH��&�I9��NE��+sqf�b�DURSD��ƚ��u��-����~�����e�Z(����is�*-J�9Ҩݞ(�zl7���#c*:��̡Zy����X�(�-�_����+��Q�L�M1��A���<{���ʜ<�+�jݶ{���z�!7��[�q�x�}��ogt�uY�r�JE��B�1V�L-e��63fD\�����~��ʚ���Eo�3��1ET�Qn�6:�;������7�_t�p�(�-Е@^t�S�;�t�R��P�v�Y�ջeW/�UAʯ3}�5|��|�I��� ���WN���D���#Q4+�4�>^����zn���������<�y)�vy�����7��r^� ��Tn��<ߝ'"E���9`}��������#|�b��S4^8i�%J"P�8�:U7��n���7�4�>_uzѕ��Kc��G�/�D�Tz�d5���dqk����?��(�-Е@^t�S����3���e�6�6[;�,w�ŀg�޶ows �}+mӨ����Ħ*̂���y�{��W^}���^����M i@BUr��\�U+�d�a�w]�wԐ�ꂅR�PD��S��ԭ�I)�;vx��\�K�m���~�Bl�A଻$���=�J�@��[S��JT�#��+��!`]1�;|�?~��{�`g�7q�{�Ң��!rY.@�VlW+6v�K�p!�M@[�����n���[�ڔ�w?Dy�i�s.�[u��W�����}��{�����wm��x�棄v���#jb(NU ZJhΖ�qr��xG3$��N�`��=���ʼ�<�����-�����X樴�Q3E��b1A$0��^s��8M4�>k�xf���qp��9D�v��32�T�Т˃��^Z�a�l�A��I�ó��E�
��z��6��*:��՗WCtq�A.y�a�] 1�ƙ�ՠ����b�f�m��n�x�����d
u���Ln��s��{����������m9B��ժ$�*Z�v�-̬c��t���@��c����G�B�ܩ߻���f�0=��gy�f���L�qU�cT�jS9C��T���I%w�}�J�A��q�����Z=��R~	Q�W!H�b�1jW`b�eNc��zk��ܮr���_�?E���u�j0�_�Tz���<PWR�7�w���34<S���%Q���Jڀ;]*��w+��\�+�����,=�W�~�Hf\U�)�0�{m����]g0�����*k�Yq ��&���������t�ϽP5��$G�ٿ�L��u��� "���b*��/������o�n #���
"��$PP�ER�T�W�‣H�s���?�?�AU���w���?�����+'7�g���������_������������G��������7�3G��W���x����������@EU�Yq�7�'������O��x�����?������]����<=��?�?��o���g����C��
���U@�"I!D�Q �%D�TI!D�eD��@�Q!D�Q!H%!TH �!D�IQ$Q�QIE	Q!T�RaD�	Q!aD��RRTIaD��X aQ&HITIBTHP��!�RTIEAVIEQ! ��R@�T�D�`�Q!VTI !D�BPT $T��BH$	��HP�%RB$$BE�%BBd$P�!��RXB H	��HB %BBE�%Y	XB �����!��@���B@��$P���P��A�$D	UH@�!`!�  %�%�&	IBd	R@�$!IHBQBT�$B@�aBP�!YB  	FB� 	XBA�$�I	YB@��� %�$�&@�� �	HB@�a	� XBYAYd	!R@�@�D�dDY�%E�`@�!	de 
Q�	FR �`YQ�$�!!A	F�fC��C`R!
A�F	�`V�@$@FA� �`FA�� �`�`%$B��a!IFB�A��`!B�FdPeA��`Hd�bDTW?�l�o���ؠ"���?��sۿ�c��C��������"�������:��]?��q����;���W��_����_��~���� ����PU��"5�EU���F��]��*�f��[����?�������sw�ѳj*�_���������"��������������Cx�"�������"���_���坜������xk�?�����s��?�n(��:.��$�����_������������"����������W/�������������J�������e5�ߖ� �e�!������������ 
������.C/3�*-a�>{�  E( �U T��:�� ��.���e���wi���-ۖ����>��
z(z�^�*)�ơ_K��lez*���J���T����� �JT7#F�����2}:������t>��w��4.m:�G�u����`�ɠ ���C��>V��5@��GvW��L���� ���uҁ�7�cO��y�N���r��u�ݝiBe��:|�>� �wז>�w���u�����zz|�R��P  ��U 	P�1ER�� �hd`h0 ��BR��b10 F`�  ت�L�M2 � 4�   �I�))L��  @   �(C�	��M4��ji��驔�FĚyM�HAR4�jbmM4b42z�� ������}<��nG�UC�M��m���ـ��s�C�x���EEE� 6W�Ӗ��_��=�( ���QΟ��ݟ˻�?�ٱ�g�3�����?矣c;�gfuy���lgO9ǆ��#���z#�(��=�.�U
�V��p7���������ET9T�������D��!�n��T�d�j6^}� �a D5�]��x�����v�3ǻ��������}��/�ï����r����ŮC�tۼnۧ��1�7P�6�����m޶�9x��u��7Ol3\���9yN[��%˞7Q��9m��t��Z�kZۖ�PjM�D���R
jM@�Ě�SPjMB����RjQM@���A���CP�jAN!�(��SP"jDMH�J��PԂ��R�q &�DԠ��SP�j  5 ��AԈ���5(&�DԊ��R�q�QH�5 �j���]�6�R����RjR�]@���5.�5)�K�MHj]I�k[&�Q�թ�7P��n�˗M��9s�Ss�9�5��R:��:�P��ֳZ�\N���Z]�����������g��~��!�:�?F �	W?m�����a��u�[�D�JS��V6���Q�w-��M������tn�-���e҆�4ğ8�ʕ��o~����7q��-L��0�!�Z�VR��|PX�q�L]�q] H��,��m4��P3�8LD��8E�$�q͆�J�l,)��
��4TVF0�vBHa.uD!�B��M�e�DHK��C�e�e�����PR�6h�~w^i�(�nt��0�j%	\b+d�6�-�9�n���G �NGI�$���oYu䭕ش�ā����(t���k2����+F�*��!���_!u���f����`����p�%Y
���0���^	�<&v�P�͠�������]�th"���ٽ)A�Ul�0��<<nr�Hr�"á�J5�B�
2�	٫2�T��̂A�Mh��8se�M��&��ʴe�	Dq%x;.j�2FH�Y5���m9e�����(�;�d���$ȅm�hA:���9��-�3�y���󷷀t�)����4]��M�I��!M��y
�I�w�w�7�9�mqӐD�IlXA���ȖLr
-�"-�����#E�� `�t�D
K�hְ���P�vGNnC���9�%]���<i�4��4�=-�,�57�6��H��Ŋ�ꀱB�uh��c'��W�Y�s:�LK�TH��)�$K�q�D���Ͱ�d��Q+���7B&�+��/���ab��/M��&�F��{V���U�ɍ�D�."y� ��l������B\!ڮP!�Ξ��'Fg��m�� ���6R!vS`��J�E%�	� �!��#7�J��y+5�X( �F1��!EF�5��� v ]��%p�%��+`u� ��]g<�%w�m�F���O��FFB���mK5�Y���0�qWA�x�W����:�:�����ך-w��`m/�풬�t^�*텴J+GÜy<���!�Z-2܁�p��6�O;��|�
.�4cf�F袃�7�=kD!EmwE�6o���Lo���!��a�;� |9�&:MA�8/�������7����1�4	,��;�`�TB{lf���4NՉp�`�Ѹ�X2sK�_�f.�������c�a1�B�Ie�ة1h���"��a�/�(�]�����js0hchA���D!��E�؀X�V�@�&�A,dծ`�h$��9|ƌ�y��)o�o5�Jā�X1� ���X�I�h��	�;�=�]60]���mK��;A���;Om�4����s���^wn�9٧a�n���=��c���{�n��r7g��{k=n {��ĉ99TMtJƵ'Bn]�Q`!ߧe�9�&+7&�k���K5g69���a�U4��wi$��f&䣏�0�ph0��:�M\F��eH��mS���P��`bu�w�{4O2%��Y(^���GSE��,Y���U����Yxuۛ������:0���g�ݞ^}�����!��M��5�/����{��kz�~>e��C@(�8�N�8�2�m��RCZ=43m�n�ي�dK�w�7��V���.@&��b��y��+�LM��qX�<j+V/5��-�o,R��t�cݸ�����`�X,we��`�X,��m��m��`�����I �7wl��`�X,��i6�I6Ҳ�/-��'�$�]����`�X,��`�X,��`�X,��`�X,��`�X,I���	�`�X,��`�X,��`�X,��`�X,��`�X,��`��a$�ad�
��`�X,��`�X,��ũ6I��ݽ��X,$H,��`�uV��$��`�X,��`�X,��`�X,��`�ZM��M��,��`�X,��`�X,��`�X,�͒H$��`�X,9���X,���.���A`�X,��Q�b	 Z�)��d�]S����� sc�y۷wr����'�9�/Uf{Tۨ�񶕝���T��β��|�`�Xw��@�.F��Xl������ai��<ܩ�#N0�`�4m��Jpog���)���B��u�L$ ��Y�Z���k��6`�wxP���5O)��j��`�Xd�UfĬە�O�����]rO����mf`�ff�=�y�'u�x.;�3��:s�$�wt�7yHy�<��t�VbԎ�P�eeksyb�Ns�^���:���R����W^1��5�{�����ν��ԒZ��pb������܉j���)rI$�����۩�L�cy���̢�31�6-��̻Tq6L����z�t�I3�s�/��K�9ޒ������\e�i��5��ev�_s@�5���j�-쾷�p�kΡB]�st�HA�޵�9�-�xec ۣ������Z�N�D�3���Yɱ�����y&q�7Whؔ��*9�9�>O2�9�n^��Zӷ����h�MGB�<%�̝HĔl3�$�ۨ�#,Zn���K�rpTh�([$�{�cwY՘N����ng=�웧1fq��.��u��o.<����ii˹�2�)IQ�=֖Z��N�#��ws0�Y�36�,$�� �^p�˲��6��ի1�QM#�k�g�����]�/]� Eմ�$��]��ҫj�����o��\ո�^�ze޻�1�cǸ�դ��Ӕ�̣i^�vI7�,�q�y��<͵��{*�
��̼}�K�˺l�����s�"}wdݽ�7�_h���9{�gd�"��ꔢ`v�v�VovN��9��M�,�F�o9�<�$���7%��9o����R�z����f�KU�љJՙ'�i+'P`�*�����q�=׻�"CW�\�#�y�0��]�v4�V���h��8Y��H�y������e(H�3]�ۉd$��.����.��ͽ�]n^൮��XuR��,c�Ӏ��Vʻ�QWÞNHM}k@$�*n���V+\�26ի.U��@-���D�!�#P0�(f1��Zy���S�V%���cדLθ����r�M�����z�o^U;��G5� ���		��`�XKM�$��m��i6�@�X,�j�0��[,k��`�$H,9jZ �L���s,P�]׭�-ַ�6���qa
�Sy'ň(� =�@�{(,a�[ܒS�s�y&ծW�n<���wP�{�l��d޲$H-�N<V�N�ܜ�^7qe�m[u'GH��fW^k�x�a�[KKLvi�+gVt� v��Gf��=��ۉ�x^8��8�_h��h,��O&�ǇD�D�;��^�]Д6�f���[�z�=�����v::�}�dĽ��-3��h1�����!	�$P�"e8cz0����D٭Ʊgw�����4^��dw�
ʔz�S��d�n/k��*�k[\Y�{ �˙�ň��[5n0�)�{���vv�{q��vߌ�K��<>q���-��֏X����t��GA�aʀ�\1�c� �@D�>6l�h]��۷�W�����]:�������"B�I� ��3(��q�������?���/��  �������͢"����kH��9�A����ǰ�v�8�|����P|!AP�J'��������s��Ўz\S��#��C�(;��$ڂm!��L6���#�����T���$bh4W�����_��Z�"�o2�H�4!���xP�k�AE ���"x ��`U�i�+H�YOC�x��|���8�������z�	$�F 4�lh-*�(ezz�uX��.���P�`T�mb�hZP0"b��U0 � ��*b)�F��A�pM�p��lU q1X�w|N�W�b�<#��l TxC��aPU	�a��w�������Tu���@��x���x`�so/�� ��A�)VK�����)Ͱ�,���-��"��QD�E6�����2L�9��wq_2���蓰H�$4�F4���j���Yxj����1���K&�P��ՊtuĮ�Δ����n�un�WOc�����Z�ͬ%�*��ؼu�+3$��n6 �����_n�7[k�m�}��n�o�||gY|��4B�/��f�_Y~C�(UСE�N�#�:�")B�<�6�z��]���R�v�J�Rڳ�݊qF��Y~ľ|�W;�RZ)�<��8Ԣj�k�g~k/�7���\�u�������{�m=ݷH`d��sHj�h�-�Z@�{���%Gn0b�7ycyَG���py�Gb6���ت0,ܐv�g�ܓP�m3�Yˬ$��@�[�təL�A
�)����K�UUU	;�V���7z;�*�7�FD� s��Oq�0���
޸ws�:��/w�G���I�\���e�PI4L0B! 1V����`,�u��5W�2׶_��Y�y����iq�ڐ2�4��2a��;����y�ݘ��^��
��W�䰰��^���������M�\jfʼ1 �j�HnQ��}k���L�g)tQq������i	B	��7BJ4��T�
W|���Ɗͬ�L�d��L�)i4f'�cRћ/{�*���`�syl��[�3���>��pOx��#y�{�􍴓T&��x��>������'{�{�ݸ�*&�D\ ${�����{GT��0-U b$"����.���[�=��5Y�͡�VdT2����=��E"B�aJj�^d�"e h��83$:�3a�&�`h	�9Ȅ#���Z�UM�n�v��yÏu* �H��3��F"���w9x}B�@�����s�ˈ!��@�·�O�w��������
�4�Wm�ڬ�{\�j�0�h�H��
�y1��0*���2�>Z�M���$"�f\o)�B�[U�3Y�^Mŋ�x��j��DINh��N����w���緇�<�k�_]�m��"O;;@}>��臲���v��#Ѻ,/b �E�A7n��w]o6Cm�Lc�go�呓.�
υ
�YG_F*�d��1�����q�1n=��D��{ˬ�(L �}#���s��l��q�$v8j���A=�L��U[3:��;�8B���a�C�����*�*�ag���;|&�F�����"	���i3P×�a�VI��,4��y�Vkm!_��A�*Ӥ� ��[\d�����a _��Q\��"����9*D �N|�(�7R���?�(4z�hYI+wC/�dMQ�������,�%2F��s��^�Q�Qx�D	fR�!�5twP�`�%�@Y��5an*v,�E4TMD�{��(���y�D�)����j��s�X�(7=��d����""" ��1���χ�6���� �����g�VB�tp�c���qYy��g�#q6�j��&z��k��nF'b�[��0�p{n���q�P]�d��S�.�z���n�D;���nªxd��k�&� �{D�Uٴ>
ey؟n�T�.jɊ	��t��G'lG���Ǟ�~������x���D�T��KA�|�w��8��9RX�C6kv��]�� ޢ�����(�F�;�!�h9�/s-q!�=�Ԉف&���N��CO�P#��t��Pda:�@�|���Ui�ADx�o!Z����
��>������.sS�V�P�
�X�N}X��9 ���!Fd�;�[B�y�
 M�Bx�jCslx@�H�F�Q�"���-���H��0�y�+��fV�Ț�aZ^�B�զ�P�M�ے�pi�q|F���R�J[��ڠ(I�B���ܐ�}�����οP�(����*V��T�λ�7W[�#�qU��G�U@~J1bF'�m�Μ:E�>H��C5�PeL-��v��>���9����{x.�9�خ2,�{��éaz�#M{����b���W�|m��#�F����X[� �l�څV�f��+��|��U��G"9�Qn�1N�{�Q�H�,oUY�� ����7z~�UMt���I���46B!�C}�m�؉383��-����0U;T.KgPj��<?x�g�H��a��|��g�����rg�H2�G�\T5ҙӿc1�g�UG�pag�C�b�`�m��:A}��*�$��c6�0���-�`�B#
h�acuS�7� �d�\�xN���+��ϕ@�p���k���ji���>(��GP�=82�e\(�qD���������9�8�-�ت%��D�J2Ôj6`rT�!�[|F*���о�a�%@�=�i����`D@��W:Q�!�7��iwɈkO�Fj`�w�w��Pp�"�W�V�j�nU�@��,�`#�!��}�}�%b��V���e!����+�#uY���Xx-s��B�	����n��Za�T����g�|��n��;An�a\����U�,�1� �OFzeLl��G�F��P���Q�z�"*�A��k�c:�rK��i7�J'�C�CS��dn2I�����j�V�V�6�PB�U�w|��3�H$7*���B�k���)绣\4��>X�2���§�V��Oz��n48zE�AUG�b���ЬԊ�{;M�Fye�qX=�=���Y���׺�3�i4LN����� ?uW�;��~��d$S���h|�a�B�|��HϹ�']�f��B�[;�|�������\̗��5I}�7`P�K�Y�`ദAaR�ⳤpuVy{���C��|��G�8K*|3���+�`ݴh�D %**����5*�D5�3|L�뼊��P�����(�z�ָ�*���Y�Ꚅ3�w-ߵ�����9*�18�n�A{۰w�����)\��p��];K�gv:G�V��Ln��FFdP�����/]���;����ah���2�Lr��NAB���$�ʖ(Z-#���Y�����p��˕�o���O���� !���W��t�#�Ǐ�)^�P��G���+�*���=�̗!�T�}s���Y)�ϋ��H��<�xV��w5��j��� <���C�\	�IpO ��/�W�Zc�j�
�,%W �&���p	��w���42�r��>E���	a)���X�G6ͭ�HU�N֌��^����J`h��#^� �ٛ�	��̽mn�,�l����F�GYE|<Y�w��,Ӏ�Ҿ�.	2� ޡ�U������ƮZ��8��lst��s Ƕ�b�;�3g4�v�[��]���E�b]��R˦�6�z��;�.z��e����!�:�iU�Mջ%����}�}]x	�rA�����X�%L"�(,���@f~xQ��D�ڨ`�+�| �<a�^}�s���IG�n�͙*]�Uf]U��q�T�ڛ����U�D.3�E�68�uK�"��0����"�4-���y�҉:����?�we(%��'UTp֖xk��[��;�,M���K�?'|��3w9YJW>`��z@�/��h� D���]|�YH�J�W�o��QH%��	 �`�|��y��䒉(��_2*]�J�Mm�`RД:���R��� /�;�&��Ը�*/n������\^�abb�7vh�j�C��$��H��Q
�e	HRj�`mr	�fT>{|�K.���$R@��K�H���!B:F		!ߌ�" �t�����"o��ޓpI:
JK B@�Z��w�$��(2	 �U	" z� �HEK��5��|��e]�1	��O��E?��p�m��b;��(R����&�&�$(���$��E�v���15�<�H���l���)HE�=�m) s��p*<���JCY5�H$��rE�2�.V��JMm����r�� ϟ|8h�K��A$��(;cqI��. �;�7�z�G�" *A�$@�) � ĂQ		�Bv�I�u��|�w�&����9��j��(J�!���A�$� ���y����Vf �UPտ6�l�9E`P�+��$Pi)"'g`\RBr���ڒ�_32���B\R@�J�H�U! �'!���A��H$�إE�n�H���e`j	 ���>@�&r���	�P�!쨝�QQ��w�f�WY�JN�16��9�OX&��$�v�	��7u��vCq
�+��L���&JR������W������4�P�L�����k�9�#cQOnv��,���˘��x��R\RG\��t�5z�$�����Q	���Oj_ˢ�]�^��`G�
RA$MM� �	�;��oA�3P��fQ.i7�I�BH��Q56��|��J�R�0�	I�J��L)k�o�	�I�R\ O �	��J�R�!�̠VE���"\���5��) 2D�$�Iڤ$D��i2!#=��4�om�9 A�jL��.V	BH=��j@��ˡ$C�ߧ+F�\��N�H$�H}�~_˕Y,�.�V�紜�	"�E$O"TG����$��[�7YGfsN��\�� vc�V�;\�`-
1�J� �!F�S�ؗ�����hJ��d%'H4#ndRA'*���dJ�N�;�P���rB���)I�kc�����$�rRԗυ`�	 �%A�j	R��ȗ�p. �5<�T3VdK�>^�5��0JR����t�23�
NRTND��ߜ��T��E$'��d�zҿ!$a6��Zp���dR*H�'�J�����F�jYZܩEU/��RD'|�.# j%A$ʩ$D�(n	"o��t�P��.!"vy<�C��Ќb!uR!"�&���H&���]��fA�����		���&��L�t-A'��qI��.	#��@o*�,�$@�����	��dBU&�\EM�BH���u��7�������z{���Kʻ���}�Ț�! ��)Q	���Hr��\�F�ޥUeT�z�&𔚓!(N0�)JN����)"��@5��JѸ���	��hu�d�$��PuZ�iJ䨄�H�A��������*��9yJL�A�%)�b���"�M�u(�0I�rB�!Օ�%E��9��^W�����R}Z�@���	I�9'92�감�)5q&�ݖ/<�ߞ�)�%/`TRA���e��̙2�H!��$C�jC%(8�bm)Bk0J�ݙ�ܹ��We�%m�"k3x�H'h�=�D�%A�hl�5�;�/̗Ug$�Wk�� �B�J{=�B��h;X��Ͻ���kY������53�r���8pW�
�
.ޡ�A�h�q}���~��d��5<�m$*�ˉ�`Mtn��WD��2D��2r�P�U|�r�1��#Ɖ��>�K.8�>d�#Zj��0"�A�L�poUi��PC��������䯈��T=����&��|畗z���5��X~�+T�cX�cI<���)w�w݂�`�#F*��G����ꮰ%W9Ɓl���!����f�`�6
6(^ø�{���ADȺ.>ph�H�Aj�<Є�Q>�vt�B�ul潊����Y򎄮�C�L���cw�c����!iUR�=�th����4�?|�a�8�!j���������qBPD?U[�����3�N��K��;��3@B�4�u:�+(y�c���k�|�W$6F��P�z�5�Ϡ��/�URU������@O��64�|w��Xm�O�Wp�tx�hഄH�!�dM�8�ZI�*
�}k7˾||�X*Y�-kb�Hߞf�nu�QBP�Ag�燓G�+U:ZWN��P"��j���'a�I��1#	��c*��A$Io^���=	~~��s�^�LPOEBɎ��d�����"""0�DJ���DD@%�U��=�իE����ϰY�n�2�Y��Y�aI�u�E���1�2�G��#��m��`�qPc��z�G�Ϭl]�e��u�4��{�璸��C�[cg�n'��"մ"&��&��^c����ж���;_^��O�#������c�R!�>+�~(*v� h���5���|K�#�B0�;1�@���9�:������q�|��Q_�l��|�ԼcRv�$�A$Q6�|d��H�w�?o�5��0X���gM|sU�w�}�C,Q(��#�P��9=��/'ǅ��T�X� 6����&Re�4�ۚ���+��de8�άV�)�n�����9�
���#����1��ȼ�F�&�+�"���̶�c<m���8�%:����1��	=qu<s.���ڃ0�V�IcU����Ma��FB\�z� a� b�{��r�H>�5	&�$&_tz�A�j��J��(w�d5 gw�%��	��m�����S6�=A�z䓄��g�;�|[�����꫾rݑ��G�� 0��^q�ϔ�=!|h&�]#Т8s�˖�uZ}�O������"\�R�A�:@�c�H$n*�C=��e�<{!�cM�e�&�h� A�
q���2��ֆ|���%f,� ���!F*�%kF�(�Q��h�O[��P9�D��L�F�}�*FCq~��t�u�����U��W����Î'|탆�E�ռDU�S��6��O�#g�ب1<�[$)s�1n��&����Y�5qi�[�%,��s��i6< =5�!�\"ߟbL 9�ymO!��s�^ʆ�t��kn�QQ,��(�F� k�_��e�b��E����c����۱p�]8C�4�#��>�| �7U"B|��&˞�^�<8��p.6:�f�d�<���Q`p@�@Tݪ�E���P�N���mu�\m"�V��Y��y�1�J�a��H�f� �a�V��M;CY�: m��eD3q�p���:G��Y�wc�8kH���'	ޏ	:���Z�r����9��s�x���o�eU�$����W��p �0����V��7m�����݈�v�����c��~��=xjb�Ƈ;�p#\ҁj�|�4����e�����Mf��a��:��~P�]�|�a���!��V�q��2���>#U���
�	6@�Udg:�]�>��b�O0
 ��w@�#!�󻿕]�9r{��Ԃ�������}���ψ�?Š�3�d���y6�w����*��\ld��)��$g���!j�oP8y��cJ��H桤�;SDF��(��f��
�!����-0;�8>`��N�U�5� +8K�H
�}^p�,mf�]
Y*��1���{U	Æy�KcH
!��tbTD�܎VXg��K#^�t�^<K��I��UT"���)'�qH"���)�,d�u����F�d����J�IB�ߘû��W�R��Ͼe(J�(�O�n�Ŝ��9���� V��|q@�c�:��_S#H�_и������ZG��k��j�h�8C�&O}$���,�ޠ�b��>���� ��� T��2}U��6jFn��7MT���-�W��L�i��Q,.%���H2��B�2��LloSAARf9QAE`�7���N�L�2+�e^XaK��3�]��`��V��j���ܼ5[UJ�ն��+hݴ�wk�4��Yv���]NM=��7(I�a�qֱh��oZ��qeQX�b�)^g;��1�V�/)燱\ΰ]!�`�ˬV�8��=c�4��z��{�듢ﯾ�%P	�*kKX�4(=�H�ɢA���D�4��nȵە���\����~0�74�Y,�x ֺ^�h�Q�4���/������H6A��Bl��B����P��_T>0���y#�#���l2����I��i1����L",��H��i�8Q�0�Ďq�.f{��R�=�$� IB0� �Y@"�@lv��M����73m��JڳNxg��lP��dF�V���6E���2�>p4��e�8G��%#��Ĝlȡ���0���B#ӏ�h���Q��t�ӷ���*�����>q��Ōdd$u�a�U���7	�>:�M2:Fj���Ȇ��vt|�$D"j��m#����@U5v���L\k��:@��<��EY��C5dv���R4R�}��b�ږ��ڹ�nW�w�1D>@�+5�Ӗ��
X�v�O��(kT�k�̼��W���j���'���y|����i*�5�~"F$)1����ǝ�|�r]|��
0�����#��5�?d�*�V�a5��h;��cő�H�U�W�]�J�.��h��DX5tl����jC���kŅ�s2�G�;�-h �ow�oz��}_z�+Z.V����vF�H��\����Q}us��
�8-��8@�� ��f}�t�6A5�P�+,��B���\zU���"3Uiӄ}B�8G��]yn+غk���%0�`��C��gPg-����A
ycHFjBﳂ��C!y]�6�]PC�a�C�H�<&k���B�o�V�K^n̕�P�(����/�8x�3Pkz��m��,E�Ƈ�g�E$�����i��q�5�c���!�_U���t���~��̷�aS%��r�g-��,d������&%V�]u��W=$����3f��8�ﻑali��?��l��q��ه�4!$h	-�X-lm�7��	!|�8M���{��3P�3Ͼ����<"ؠ S5�t��9���:��<SP�����1�p��7	qH�٫3:�<���<5p�iG"rH�1�M�T࡚ �Й�`2~f�>�4X�5�� >5#�v���13jX�\ }B��!�C���@�őmO��j�4��P�����ku@�C�@���<�|F�L��HIm�'�C��/��lLUQ4(mӟ�Z�b�T��r��x٠�B�e��$���;�������3�Wz�I�y/�@���> ��4�j7�#�VsP|C����|�qm_��Vht�z��|��+���"�QH���q!�s��D�6hZMX��p�Z���3Y�Ǻ �(�H�h{y"g$r�C f*�<7�O���D�UN!���`t���*5"9�����Ǧ�2@�a��ҩ�4o��p�������]��3X@��� 7�ޗꏐL���.�-5�#@D7ʢ��Cl�!VJu[���6�JaIYf\e�%�])v�J���	"�S% e]���v�*�e^ BB��A-*�%Ы�l�N��@�Z&��x�׋�����^���
�ssa�(7
m2DDDDZH�s'DDD$�Dm�C` �BVf���땷c��x�����7bMm0�vYՈm���ZԤ�e�Vl�>!s������l��ޓ��*m7!�l'n��D�:@��M�mɮ�[�+ �Khvf\q����{������)f��˲���� ����l�6�����M1<g���v�a��Kl�~�M�e�-�D8TC#�3]��$3|�m�x�܈�y�^\ Z��J��H"ـ`!�	-�^9<�H?���a�3�{�|괐��ӥ�#ݿ�0�9�Y�ha��~#
M��I�xZ�D1*����"���݌<��2�0�O{�P�a��q8���X�P�0���:ZZ�̷�$AD�-�����Y�D>뫪�CX �+�lW���6)�0|����Ⱥ�F���q���a����ʹ~�6�A��֞K��TI���M��,��q��M��������)��A��n!a �hH�C��1�� ��>���[l���&E��A��D�`���hB<B�Y�m/00��/T(q�}�/�!]��h�c���^� i�� @C�#,p
Y��k~��{�q��6P�]Ph��#���m��48N(I�g�'��7`B�0������,�X�CB�B� �*���Vho3�l��("D@0a�C E���$�:En�,��9�r
�o����:�#�c��P�V���y(ea+WTH��P���C�3��N ��0!¬#z%⻑�QW��|��#�Ѩ�$�����&;�����P�������}��b����(�rV�紧�H��(E�;d�.(
QB�� P�!�֏aa�#�w�"E#���8��8[ztp���K�:G-= �x��Xzf����a?}� (�|*�x�����B�5�P&���;@����v ��߁a�ajL�ל�Q��'瓊@�XUR�U@��$��;�&�Ȝ��')�� ����	/�9�i�L4�-�P�A k��W&Cu��*Z���_v�+z��A}�8-YH�C��V��-��,3��C���A��R
c�)m����S��L�3#H�r7Ѡ1n�ЇI�x�������Mss/ҋn��6���2ʶ0���Ղ�B@�p��P���fIA�im��0�X��w��]�D�p��U��x��j{4�މ)W	#%Ԉ%�J+��ٱäB"q��'�^�:<'��BF��t��L-XW�v�E+(8�X��zO}fG�j��6C4��Q]�E��>����"����?����T�۴�<ty�ƕ�ڴ��g�=P�$($�G �\�$ZS��lVa���'�.�X�����dΒFlP�n��B8t��>�i'hdU�g��h"��BO\�G��^i���x.U]�C7�(�t��>&k�����i��I!K��"?�o�F���`�8IʢA�[p� V��)��jP��H�M�b���sm��x�݈D`�L8��d����q�*C����&��/P�ITB�F��|�EQUӆFAm���@�L
���cEH���R�T�$��R��E�ڪ�(�ƮZ�����Uy��a+�����O'[p�u��뀬�NQ�6-{�����Ծ:���Clv�\Ǳ�����=(N|vrr��v8,>͹���7k�zU�c!Yv_��N*���<�f�)���]������k�����x������ۦ::��|��j��Æ6���,�� �=�'�J���=;���
#Ɨi�8@�[�$7P����܈y�8E��[���@8F%Z��D(���v�4^�z�A��e��ޏ�`��z7*��k�OB]��C�<˯�Tj���i> ��P����xP�G�k=�@�-�ðU�_9�N���e���\"��f��3Xa �7��]���H"�Ƈ��HeC��V���{���q�~4=��P�I�W{��!�7trP��Eʠn�P�Bo�˵�s��n'�ߔ|���u�]��%Nݽ6C��}v �8F19,ޞ�bmFk1L���iF��y���ҝu:�J-I�K^�w�HqY
ۭ�>Ľ�#�ғ��A�dr���#eA�m�8i�R!��е^!j�*�3�H}vn]Y�\$�,���r]9�CZG�t�=��2�k�u�C��l�'`�jo�u�z�s!�@Ρ��n�0N��z�N׷V�w���G�I�D�c��p��a��@�e�5g�T~�>(�Gz�iWH��ȇ�<p�5S�x��Ґ`a|�餤F\/.ԠP�l �L$`P>��`�3k�B��Q�D5*��%��@(Q��ױo�r�(B���*���A>�Jmm��}�� ��{���!�B�τ�XSH=��S6���E�w���{�-b"�b��n��b��1U��B͐��@1�%���$	F*�$��h���H(�'=T(U���LoG��G��{��r�o���A]yПUd���ϝ��v���=(BP5k�O7�<O>wYv�vf���N!mB�<�@YR������&��i#�lW7��n��J��3,��yK�{g���J9�hܿy-�kX����4��w�P
�I�_|yΔ�N�7;;Oj�� �P�(�I��WcNx�p�ذ����2E0�SH㱮^WN)����_s'��^R�{�<Ku�ۛ��}{�,}�g�>I�!��`צ��Ad��D8�4���zx���M $ 9�r����Z�Pŕ�%��g+}��3{��\V�F�u�1�8��Sdq��Lc|u�>������n� }/Y$��Vtĉ��}�i2\���ɯl�N�I��-��kTi�搖k����� �	R����0 5@&��h�w�|\��.�7{��a�
"�*&@mQ L�DDD@E���DDD2@%�^�Nmqu��k��m�U/6��]��p���E�Gg��_Y�=l���z2v�ʆ�رmƺ��lr�r�i:��he�\#WK7��E�C��M]i7j3��G����BC��H��WAV�U=��DWhxG�ĳO���� 8=�z"���`\s��s����؆�v��f�Ϲ~�]$���&?o5Lo)��N&�U���*A?:��7�H��Q�7޺M=uxe��I)��SD�K �;Hz�l\�#���dI,(ڈ8Y�6Hr ���n_3S>��C��a�BH���pI"�!@7;; �v{@�rt�b997oh .I���K��B7��y�S�(�c6��M�A����y|ɐ"Ϊ		W�F��)�'Ja@�K �q ���UpW9�É4�mc9���TH4��b���i�;�:@�o޿aig������桖���D��%�����).O�}��ﮅUp���FG!��I�UK�՗��دG#��4\
">�s�> ��D<9��ĚĉP�X�����UM��1�:�/EUP��^��������y�c#qπ�����W7�G6lih�>��L�O��,bH-ȣ�z��C�v��Zo����gf���e���{�@R���@L�nݻ��-L�\�j�[iia�u2''b��trgW2�p��R`�T�B�>�ʹO"��>��}S��]@�I
H��v=x�����ewu��;}ti8���*�}�8�}�>_&�J'#1v��g3�JRH#�0�H\%��d�Q�][8:5�<������p�-�HX�����ř��rQ��of���i�[W|�"X����
�s��.꬀芳�*�0m�đ͠9e'��<^��������?}>��g���G+�,�,V7�%�EJM:�3�U�����{Hlu�>�p�]^���s�"�� �Mi���m�� w���O!�	�Y��T{�S4
d�]�ɐ�*2�
%�0I7���xF	w7�v鞀�n}�B�p��� �B ��z>L��d�%3�4䫙�r�9oK�h��N�Wk$�5�E�_s1�Y�2�4LO�dx^a��h�)���oK�{ޢ�f�k֙5-T�&�R�Y��~|�;=�Q[xx����H��7����|R����"%A�DQ4(�3	�.X�ҼRj��]W�1�I�.ԑ!�����sy!�&k��ؤ�,���$]O%!3DY
6n��@$�7S�L����df�VXg;{3\W�l&��OMK���N?�2�-2=a�V�����&ꚫj�]��������a:1����]7k���7k�n�E�ُs=��������m���;��sdL6��և<ij�%uq�]`Y۵v�۝�۝�mt���Su���0��;�����7��	��/N#GV�x�V�r�UV��W�����9�l�hk�1#�D��hA�rZG��j�%������|��9-`����"u�{]�B��}}|�y�v� (0�B��p�sl�v$6T[v������},�}��+���0��«P���v�Tyͥ��j/8�>����RL�m�C�Rm��,��9������9���xg�X��u��&�S�$� �\^��3s'�����I|H��V�BTR>D���32R�-�t(�F`��9ۛ^Fw���_����2V�r����
�I�Ji�N����T�k��S)�72["���Ub��N��<����P�	��3i)3�>X��n�"���Qu$Ǉ���E����FĂ��5��o"E>�/֭}��uu��k������q� h9�m�j�d�v�Y7Ҙ�ӟ(c 5]��E$�b03:�~�y��`�'���r#�w+�&9+0{;�(�J� 7g�~(�����f"?h8���_���CKi��<��6�F�=燪�@�t̳ե����9ޟz©��e��w�:��o�T���&�1Dh����<��aBL� l)��s~���n�v�"���%�T�� �Y���8Y�ɲ����o˱/�BH�l�=�}/3���!�qw6�a��;��si�GvŤ�6�B�R�)�&ߢ9η![�s�f.�6(`z�q�n1�;�x�-�]a�Q��^(�|�w�m�����~������,X�*�sj!Ծ�܄�<����ś�/O�"&��f���d�&,�˗k޻��ݕ�Y�o�����I
D�)3\�����U�T;�����o�9~���N܄d�ZXZ��e|v-�ߏ{�w7���ΰP��mŰ�<^i��}۾ܽa�r���x��/c��P#ޥ�I6A��r�:-��iҢ�O���H��UR�"ƟG�k�ʝA��E����$Jy{6�UٽKƒ>��0�����3ٛ2��)1[Mo��{��g0�y��{�fMo��w~&�`I9@=���� )i)�t��E"Hk�M�3d3,��Zd&��) �C��	��!^u{t�F,&�\K�5u�-ʲ) J���d R!$,ʲ겦�*�iF��, �4hh�fD`�.>�Gt���3��frL��g"2DDDF�Бq̛DDD Oʀ�Ei�q���s�z5wn��Z�SV�屵����ۢ��Eg��n�j]=Y��n��*/ccۉ�.��{�WA[��v�ڏA��{y9T�X �� t	��=����󽧳�f�j47g��F���׽�������}uB�.�M��ؖW#��nt�혱�R�o'�iu{�d�'�hn��O�D�A���m�)D4E*h�Cݻ��g��c���xC���m�t_8��V�w�u�B������+�M'�KK9�][�������P3̵�Î�t4(o��/u^�;о��N8�}�=�d�c�W�E�M4ˤEf�gvd��H����ɖ�}I�	�p�P�]���]���;�.��\AĒ��,�h�<�$�←�2�(��W-��G=��tQ4�
t��F�؀�<�X������x�����)�}����R}Y0�E�M-�sz_���[��ˢ'y�����,��,�R����39z��h���n���}Q i��the���9��#E�}�W7VƏCĺ��`[�R���f��5ۨ�"D� �M�O'oN�SV�	�l�W�����m�3�)��y=վ����b�s���G9�-��33 ;r��8Ҫ�;:����}�B0����'2���$ңH���L�z*9�&�Z�@�G*�͎����e�W0�:L�[%�jy��Fx�ی�Ӛ1�G�]�����GFuP���� ��=��0�TQB���fs.R0��HW1��p�y�!��f@z�;:�����b��=°�����J�Tǣ`��:�xy��"� �"�=����a�;|��m5]�6Ol�h[9���l����|��1��Z��f�I��%+=��[�nƘ@ f*u�~�r��Ӫ*��vWD��DQ[O��c�A$�K�m[��z`t�r����[�Do#���r�X�~��Lsx���L�ٻ�m���3EP�?�=���C>�E�+�B���֞�H����61[;337��؃ա ��&���������Vr^s���׌w��$�B���Wd7N�*����/=|��Z���,����'m�u<���+���:
�� �cwv��(5TP ]���q��I��l�ON��"�vޞzmԙpċ�-��ET����(�N�|���$b1Y���D�^�ѡ@U�T���������<[�#ל�ioE��[��*x�P���
��k��� zV'{�9�������@�����~��*=8�eEUQO�T-��EC���}`m�n ���������ɪʦ�������|�����.p�#[\��	7V%bLD���A�	2
� ?%bU�A��v�6�RDM���@a
��2���(�0�(H���J�"!�P.PP�1P6�~tP	�&,L�<�$^y����� �(��LZ�$(�X �G�x�J�0�(�7�	
6�����,4"A@�[�*�dS�~`e��:����E��r��-]��|-�8	J�(-"!=u/Mlr߻�g������:�۟���v��ç�zy�_����;l�������8�>���>^~�~[{{��N������|��՚�Q88�t�Zw6;O.�wC��_Dlm��8�v~�����y��my��T:������~\��������#��ԔѮ�����TD;CyI�T?�8-�������3��_Z�����O��h\� c�s<���J{��{}���R(�*m��v��{^Z|#��A��@EP������w7>�͔�_ğy������}޿+��������$1SF�MI��xfӾ� n�~�<�%��Ŧ��_��5�NP����^������S@{ߣ��������n~&]���rȞR��~������������yuf;���UD�3EDQT@�M5�D+0
ĠD�!H�KDE�PC!�1!���"�"�(�B�lb��)��6�
d�D� ,�B�(H� �+ $� �+ $��	 ��� $�*�, ����
��J�"����*��@) 	"��@	2�, �2@ʨB�@�*�	*����C $$ $� �0 ��@J�@B���@B�@+ $���

�
L�HQQ)T�}x�!04L+����
LH�D@���R �LL�D�A1,�0K*%1D�S2J�!1�p�	���u!�J$��#L�00H̨���fuj��h�҃��6~��W���A���Ϻ��ln���~���"�!���@^���$�2�(ģJ1����={O;�G���᯼p�"{>��r�}y���h|���w�Opw�17�>�?7q�ۻ�7�L<����������������i??�(���Cbm1J�|_�d�����A�/���_�u�ߺ?6�twd�п֜�?Yv�77�#��7���w#�}'$��YO˟��O�����U����[m'����О��g�g�k�ۏ���$U��.�"T��1s�o{=�/%����C���x�|N���lu��=�w=0�$#QU}����{� <0>��?;�����o���f�ѣA>����
�-@TC`p?v�* ���c��y����69=����֏�l���c5�QU��pC�����wwȨ"!�yT2rh"���4���~����Y��!�JZoO����%�����("�a��Q���}%�9���M����9�����"�w�c����8��>�������A{8�Iۮ\�;|����ܺr�?w����?q���������'��O/_��o���={����(�~s��>�غ��Qχ�'O��x�V&���C6�������������r�?�l��{{ � ��U�~���UG�����{���y��=����tOh�~n��{:���oFN��=�c�6'ן�����n���|�B��O��/�~���?QO��_�k��ÿ��wb~P�O��|v9E�8��M���� �._��lv�A�t@EP�Ϸ���	���F����bX���ԁ�6���?y�t���u�طoWaO� 'k *dmDt7.����o��8y�����@�����O>�Hz$ Q�!����h�3��lwH��U���k�l���o����t ��?Y���??G{0����-����v�ޘv$�?�=!�=���F�tz���G��N��|ƽ
w�rE8P�qG��