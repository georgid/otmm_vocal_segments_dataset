BZh91AY&SY��Ǎ �_�Px���������`�\��5�B�  �Aq���n`5FT$P�OI��i=SM =G���� 2Q#�D�� h@�101��&$�(���5@    �"�M�I�1hz��$�F�P�S
z�(mF��4OQ���`��� �J��*��F�g��?г!x����(1��'��$���
�#�G�7� H 8Ѓao��a��o����C��G�̻�������������pn�:t�#N8p�,էw]��ӻ����uiØ�bØ�ÄffFfffe�f{� �&T:F�էN�#un!�f,;�i�7ww7y�=׀�r���A	��>��<#��ϲ=9$C�XI�^�4_!�ՉJK��umUo���/i���t��&%�������(NL��u�\�	X���T<*�7u�!�8�`fÚKS=�,׌�ON҃ɛbV��Μ�6u��^ĭfXb\�
�ٚn�&�L�r�ݴ�v:X|����<J�������-��i �v!K��V�/4(��Ӆ��-�s*���nn��Gv�q��U����Z�\�q߻V��c�qM8WǍoߐ��d3/q�}��I��Jկ=3濣��wgs2���V��f]�����fff���������%5��MuB�m�K"���&/+4���2�X��tS�g�-��X�H��ޞ�:Z�߰��@+�<W-xp 9����Ӿ��'u�aקob�[���"0��<<��.qcq�r�^�
���(g��\5ӧ�~���x��~�kd�s^�l�y;��j��.#�2���'��b2J�E�<z�31{QoWk1(��[�<�zC��v}ǝ7�g0�R�vm�;m����؁XQ��^��B��fx��u��PYЙH��1*Mf'sl�z3���x��x�@�@���5(Y��z�1�T<X!Y���x_&�h�a�� ��P��p��$������O舚#���6\���֬.43(vFy��V�� ]U�s�q���;�s�{�Ĵ��_ ��F���NJAS#9\"�i�'�@��et��ީۄQh���n=��0G`�C��[&K��!�ô����f"��(����w�X�dIGe�J9���� 0�i;Y؆l��S���x^ܷl�9��u���pHD[��^p�V��y�1���I��R_݆YItb�䦚̩�A}�|�����-Nw�����f�x�b'��$+w�s#V 9/0��Gz���.�mq�C�L:���GD6/L1��`y���t|����LQ>%0 �"�D#R���4*D��z�l�ʩ��^�-�pD�#�,����.�2]��;]H��"�D���NWwgU�	ٳ�#+�\�[�ELL{XK ;1u��+�v��δf��x�0R��G$Ç���t�݈q�Pf�!�9���>�;���"B�WJ戣'�"�K�y��p��̂�y��ۈY5~�X #ѣ9;��4�H�!�@��չ�Ȩ�*&��"BsY������x �b��[�
1��rw�&7���?xx��-�Hp	<ˮbk�`[��%�������\����"^��~;$���ob���w��k��;��y<�}�����{z���`��Wo�;x�%�z���o2y��E��&*��m�L�I��3���D�7�j�:y�g �2 ʐיTO)��fWb=wשy���Ȼ���ʹG9T��>���5�� ���g�G ��4���s�Ǘ��g��n@���%���M.m�S�����mv��.mk�]�n�ʙ��8���:�:��Yx+��4�`����vk:4v'�H {�|Fpr��C�*�ޢ��t�Ղ���j�A�da!9d�I$�A�C�9{{��s���=M4���Ӟd�&�u��6�q1Â�.��Q],��J���(�UF�����!�2�Hj.Q���ˀA�-��0�A@�*jk&5T�B���%�7��9dSe�[S��[E�(���Ղ���R�V�j(q�M�Hɀ��&d�,�FN6��:P�<i8�����&�T��n�9DdYSb3��Q#S��ns�N��*��#�v�?Ѯx8o]��I��83gg"��6p��e���I����f�ٕD!�o�@�	ލP��y�!jL#|A-(#��@�Dނn'6s���>d�+H��{L�.=o��?�:�;�i*�E� a��,%j�2x��,���a�O�;�\�4L�i���N�Ǎ��D�-I^b��?d�m�>�W2$.5��q�:�O8�ӥ�h��e�2���g�C ��I&"���"�Tb*EUX��"�QDAX(�b"���gP`�����`1�2 ^�_��d�1�Lv��!�����35��� @��A* B BH��2�cS�<�L�Q�W��o@�L��Xr��,���H����)` T7I'�J�o`�(�x�_*����5��ȕi6@ݨȭ,�z��ge�Q��Qt��L�l@!R�<�((k�>~{Ksde�G�� ����"�@�E��� �<�'y�E�F�y�`(_{3#�dwA�p��Sh�k�#��f"��P��3����4�^�y!b�h� '�� �,����N��'��)h;���jсS���֡8�P}���0G�}�'�AI��(�l2\o�!�JN�J��h���v3�l������w::yG2��u�C p`�Ph3�$�Y�~�=[]���rR��7h8�$0�,X�d�*ن󪟐��N��h����V�ɓ|C�5�tPp`xV|HT!Mj(�ƈ�ÑT(����V�E�����WA0 �C�i���+��1� �ŏ@ە5`����s2NH�R���o6�4^�"b�c,�>�0�gR�M��(m����rE8P���Ǎ