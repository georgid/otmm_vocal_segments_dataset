BZh91AY&SYHj�| �߀Px���������`z��ǹY�MW�  4R@���>��k�ml�a$!4�b��i��~�z�S�=G�ڀb��4h�U5���M!�  2)Q�      &�DS�    � �R����4�6�i�  4�D�!�2�O��OFL���C 45�Ԩ-�"��A��aS���U�	�$�B��}Re*�~��P2`�1�@�E1��"ޯdz��}���{ߓշ9~����������������%:(�B*�"FS��D"):!T�!�F�!QY�!���!���Kwwwwwwwwwww|��E8�^���rH��~��p�g�3甮 �r���2��%V��]P2j�`=��TB��)G�1Ѱm)��(� s.��f-񟀌�sx^��ʨ�;�#sjb^"���'
��T��nL8��)=;��L]�ۻ�r�)��VU�YX����Yu&q�?ȺN}L3o��L򴂥G��L����\9ʣ01�ƈ��y+N�ܥ��D�V
#X�bV.2�����L�n��iF�g������(��߇�񠄐�0���i ��~&2`�?����=��޺I$�Iffff$�I$�I$�I$�I$�33.ĵ.p�*WiQ0dӌb���tHT�<��b��9����<9��
�H0�{S��r�
��ֵ@�"�\�AJo��UO���ǡ�
�X����#U<�J�d_:��R#!�!�S�R�8�k���C�̧�˗�O�YER��'}�xF�U���Ã0h���Z����΢yX���@r3������i ��"v��R�M�mVn��J��#6m�%��mZ�]������a�B�PL��`��@0����raٱ;Af� �vi��fT�ACqw�.\Yx�#aـX�A.E����YӀ��0���ȗ�{Ȩʡ�޺XM���p�f+8,�ll6K�O_]��.����z���b͏΃;- ���y;9 �ah�佚"H�؋��C��q��O���Ƃ��+���ia�F'�|HE�^s��(Gq�����X�l�y���'�sè�T9~r"�y�yZZ�t@^�����ę�yI�+�<�ѼJ/�sk����m��v��8(	w�a*�6(»4�< �u�Gx_�F"i�0�$I \@|y緼��p2Y��Lwz�΀!�'��t�G!�Z3f�]0h�nC��a���jp
��rq�)����iNpnm��X��[�4�q��D��k<p��6��Y9����**��ݫ���(��FP�v�Q����5�t@N/Q�����|y��3���SAEb��$�f4{��к�ٓ�NS�������Q��dxn�ۼ�c�'F����a�-�C���[�jf�h�X[v�ri�UZeqW]�� �f�S���^M��r4u�1v�w�َc ��o���&�bjK�kN%wT�iü�3e��4�D�+w{��	OZ5�q���g%���;݄3���[Eޏ�x���W�'x��>j�B��=:��I����{e��Ar`��A�D�w�w���s2���޿��{��X���D�VY�j0%S��mi�4��aC��[ws�ٶkװp� �0z���:{��+<�G�+�ŃtY�֊q1M��d����0�;k�oa�;�ó6d����$@r
��\�9J���u,��q��0dg�/�B_(�J�b�����~�b���ı���I�I$�T��\|��c�� ���p�P/�&�P SC��C("�ut(&`��68�%H��
(��UjF�X�c��#�e_�(�Jh�(*1EUX���\�"���E�
(,m��.(d`F!"�V@�"��%�����f�a�KJ)%˼�C	-("4U�7�F�.�6� ����L1��:�٤$�d$UBD3���/[�֟I[��~�H�G��O�.�C?��hRmi�<�m��Q�g�����r<���1�+�c�^�[�8R��hK���Wht#VYJ6�`
u�C�h�R��;^�oK��N��@�Hfdq��E���Ӑ��861'b{��`U3���X���b�"0�4�-N�	��>w�*(�%�S��k�\(_�<ճB���_�� A����tJD2�unM{�k�x�a5M�V�Ո+X��X��
���������"�QF0"��$RBE[A� �����f:Jŋ�	I�vkpRx!��3��23//I�H��a����T���&
���v��ln�-GE��CB�~PO��{'+���U&n�'s��Jڗ
;��b:x���Y e"W$��b�t-�}���L~X�͉���̿_��f��k�|Q((k�><{���j�j��.)h�R� �z�>�`'���!�xQ���ب���bDy�#���2b�4�0e�<(�B�6b� ��x]\�f]������ 0RY���-�8K�O{R�wL��3R�@�:x޼�'N��
����=�m$�`	(��\��q�1M"�i:.�7v�3ZiϚo�P� ��e�;�k>�X��H5/�0����X��'9�\�/�a��蔆��0M9�@� C��
 a�I�<X29:�ɑ��s�"Հ+�\���.R�L!�� I"k����Ӳ�h�H%�����3aw0�ɀ!�&NWA �����T�%��1� B�0�KD#XxN���(
d�@An����Lȃ��X�����C1ڟ��A�m̹���H�
	]�