BZh91AY&SY�!� �߀Py����������`�kC������� � 
 ����ɏ�pNCa5L$�L(b�`MS�1SM4􆞡�j�I�h4�R�2� �d � @=
S�)4�ژ� L  &�S'� ��      �Jz���=G�S��ɧ����$��j�=O#Ԁ�4 ���`QB�����	��,�
?���z�|��5�"(�U�@�zKԔ���A�E��A�d ��tQ�-���~<;��؃qb��Z8H��0�Ç��2[���d�|9�HÇÇ�X\��0�8s-�c�,��f f	�&ax9�f)�CX"�!���bd�9�a��jA��i���bf>�(����o�q���~la�̹��*��B�H�Qs�Y�%��c�7dc�J�
���!�r���7c�]�5�`O��<�]�!IE�xzJ�⌄���[�O�nj�B�=[���	��3]2���\�M�T�2�2�VQKdn�9j��;�#E� vYlbv�����J�m�ȋSq�H*�$���JD9��(y�(����8�.M��ء:�X���ẩ���r��*5���Nm��"|oa�^�I�F)��1Ld1c�`7-�f�n��CCp5;,꜕��9�
l���ae@ܕ6�+!���!S�
P��D�e��Q#n�8�U��w �@T+JܥU7c���ۯ�:�;خ���fb�=*��"h�-��h��BTh,�3~�UM�翺~����� ���w�9���M�#��ܨhHmM<��+B�J#�T�����qAH��yXi�#5l�/qŊ1�c�s:7$T����ԫ� ���1Cn�u)W��a���B��f�|%�BCko�^�}��s�G_�:�]S�&�ؕ�(4��R�n��Mm�W��R�j����ڢ���\)�=e'8NZ֒m��'Z%�/�_��w���3������Ǩ3++ꯙ.�z��������NP�H�]`�h��'��[*teQ�]W����b�/� g$��Qgw�`�2�+c&;V	A��c���l�Ë�܎G��0���YG�;�r
�-����~�Q���`�2�!�D����_N+h���� [�����Q)>툶��t�zX|��;�T,{����w�$���م��6PQ�ų2��z1���'$..4�c4o�H�q"��fN(٘���i���gHa��'�b��H�L �B5D��f�83<��ce\�>	�޵��y�2{vH��!$��p�pLɏ���ٵ��i��L,�\+%aҀ�$�P �2H��)Ao�,=��?/
|�!mX�B���[.(�t7a.p�/g����5�Ъ�f9�l��`0�� �l�;d����D�Z��<��oRi�db� ��P@F�7�92Z8m"ib2EB�d���d9�^Қ����Y�0���Xd	��ۘK7����{"H�����N_����K�QO�DWh�1G�)�+��!wO`����P&v6o�i�Ҁ�ͥ���>�H�X]K�噇����� ������U���}��%�ge��{��!�-BO{�r{Nm$�8@���7�mhq�VX�/gxEk0�H���bn�u���Ҽe{�5rڀn�Ge�H�1Q����K�	t�� aDȹ�3J m,��|wp��,R
�"c�����|N4������P���(ZC��T|ȶ��lp�Ch�,���%W!�5�o�}����0��g|!357�S %��C?����"l���{Ч��� �\�!���羯N���x����$ǷHh<�Ɨѣ����X�g�0Vh�S[��[��BI>Gg ���}� 2'��ˈ�2��H�^R��P��HH$���$�L�}F���3Qyf�/�#�f�~H3��^��OP���F���I0������縗�N�_G.zOd!�c�2Nx����T^=�c9zF�C���pOuY���C���dR�}V�WD�U��,�UW�a�s��Y d���2�!�JE���I�;T�����[v��{�QjȚc@�@�Ne��+y�L�1�yT݊0�z�-5���-~�@�~�Q���,��K�d�n�{�d��g���.L��!9��O��_��b�v-d��R�b��y�\�a�c�G��8Z6�=��焯�Hv����[f@mک��r9����Έ�}����Q��Y�C�N����5bn7欭��W��]eΊ`�Ѥߜ#��Fz�t3ޘ�G�ǃ�Î߼���pzSC��?���T����a7��m��ٳ���!g���4cE\�C���#<�u���8&��3	��s�t�4ڛ]b�Oo���1H[77\.M�M��Sp�ȥra�Xq.p�N�ʗy  IƟ�ƹ�v�����0��c޿+���H�.���I�{:&�X�a�#Ԓp�&���fU'��r#,�\q�J�^��/���y� C�P�q��*\�����`#��iO�gse[���Kz�˞f� �/���	��~v�t�[�v��j�#@��K	0v��|D5OAt��Ɵ6�����K H��c��#&?�ᗝN�}"|��g��En�T5f>ԓ����9̆X_\�w٘vr�qW�oC'���?I�1ђ�<���-�1�ͬ�tױ�=NpwN�Q�U@
� !K�aõ�����r�&
��r�Cݪ�! I�X%�(A�ԅ�UՃ{җ�v0�@/ �0h�X(��"1(�B41	 
�����"	prU� B*D�"�`�@`@?Иd"B�j�2�%(�\�' �0��D�1�6��k���/ ��}k�gJ`h6�<��;id@7ޝ�3_����O���oV������=���{k_/6ת_+d���t�"�͏wf]�ڏ���zZ��`lF���9�iSݓ��;�l��yr�S�_i1$A�;974A؇��R�@F�i��"J"�I'�k|����Ȗ�� �Pc�ڲ'�Ѐ�\�샔̉�����zUD)����G����#mQ��y,�o�:�ߛü�����Hq�c�8mt�f�|�h �Y���x	��h^4�u7�C't�Nq�`���I+���4�JJJ�����%��b�
J � ���)
J"���bb(����i�]� bH�Z
"(��"� ��8H�g��z1F9�cP��L�BV��6;�H;F�T
�L����Ĳ)�r�������F�;T.J+Τ}��b����J��<zHkl�����	H�K���p�9Sj>%6��˾c��}E 6I���j�IhYƊ����yp���������ڕߺr�"4H�7NF��O�%[6
i���h/&C,-p�	7:��Y�w��F���3W���y<���1%��6�p�2B+I(��&h\�:l6Ӷ���dn
8��Q�$( �>r��Er�$.�-�K�K��:P`��ar rL01y�w������TC~��;��DQ��Ӯ�=�_�u'e��`��̭,#x�R�\��t���@RI�64�]�pB���l����Ri�$�A�#G  B÷�P��߆P���|�C�ĻZ��]Q�I��0���Pq;=��9�ӂ���we3�$����`�����-)�m���r�!�8W#�kC3��5V���G3�ɬ0����-t�a���-���
�����z�H��~I��Ȝ�%��&X!h Bכ|�TԤx5�Z"���.�~�Kd|�S����C��>{
�a�7�+K��w$S�		�|`