BZh91AY&SY�Ʀo {_�py���������`�|��Op�PP�  �m�`�۴�%��)��Ѥ��<� ښ�� h ��@�*=OPi��  4   �&M4�dd�т0�F� JzET�Q�L�����0�CL##j0$�	z��4�224�h =&�D�i4�	��M�=2�� 4��SE�A�O��[���� �FW��l�]�BDU�P@�u!uI%�C#qEx�]b�@BT���k��a�]ϗ�t%O�{^���;�@�4�t�#N��it�:t�ջ�4������;x����\t�:t��4n�����Ϗ��������4�:wwwv����>>,�}��d9�ܚ}
���@�;��a��������&vDMD�y������B]�p�DaT��K�b���Y5_�:x�JPqV�Bj ��{4 �O�0��V�$f@jN��)(����(��V�eʪ�K�����S��2�fU܎I�L0�d���mbF�.�#�������4�y��>ӞQ�����3��N�d2[�����b��丈��sI������+-L��¥H,L�i�����ȡ��C�����.	�}8y�,�  9U��vE#���Ok���`��t�����ٙ��{��{�����wwv�����ܻ��̙�ݽ����˻����ݭ�2&`����۪h��$nc�l/HF=3��nm��x��6`	���[���� �B$8�K�~\.�	䢑��6�HvR��v�j�����tZ�ňBHZ3����xl������.Y1�á]��e�W_lqn��Էw :.���~#����5������&���x�X����a���v/]緜��Et�O�H٘�Ǿ����9�:��Tr��#������NIj��F��Xo�-��+:s3�bXְ�3�;A��>+V���86�9tȀ��0���N<��@�F��m�8�:����1�L�%�!��2�-!�b�Q�{|��6N�]�8� ��Y���܅�p��.�a�C!�"4��P��O��n���7�a�àz�ׯ:�x�,I��$ \� �u���������07�n�``�t��d3a�N2xl�?�I��uې$�Hm,��8M�2t���f���as�Q 8c��$�C�4t'pi(��B��H�搚3F����c��@�4߆b�jYi��sQ���ˊ���V�t��{������LȂ7��-A�N-ô(H�q�g=�݀�~���-8�5��	�0�9�w�D��������G���!Z}a��jذ��5�<@F��}����(�5�橁R��0�c�aY����!cM�!�"�mժ9�i�Z��M:o5�qM���a�jM�P:-���,� F��-��0cH��O$)��0���lvbZ�'ӌ=Q�&��DI�hQFC�h�����(��IP�a���6�qz�>s�L?�ك������؍?>87��*��u9� �MB!�]ҽ��õ�>:�*%z�]��3/Sl{(D�Г��}�y�B^���+Ѧ5��]^����8[���5�P�SV������4D��<`���xbA	%·!�9���SjKA/]!�+S���G����<%+xq	,Ƚ��.8��dG��Π� �0�r�l��U�7/�P���TZ�|����ҚˋQNv�z�i�^̙4�zdR�-�e��j(���g{�J�5��)M2�B��I�\X�4v�����Ua�>F��]o��0��,���鿇ma�2�dB	�$�o�Iy�~��������H�cad���_Y��Xk=�w����1�!^�\b���om�4�%/9�f[+x���|�+@�N���K\m�}`6�}5J�&�3
��>��o&�-���ˮj�3�UQG���=t�9ٳ��Oƌ�-˽;�ק����p΀�xr@��D�C��C��ǳ�N�w���VD�ؙ.��CK#	Ʉ�I	$X���������% ���.K��-yq`�	{Pw�]K��7{a6�IU%`�!��P�EQ�fH��ҩ��eAUT�eT��H�(�4���*���i��U�(�2B�E�P�@�S|�e�*B�%`��$R�me.��д-Qb 4#[(���)}��j�)b�R���W4�T[f�s������Bh���rHb,v��Np��O].�u�&�H�Ǆ�O�j�g�q	3��
��֟nu�q��,e1(���}�ⰰ��U�L�5۹�ԍh� ���4�Ћ��Mnt����A΂��0�H;c���q=�s�n1�Ҵ����0��ѥ�!����IН	��(�h,R[�:yl����6d�N�W]
l���MXgA��%��e_\���?�.��.RuةA ����Ym��&��.�nx�q���$-�
- Qj�j���ST�

 �� �R��;� H�
 ��e�*aP�R�.}=&v���!��f��f/���(�@�� �Qj)�"�)"��2�L�|6�1�4���8��L��c)q��Xq��W#���xS���3�⩌�����Rd�gAx�����GQǩH{���s�*��P7�E�		Y��k8�v�i{L�>注P9A����C���b�82<��Ӻ1f�lh�E�� �����4M��GL"蠼s'xd*�jbb^EvG��@A�`��0Ε��6c`��E�Q�p���g� ^8�����j�"���o@�
�F[�@�p	�D�K��"�s�]E� б^�Ǟ ��ù@���,����6F�?�?7�(s`�x{\�G��_	�T�2��ٱ>�E0F���1�YV]���	�����J ������&�9Z���aӭodH���T�Fk(�Q��!��D���ǁ���i,��H�ٷ˩37^J��P�|���h��RH�5��Q�WT�oo�=����C�;��@�9UAD
ZCٴ°lJ��̗�  ���*z��@�Ev���;L�����U*\�>�N�xj�*t��3������,��	�mu��rE8P��Ʀo