BZh91AY&SY�pB5 T=߀py����������`.�  p W����y2 �n}�5R�5�`T�غ�
s��U�uǏ<m��nN��k^;�)����m� �=�����
 � P   eS��Dj�����4#@L� h�IO��@42 ��� dO"�jz�A�A� h�4   J~�$�eH���      $��F�LЙ1'�Jy6�L��T�FPJh)MTz��  h    p�9Γ�E��ڪ".(Ѐ�n�"�YRQ�O�����1�3�"(�� F���z��J+�����!��b��C�~�g���������l�y�Ljl��_ϝ�,,c�g4�c���'ou3�s�鏏�4��x�j�Z�ӛ�fw��r�w(�O.y<���q�=o�֧nkW5*�v-��[q�$�JԒ<���_�f^I�Z^[��ʝ��m#��9��އe�v^J��&K����3����{��fw�w]�.voZ�7w5P�gd�g�Zs����L�7�V;s���l٣F�Bw\8�K,��"hDF������t�8t�9P�&�DuH��������Z%�"'�jr�6"Y���lDDDL0�@ �!�p�4#�������P�����Љ����8nW	��DCT��"hL2�GN�:$��b":�DDN��<Zٱ�NWIʆ�R�v�ʜ��e=������o�I7��5Pцk+�a.�DD��{^2��"&0�IIB"&Μ��Â"`���"tL�Xa��wX"&�X��4"#�N�X��v2%nv~14Ώ��������C�~��}��?R���9TpR�N��Ns9%�ƑRn�Q<j�3��ɘsp9�0�d>*�R4En�ֶ�ԑ��Ц��	�}��Kt덈��8n�V%ǫE�̺k����'���0yr�zg' �N,�z����Ӊ���N]d�=M�LdA�i�nуc���7bOn�5�"'a&�L��񱵕��n��os���bLh�*1D^��q�F�˸C�R�p�B� lX��Rw�։��=S�#i�M�4�Sq�X�!����ǽBNBpP�BR�H�f�$i`s+᩺�6��М8�ӓTPyZ�������ȇe�c@���<]��&�+M]eB6�ݕ�xq�t�E�	
���H�(��V��]��e��e6��7R�(]�6\�$��]�0���C��IX��$,n#��1�@�:�Ԭ�֦�t�ܘڳ5%��-��_���u^=�J�޼�}�<�#Z�!���?5g_�:���ħ��Yc��r�Nr�Y�o�ȻN�g��i16��K31�';�OC;G+�M�;^od�OBj�2U��_�ʩf��W|��N�V�5���$%���977�o9΄6߁@�T��̐yfI`@��&ƲԩZL�SLKH*]L�b&�����ݔ��śkn�k����c��� ���X]��h&ŗV���\S�,ի,�]�Z�HP#M�Mu���n0�uMk�&$��KB�F�j�8�	�.sd�U�TI�="g��a�9���s� �e�>��q�2o��p�y�ˇu�r4X��QΥ�/D�؂��:��g\�{*UTT��KF6f�F����kGZTt��B5ED7���֭5�h�*($R�$�*�$I�k�����e�Ћ`�/�f�@�L��-�!��+akף	��m�:Q�K�� S�5J��j�jhn#l��J�\l$cŻ8�C�H��"a���!�b����(�]a��f�Z/M&\lkv�����m[iX�d˫s�G9y��.��u�D�\�]n�q��˛[̋%�v�%i6��D�ܪGi5
��/���
�J��?X����W���3����W  G<�3����,w�)�����;B�0
( P@��@4( �J��1�0hBC@��44�ƘƆ�4Mi��D�E���O������zcb��ö�Gi�ٸu�-����V�hZҩZ�B֕J�Zh�^PD�ĉX�T�\#��V�f���:L���Kr�;I:m�v�a�p�h��l#�nm�m�v�í�7M���ô��6�;7�a�ةW�Z��ǂ�*cΥs�e�/E	�	S�L��3[ �|�� ��\� �$ FOG�=6�WҞ2�wڶ�@�s�T��KP��T���m�5��}�6LD`��:#ǁ�9�r��Nn7r���ֆ/���/��˶$$�$ɑ����:��%$U�+8�j�ãā�`�B��#���g�Ӄ(FY�����M��Q�5	B7`�] �� ��nb��M�����8к��#\�SR֕B���3�c@ ���0�;��9�L�ʦ\p_t��}4��s��x���xq7k34aalF�*�(|:�))�v�s3 }��B�C��_����0F;a�'�0�y$�ݺ>h6ĆYp��ʓG2�<������S���G���ApB->!��r|
lT�adq2iQ�}	�GG�;��<��Z9�����m rɱl�I*�v|p���T�����H�k�AÎ9�%��3P�!�tx##֐���CX:*řO�L�38�E�7p�nn�+�%+�"$Hm��)�P�1������	ćBa��d��1$V9N�|y瞹Q���O�;{���7�aG� �;�pc��a�?�/�;W�Y�����O����_&pL��\��1��1M�<m���9c�v��G�2�a	߇\��#��0,f9����>$��!L������3 ���<d�pEB5R ��f.�(�8.2c��F�(�8�h�D�aP��!gFz��_�8<'hq��`f=�x��k�;Rଗ�5�YU�_�ȧ,�1��@Q�^#�����Zn�pF-%̧�5�:�?�-G����
R�4C!	���.����b�x	�b�g
v�
�T^�k�2��C35_h��y�r�C�B��U����6�8�F`����A��e-���)�grݚ�4�GdG ��m�g��rLF�z(�qD�xxBR&�E�<�:d�D`���]��f�@3J3[h�ޛ��,�Ѫ#3��32���¢�-���Ř�2n{���m����[D̜V�"�Bď�-�mZ�Ulw��uvۜ�R'#4��-��-{h��a��f��lYC�.R*i,+��*��(�"H�(A���~��g�A    �ADA�e������
�e�op��D'�I�@��3��c��p@쾝f�8�<8C3f�����:������9�H�T+�Q�8<u�$����Pi��EF��?˦�nB�~@�=�+�� �50�`�C��iB`
]#��]Q�j,�pZ!���جS�,Pq���<���5��p���9c�@�D���30bn�f�5V��d9�3Q= �����&���>I���ۇő�-���xTɢ��l ��(hϛ8�7VF|	��[33��9��I�jy�!��� ެ �u����������qІ��af�
!�Ӆ�_�:�S���0ݝ��BC �ɝ<��J(b��Q��lc�K5X�13�&���u��,���aF�%ۡt�=F��Bo)}m�(�TN_-v�R���Ո�qo��:I#0���ʋ*3(�v���Q��]��|(��,5x,���xێI�������pPCxC�8�-d�<��P��zxD=�#�t�r��8m�6ft<R��@�RJF� �E`H���6bYCCJ|����$�܁�s���L-��qI_	f�>p�S�X�l��ɂL�=��C�1��(W�6��C=�
4ӧ��$�0d#��P�jf����� .Xxx�þG���G�����§�v�š�37�����<2H,HP�F�
2ӿb<c�a�ؓ`q!f���Dm��|��s�k���<i���9���҂�"t��l��c���C��Y��I�a�.�#����s�s��v�0h��9��"��8��031-�]ʁ���N(^XH��$��n�b�� �D��I�����/���bI��DaE�sDQ��u�������*M�'��	0�!1i�$2L�ũA�Qɞw���s4�l(�wK���ń%�Y�XJ �C��2;Um�l�<��!�	�\��gםڿ �� ��(p���v� ��b����
.\�q!A��M��T�Cq��M���Pf�1�c� ��z���}�i�k�.����.�1�4�fdy�dcq���sL)qm�X�I%�侈��Y2f���3I	"3$�?-�u�Ĳ`fc���$b�0� �b�<�A0 ḷfw&8�D�X�H!���	0�C�2�a
A�<� <T"�,D�8I����0N#�لG\qA0C�2��K��ا"�wKn��Ft�MGK�8@�0���31R�Z.J4��2��G �331�1�;z�5�0]?>eX��#��'�*A�@��G 8��r���-����y�J�|��4&t�ι�,]t&yX�������,I��i��z5�m�ڠ�z�@�}�쏷�^���+"��Q���~���>���1��x<[6`��w��M�� �!lƛ`�zp�T -���t;��/�G�i�aI7�uO
�lp��]N�T:2,��.�ԑ؄"B���"�ho�G������f�fh"�p�]����1F���>�p�9�t��qd�df>Sbh����j��4�֮(}�,}�pq�7�t��j,�n�Z��3el�ՖtC�<r��� ����=9�)��!����y���Ց�C�tis��f�ҬRh�I���QP��@��DY�9��G�:�#M �;0���^���������۟3<s���mkQ�@�-��UC�hu���ГW����=�u���6ճ
su�ЁБ��eO̗���}������ga�l��M�k�h�n��I#	uҠ`�1�,�F$�
���Ckh�cY�f���v`@�]�	5���`%�iDPf!�4�B\�� ����B �AC�(��<0�$�ã�^4r�G,]$|3�*JΜ�L�Ƣ�Yps�զ:�4�-#�31�8��;/�X��Fh��k��A��%��*���P�V.刁�t��d�e�I5ӶhX��0�;�ɨÁ� G&�F�sM�eÆ���4D8�B89�X5bD����fB-��Ӳ9Fқ�|��)z���z1
�����f`(�v͂f�ü&`��8w�G	B��\��+�t9�,�kvg�����1D�� ���D�Musu��s;�LJŊ�**+;��f%��Q�R��n��濊�dS�8���9��o3t�ϰ7�\ ���׉��d�_}~$���k8FIFˆc�n[q����0��y��dV�1�FS)L�0�i*{�^�;��(���ن�')��'N�� �K�w4��,ÿ��s�a�Ê-� ���H=�&���'H��t�Hk�-�i�7���1uh�m�e��✥:}qX�^��#��"E���h�8X�-�"��V�����3e��\�����g�PJ�39RW[��A��j�.�=��(W�XJD� 
zv�ݙ��m��֫z��W���Fљ�E�EW�G��ڵd喜��0���I���>�E9���)�v��уȆ	���X!a����)���v2��@"M���"���]\]tnθ$�K.R)RJk�������0�39�����L�AQΌ.D_���9��,��>���3��4��8��L�L�P�+�*.@f8!yK>tI೼�$N�!� ��sx�a/b�@�h�z�+�E�H���II��V�U��EH����b����ĄRB��c$r
+�3��5��9ä���pAh�	���ν���?�U[�=DS��N�w�l�9e�Y�oG��Ȑ"Y6=�N"$�4E
��t�=@D �����1asz,CԐ#	�	���6��J�(���� ���s\8�$�'�%���Wy��6' @�	� �[j[��JL�%T�|�'����H�:$茂Ԣ5�,Q�ȍ@I,ִm����sh�jhr yOo�|�tA���}8.��1�:�B�E2�2������88�D.Z6�9I���z����PeEg��fRYe<�ŕ%!HA�D��e 9��g8�Y�D�ޞf�P�	�Xs}қɹOX-�)�1�t^ΡdA�EP��"�fb�s$c+�ZE�(�k��δ��Ɠ�H�MJ/�\�#S4� H�i $�Pc$ÐK��M'e(Å�Q����
88���%���9��{X"��#��|n�0��s}�ܙ�N���x �`u���\�!#-ߢ4�"CY��b���J��` ,��d���C�=h��� X�*��/ǖY�a�󾤵�)٥�D�^ ��ڃ(Zڬ�b�E�%�	�P@"��*��K��[Z�/P��������L���R�B��d�B�dDUҊcR��K�J� �)�Ű	"�As
W"�Щ�X��"�pX�(�@G�
"�e\̱U���ʒ��Q�:l�V0B�l���d��4�H��b+h�dKƠE�4.��8���z\���AH��y�R�H"���m��[j���I��g����D}��uA>@�AP����w��?$ʐ�r� �������AP�P����a~p���*����p. &ώ[���*@����=�#�AA�AAAYAAffW��'�><{�?G��!������ys.�OC��D��X�&F�+<�ň����}^Ng?�������9
 ��N������C�C�)�!�T�<�?�4�O��y��x^��2b�rF�#���>��l D��(*u}�C��D���S�|^@@������{�got����1��<vW/�w��b����#3O_�#�f��u��[2ƴ~��E|&�OY�&w���)$���7�8���0Y��JE�%(�@H
AH�� �U�D"�"Ҩ �$D���*����fd*�J���V�<�#1�fE�va� �lL0@��6��ƈ��hX�TA*ظ�obf8��5}��!=}UĄ���b%ߖe���؅����̺{y0" Y�A�K'K���;r�3>��1ğU���K!��`u�	���0���x������8[�>�ۖ�����#�6��UDAR��������!��%[���6l5�C�wӠ����B�>������y��a�"�ug�!tȦ#�Y1�*��8p��FAF�d��E�b�P�Qgɇ0X[��Q�G� Qj��DI�

��Iي�4K�J�����`�lR�����LE B�!���'ר��q�f� �!�����zu���̀������3�8y_}ބ�;�������$CɊ%'�����}! B��5�[�<��$/(/�8�� �>��T���?��ga�<>L7�ބ7��i(�HQ���/�q��K	R��à�ۛ>�щ���g��L�����8nL_�2S6Γ @��9ŭ!y<	�%	m���Mٺ��:��M�D,d[J,	I���7� s�oUF8�K�P߇B}��m����{����y�U@^VO�����݇4����9�G���C��+ɌP�6��q������)�s��