BZh91AY&SY�{� �߀Px��g������`~�!��@   ����Z�K�R`�)�Q�h�� F�!� d)ECM�m@�#M2Mhɉ�	���0 �`�0�&�B&F�z��4d=#@ A�~��A�i�?E�y���#I�z2�d� $�h�?T�Ȟ��� 4 
�(�5Tf@P.�#H 2{��qL`,X�	)����Z'�`tHMXN�2��CZ(l-��@����>�g�}����V_ۙ�����������iiӤF��t�-#N�:wPߺ��.#�t�<G#L�:F�2[Hӥ���ݑ�������fffffffffff}:3�mxD2����>�,��+���?_�
p�F�*Z&>�0�Q��*�=^[�"&�Q�\h��.
w"�!%3m�������.���*��l���P2�a�;�i�x���ə��|�t \	�)bi��(C�xh�" ]e]�t��ymVUcEUשۢ���ǳ�sNiǇ���	}��C�][p��	�q���5�Q���j9iW�W�E�x��T�̻n�\��MM�wHmc��}U�툐em���$JY�4a���E��V��dc������˻�ۺ���������ݻ����8ŝ�7S��
��I�bCN���cyY�O�5�OB����	��υ-���2��e��U�Qk)�u��\�6�N\�d����5��_��~���"&O����稘�B�3�a�+�5�<a�d-���$��U�G@�&;).�����֋al>|��I'l��N͆�%���ogY�gl �b�Ѹ����	4����ٷ�n)�3�p������وl�.�C�l��!D�
�[�ԅ&ȏ}�± �7H7)p�pȋ v�2�Iayn��5�����C-A�1�`0�3-/"�"��߼���	�����ǫ�d�f�Q~L�1ʢ�!�A-N�P�eБ�vj�k�d����,y�I���:0���L6EiVFgM��a��������E̈�1�A�kޝ,-Y� ��<�́3U�@���Ϛo������Y��e�q�u�I�_0|�fލe&7k�£3�Ue�XN��9��iu|u�!���T�`t��\��~+�%�%]�bA$��AD�0��/�P�°g��\�s�C�2U��O��/?c��{��lӂ��>#g�q7��5k�����%�����j}����������u�%^
��'�ܟM�5:F�"h��SP�R��w���L��^	�ǃ��^�ʈm'o`xy:
��$�o{|��;�.U�!9@�:vA�;w;0����->�92���A���WM>fs��8�q�q�&g�K�SOp�M���8y`XkɎ��� P7���yx`����>񞉈x�*��^mT�HFg�,f�Oz�O���[�8�\S�Ql.*ߗ�=�b��g졞��@8>y�2^�Ư�63H�?}Xs柳����@�bP��wr�x$��'ӓ+����.���=�y�~��Sa��.^����8��w���}<�f�mü6�D�����> $잮�-c�zÈ.��|7���:9M��dD��7���z�d5���2\���@ve���F�\��)�p2��-���ȣ�P�B��Ί���Q�F��㶛�aPۧ�x��Q�ڪ���! П'�������s@z���fh�j$
,�T,T�	\� ���h܉9��

��܍�1M�J��kZ��@�PX*"��V(��R����DUPX��c*,$���
@ђ���]�	y�*Ii�,�ip�b�	ma*̰�K+��YD��'6f̝��4C��Mh(I�}�s ��$��H��i�Ջ�g��Yb�YW�}q����?�_��q+���XX��a�j��U��0��*Aƹ핪�+c+�Q�Ί�ȈLjJ���5�)�i@<HH�!��D$Hl�M���-����!��G`K�T��o�� �d��S�)��ALw��V	������RԴ��w!S�ﯠXŒ�+���g���D;�rD��Y�ϋ�
�#�i�8VWt��tKY|ވn���|���U�,QDPEQb��T��`*��X����"(�"����)�1&�a τ��^��M�3(�'�p�8COI����d5��*��H�QJȌ"2 	-�3��u11��> �1Z�5�
����ޒ� 1ݚQ9�����S���T���{ǻ7ޛ�6'�����q�Cw*<��&��X�}�I&Êwk�Oa�� E5郾 t�x���6[
i)�>=䁊�" a�:1� 03���!��h�t'�iv7��Q��,'K 0+��n��g-�:���@h�7ww��80�مJ�B ���6��S�����8%����b(���3�k�;�(F��5��'G��� BP��9����!��O�z>�uT�2v��ў#f(z�>:�&��񨸈�8R/�)�9�Ug5�
7/5/&!*���X��t!ٹ�b�!M�,���t��N\��"rp��zM��t�k
�r@��ɏ���ju�%	m2�s��:k�i.tn.,Uh����.��A]y�������a�X�u&r#�U���f@���[<yP����%�N��9ԇ�^V��5[%��rE8P��{�