BZh91AY&SY�� ߀Px��o������P��2*Y�j�56JzjQ�SC@�C!��!�	���dɓ#	�i�F& �"d�$�4�U4h�z�4(����&L�20�&�db``$'�6��i�S�4���� ѐ4ڙ 9I +!+���{�z�M�)d0��BZ�����bָ�X}��	ֹ���V\J$��h1K��l���z�;yc}�K�	֛:��K����Af2:9�ӘQ8����w�������ع\�ï~�e�����;%�Hw3��lG<2�#~h��	�a0�(�06��ٝ��Zl�N�en,b8��Hs�A���mJ��,���4�S�33��31v)fwp==��8�،�kM7fv��Ӳ��g���N�3��|N�ޚ��il�6۩�u��s��:��l��j��M����m�	�� /<?
�Z`���x�ӰZ���kgy%�<q��C��������d�GmB
a3.5[�C)؋W�~W)4�Ӻ��(��T}����o�܋����*����v�ne�����,O&�:����?DW:z�Nw���R�S�ڛu;>�N�	WH�(U��&a~S�������j�*�yEv��H,5.���\�����/sd��+�:[d��v�S5{�sy\Gf���V�@��Qd�-Y��22���iy^u�(fV	�`ӥ+"���mT5Ȧ����WY
�.{/=�G�pृr���9=lEC�������L{�-d����u�+sセ�a*^<�F�"*d�#~$0���Ĥ}�	V¥��K�4�d'������#|����&F!�ӗ�A{��\����P���04Pȼ��ar�\�e�U�m��'��&[v�"���%#r�nB��&�a+�J-���旚U:�Ɔ��h�ՙk�!��0�q�Z q��p�8dxyy�r����g>/�ͤ���X@-)/l\|��T�P,}}JC�����&������M�H��,&6<꙳��9*Yq�����$���K������p[<�$�p�K=�{��/���7`����{0�/g�W��d/�HK#z��g�Y4,��WA48�h��dwT�19�s�]��pY�D��w$S�	H+�P