BZh91AY&SY���y &_�Px��g������`?=��<wk�|g� �}   �,�Up-B%
�O@�ڠa3P hh@4h�@��=&&��h�2 	���UT�0!�   &�`I�P�J   =    D��2Fi0MT� 4�h PD#@�I�f��ze=M42 ɣL�!=�* �DTq@� �B3����ax�����P T���e*����bBr�x\e�,$�M���ˋ��{v�ԛ�ǒ�� �СP�m�k�����������]Mu�ݳS]MMu5�����Mu�v�h�5�5�mֳS]�9MMMK� �I�[�������뮺���ѩ�������G�'�����p����� i>���x�]����ZA��LHPL�	���2Z�$،�Ll1U3w8�JYp�7R-�rM���zS�D�m���U�uz�E���X��Ei\���33" `4� ,�.:�5��䕻Rl�[o6v&���i�x��N�C�q&�`FJ�)��Y��w�Ge�-T���;�AHڐU�"�tUG�]�� t��[(�������Q�l-U���RK��#��ٌ�_��׀t�:r�PP0C{nm��E@�6͙Ġ$	ȞM��\�*�I�[<�(o.�Ұ�8�[������,�Q�����j�����J\ʹ)������%\a�Z^�����s��DSBm�\�*��B*��9�2�DW}R'U��������H���R��`�Z���X�ƪ T�,*`(7"ϩUmJTL6Ssv.<��k�k�����1vq�����ت����痕:����4	�xo���@*Ny��Qcb�mzD'?�%�a��1H�"%�B4�A;�]?�]ԉF"?w���ǪԨ�{�O,�
���������	���O@f����_j[�sG9���3�M�9oj�X�tx6R`�H�C`>D?\]m�������*��^�v`��Oe}`�G+����|����$�%\���o�Y��T���91�j�-�R`�V/�7���p��%*�B���F����!��C9YC�Xx���!���$��@�Z`�0�&�`aG'�r��%0IɓTl�D���` ��2��a�M�-w�4J�٧�:�;����0�G��Ÿ������	̂J�(E;���z�� �@�mC���Ai.Y�,�	�.<����D0�ʖr��՚�M�@��nn�ȉ9�G u��^��X��BX1�O�:@���«W��1Ő�G=�(�%�`T�
(�P��si,:���7�4���E���E�%�H�č�"������ϖ*ׇ�s�C��\��&@�0G�#�<C�C�v�H
�d�H˒kcLY������R��:(��E�i��I�w��3��ц�]�f��l��@�}�����`4��T�/g��e��vN�{r'�iz0x��=؈ �H�{a���y%s\�Μ��.-��|��=��t���2�v����j�<jnC *nj�<��x8��e9֯;�0A��H0F���_�7�&�
1
��ZԳ�WqcU��l:᜷�0�LQ�eyCw��t�j��2!�#e���QL��X0�;�Go8��+� � �S���󓧝Y,*�I���DE��aJI�X�(K�� �ޗ;����z3��=?��\�yayAa5�p�}  {���c����>=��&�}:\ne�e�[�bhT��z<D�<���A7�D���\c�>��/F���Ϫ�{��݂!v6�e�\Lz�6x��j2,y�b����n6��.c���B����1I���9BI�͑f.�z��Gcd&%�E��U@�]G�1�Ƴ���q�/hW�A�FTF+����(�'f�͉��Bj7T���a��	h���Kf�`%\�������/��u�r�;�[�����8L��<�4��ڎy��.$�\��"Ƕ�k��w�I8��:a�[1�0TM�n���7�DC�,�~��t��> ���*���Ń�U�-ܤ����W����c2���M���}�$]Sz���n=�e܏�����狺�;��Cӱ�5�����
�*'l �g��]��{������C��X�	�ȶ�!�!���0�r����~��2
i�k���A�H7�"�K��̿MhfSm<�Ww<�Z��W��� 2�G?�0+���w�e/F��[��7�կ�ݎ����q����0��^��5"s���V�U��Rd�x��N�6�b��U$L�i�2��0�M<	�.����Dy�?1�]y���kPf~�4�����I��\����y��ćx��o�9�������<M�m�_m�{h��|�]'g���24Ӗ^�a^6������^Q/�*0����I$�%�Q��a~���� C��9��N%����]Us���[)(h��ĕe"!�	P `2�1
)D$�2*5)�6h0J$�@đ@Fd���d#l)���( bQ`cI�y$���Ka���J�L�$�s���	�I�L��N�8悄�#��y�EY�4�΍v��g��U<�)��NyH��~i�~���Ǫ�.�6��Է�PP�	�8�� ��s�P�]+�0�vt���=钺7%�����y�D�vET�Ié��v����9rF��w�>51i�d4�*���_'W�U> r�W����#ZF�Z{"<P�֞�ě�q)����hR��-L��<�j�9�!q�p�C�*"u��c[o�	x����l<�v��|w�3h`�hH[ �1`�D��,YPD�V1�1�b"�����(
���" �[�F,���`#DXv
T��P�1b�B�B��1��k��B����k&A�0�!������DM��A(Z�ZP(�"��Ȭ���Ac�Vf&���V��`�I�Gs�A�\KB�|20�?D���J��S#�����);�Y�`<�͗�8�lOOA|^��l������
\��*mv��jM�)��-Ӄ�2��P6j���AC]���3٬�.��T|<�2A�h���9�P=7�P`�t�t��B/Ei�5
	��31"<Ł�D�p��B�K���_TPP�:�Cp��Ӽ.���M�ST�D�Zn�%�a�²�����)h9e��Z�!C��M��&��U���n�1p"���:��Cם��u�"tgL�����.x�｝V(t�9���su㌺ �<Ȝ�0?�z�P7�n
"`}��y�V�3�Rx��;L^�ő!���jP�B�eJ2��)��2�bk�k��d&���`�����L��%�����`z%J����5��Q���A��l�4�����K��"Q���p�
s+��ɐ]��}�'ɇ"ǜm̚�:����f$Q.�hT��t��rȕ5�l����eHrk����1C]�.��]��BB�#u�