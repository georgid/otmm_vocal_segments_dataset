BZh91AY&SYV0`� �߀Px���������`�z��;�
�   ;'X��� �ML�ёL	�24њ��h���$� ��  22�O�RC ɣL���@� ��
� h  � @���&L�20�&�db``$BM&ɉ���dcP��2i�#F�yOI����iUP�T\¨Ќ�=�pY��BIG��O�ݣU$��� P��b=q��AƊD��,�K�������n�       NF�Ň�a�f͛�x��cs9�٘�s7h]�7j�6E�������]������0�,8p��-"�Y�C��������gFAo��B �~��� ��c���I�<$���Ikv�g54 <�,�a�rf�饡��]"�p�C����E��y�A؇m�g��<��l��Ru#��MѧÍ6� �,qx�e,\jwW��v�[��A��+-���9��_D�j���(��3	�ٗ.�fHa�N��}y��;��t�Sȕ�D��fR��ZT��K-���(@�>R1p�wW'w˵Y/2�nL�$�������T����j�cE��x�'���V��	"��.�R��w����7I�^9�͒�7��˶��YO3��7uUUY�Uwww����UUUY��D�LDXi��r�*�\q�3������`\��7������O=��!!_N^��^��9�y�B���Ń�Za.Ki������R�
����t玝H�&f�C��y�r�˗��n]�$��>�j��j� )�Pɬ��,8��|Cק��4ϣy���sE7H�oK<�q�a&�w�
�
Ru��C��z�zi�zWi<V�3�9��0i�Ӗt`���B��*<Ɛ��ƃ^�k	�����]g#d+�\P!����M\�����oV<�q� I�D��(�Ꭸ�h��q<
M��:�9/�yg���8<��a�I$���Ht�ZHx�6X0܆ xzc�ӊ�C�v�.CD��c��Wp Zjo{7pz��"[�! �!_F;ԠAQ<� l$𗽝"O0Φ�@��A�q2Q�'-f�U����M�T/`v�<�;1����cD6�vy,)D�p���d�"���4���w�t���J��=y�tk��ͧX�:�zG�ɒ�F����5�/l	�e��W�R�oKF�cH���ga�/���$�8-ql.D��H �S���*<�t���)[c�r�0C�V��lZf����tGs#V ;������������X� 7��~��\��7<�|��3e�V-8��|I�� ��y��P�x!��4*&�i��6��UF�/� u�)�r<���˰zO�q�����Ԁ�P%��3��w21Ui9r \��߀�E�l�"a����L=MԻ7�[U��q���P���`�Ʋ�0�U`��ȓeA�jc��8<��W���-�f�TI`�ÄK(e-zSS�=�g$���wJ�� Fxs������*�t!�@���ձ�Ǘ�%�X�"c7o��sult ]�f�<��ۇh9n��b��s��:���+��4;u;k� ��|�,2K{y��eN��q��@e#v��Q�-�F=!����^`���]�M��8�w;�&�]��[�֡��h�;��vc*�j������m�Ծ(C6��MWi�DK���4����"�&��}��� ������I�b=΀��u��|t�:���z�}�`s�$n��P��4�k�0���
f#\���43�Q�����w��0 ��#��j�9��XQ�N�mٕC�����e�RƲ�%�	��*#s_U��ަ~�ѴY�6��1���&m�݉�����.emuoz6w�Gz�LŊ�E^�HF����S�h�9����d�$�I$X��ջ�=�=t�����A|X����P���3wR�d�4�T���J���Q�cp	$"�F[	 ���haH@���A���-�%U�4[T(�&��bDƨ��Z@��e�-R��dM���-q(�n�Z[�v�nɑ�X�`م5R����Օ�7D*�	�PP=�p� ���&�T��x���"2��$�2
1}�ǋW|:�^b�awFU^�X{߲?���K��س����,�71��2���LM�^9+���d�'�仩�$z4ù��"g�����{�N~����X���[��}��F��|iV��
��-�����ܩ�Nd�Px5��a�L�����/N?�|��g�N)�-=1�Nͺ�A�-I]�9&t�M�?W6�H\P�m�J@�<���c�;#���c��nv;' �ڪ��PQTZEF�R�TPDiAj�JQDE�KB%(
�\� uD��f<R��Dދ���2|I�y&�}�cI���S� X�TR�  ,�ȨKt��m���9�B���u�9N�#��Rd�Ð(v�1���Z??6&�l*;JM�,�09��'r4kN6��G�H3j�ל�I���ÌLv�flM(��\��s��ԀB��.H��5�;��w�k2���>�d�4�JE�̊��} �9'9����y(�s��8AB���H�dx��\�V�0��2ƞ:�<��s�g�W�i����E4I �Ӏd�q�~V�f��y�����}g�4`B��ѹ�Ρ6�;A���ݫ)��"��wL�vu�����eѝB����K�W?;<�f(y�9H�M�O8�.�<��IOX�"��w� �߶ǰ��Ey�DkxtEqJI�D93�9�'h$��{������I���Q��'Q݃��2o�`��~����Y��L����U
�q�:��k2��0嚚`��b��+��7fdG�C�@A>�7�:�ړ1� ��79��q��:ײ�rhi#d9�J�-�w��:�S�X0� �����H�

��