BZh91AY&SY�,w?�Q߀pp���g� ����at   �I ��  t   �RPF� ���� w|    �"        
 )@U�R�DP�*(�QT�$�I)B�*D��R K�        @ ""��  �p�g�X�r��-Je�/��VmzԽ����&�g���@rn��ӛ8   ���� ��� �@ 'g@݀ dt wD0 @ � .� GA@ ) !PP�
�� �@�{q󪼽w�T��]U�r�j��A n�X����}��_W�n�ky��}�P�ﾓqw�{kϽ�_ �}�W�|[�W��������۶ד�Yr��ksjv}�(��-ź��e��嗷��ռ�� DH   �� yU�y}/��v�uw����z���+w��%�Z�-9i��{�t���*t������k� �﻾��|ڥ�|EsҬ_}�iqjU}��m�>�(�*�{��Ꜳ���z综��� �|� �� 
 Yh��!b��+�Y�8������[�G�S�qo^כv�n���k�,�n�� y�,���^�y|˛R�r}yWޕ
�=�,g_T���.O\��L��z )sʜ���_}�}}w�:�{��[��  ��  �{�T�������{���;���/_'��|@�_q��[�w׫ͧ�'�Jz�z���,��_]>Mx  �u�w�^[�+���m�ź���m��z_6�wS�{�P]��ˋ�f���z���/x�+�          ?P��eR�� 4�F���h�P&ʥQ@ �  � <z�Uқԡ��  � � =��$�TԌ   &�hD�
��P 4   h $"2J��L��4�6��ɵ14�6��|	���?��o���:=�W+�9�_?�"  p.��� Z�� ?�PP ?��QA ,������ Ђ  G�J�I'�KP "��O�Ĳ*��������� j
����p �����A|���U�_���v"�`����(��+���+آ���
��+���+�
��+ب���آ����"�������؂��+�"���v� ��+آ��+آ���ت���ؠb����(��+�
��+�(��+ب����*���؊���؂���� `��؂��+؂���؊����
�� v �*v�`=��#؏b=��+�`=��	؏`���؏`=��)�`=��؏`=���`���؏`����/b���#؏`����`=��؏`=��؏b��v#؏b=��#؏b=��#؏b=��#�`=��v�`=��#؏b=��#ا`���#�b=�v#�`=��؏`=���/`=���@=� {W؊���(��}� v*�`�*��_��#�_��8�_8>I$�������k������S|c��8z{�۞� +��6������=���}]��ZoR�1j��)��BB�G�kZ�M$.4j�6HBc"z[r���t��HK����M�~���[ӻ�=�D�.�Y�N��]�Z�^WM�r5ux{�U�kF��<��֨סg�F�^ᆟ
�w�箧��?Z��u]�]C�T�>ӪUƛ��I���B��y^��߸쇵���QMͥ�A�u�>:�T��^甫Y{,�%�S�l�=2TcDi��h�Aq�%^��kz<<��Kp��竏U\[�%ssO����O�sφ�E��v���һ�;%�^+ej�JB�rƥn\)��*���
�(�5�HTKl�.��aQTF��h�K,�d�D
�$�%�ʫ.MƂIT�d�P�,���
�"�j�@<*���[�*R�P�)$*�<ۨQ�9
l3&���Y�������o�������'cG豅kk
�F��Z˼t7)��'ُ��p�Î�Cw��*�Y�40%�$A2����l.�aw�R���P�*�³~�5=2�kǛ8Uˆ���/<Ѣ��w9,�͐��|�HI)�.@�wK�S~xV��W���ܳ��9ʪ�׫�#�z߁�Ӽ�EF��R|�5)7���Hl
�IT�a��x��[�B��e��)��9`Tm�מ�<@Ǟ�!,�n�����A��0��<%��
�6֭�^�*�����Om��	r�1��F��XB��ۑ*���:�If����/F�Q�4m���ж����T�*�J1(�:|��Q~GN6��@5*c�%�T6�!Pm��DK��5!R�5HTʉIW�&z�ߧ��/�rnY�	�W�y��p��������uJ��8�+k�Nj���Ux�6[q�ʕ�Q���kW�O|���_�w���V��*R�8��ȔY�M�$e��F��ѩn:rR
����ٙ�y��6Lַxh!�|Z��1Ѳ���*%�f��-D*�Az7�a��fA@����J�zw�����7����B�:S��;�nA$Jl�5�R���{7~{�+�M�֪��[A{cl
�*��%@�� g�~�UM6a�[+{�Q$
�F�2��%�$
�],k�̳~V�7
�B�4�Q�� ��^V�J��$/\6�<,�&��W�h�7�����A$���n�F�%�Ŷ�j8�p�1�Ŧ��q�&K12���%\�%�Xt�h*���]5�����)l���,��j8O"T��l�t�yz�N����xOy���ԩ5��L��12R@�z�e���5����a!Q�X]/���QAw�l�� ���4Ӓ	 `�$�k���SG��̚�h��M�����)$j�P��#KP��~Ԥ�.��l�yLԭy{^��둫#���>�Ph��{�����i�7����Q�*^f��ɭ���������(�5����5�fY�L��7���5G�Y������y
oA�fHB�a�f���\
�Dj82�i.���E��P�I�B�
��5��%�ލ �&��7.7�]gu{�o�5��>n�q���k*�7
.�٪ZjSf5f(��f���K2ku�5P�iȴ]�,���ק��ֆ�.4\�]B�p,�%�
 T1�Qh���x�Qn:3a�ւ����F�̠���!V����᡹R-@�5�M�H7��a��ӷ�#��F�tdt������ہQ�`��*����,a	#J[.!��=�.�Ʀ�]�����Y�A$E����\ɷ�!����q��#KPm��
�H$��<��nq*��+ӛ��9
-3
@�˂Hx�U	)
��A�J$*4��R�	#T��A$�B��z�4i��R@�UBID�蹅��'�K.���J�
�j	 ����J�Qi�$��D*�TCUBBB�� X�ŅP��H$�H�JnbXl��O<��<2Qa�M�kW�I���5�Sra�t��%�MY�,���IxzxF�	0��Y�Y!.-
�%�CAP5��Q��uD�j�l�Z�������H$�T�$��#R���*%�Tam�-����ZUԄ��U	�Pj	%!Q�[aFPK�)B�*]�^dJ#PI�I���j-5
�V�om^k�2��MFܕ�i��*�YZ��Q2%�fK5������ޡ����$��+!�/B�2
 �%�\
��/p{w^Ц�����V�7T��=�Bn[��^r�Xa�fxQ�d��A�j�V&��J�D�xi�a�Xaq��r�j�*uE7H�&���#C+KM��C��j��^�q����9^�o�v���b� �4j=BD�Q�i�O4¬�Y�\}�o��Į�����o�5KN�*�S�w۔��x��R*�7R
�*��w+w���(�5�l�SA=.�n�Ʃ��efku�_V�W��iͱ�` S~T���⛞Tr�*u]����{��7�����>Gl
��s ����拯%�*4B0������W5�f���K�<��@/E�+݆y��B�Q$�5)��V�D�!��HITP�$�T��e�'�[]�%�J�*F�����޹�k[��_�'J��fB�	�y��n~�u����y�{8�T���*�5*���Z�dA��ND�����Qj9���m��t��2�]����T󆪶l��U�Hr���9�	�ʯل7�<Ԣ�B[�\
��tbH��ӑ/F�k+U&D�r_���uk�����|5�&�f7�Y���m�R�8M���Qj��������h�*�����a�U�P!t]�^ʬ�5\�������5�@�� H�"+���&�D$n��J2ay��r�i4k��4�d��NB��B�灪�L+3M]f�Q�4B��!xj\��	�(����;�3{�9S��(�M�6U��T�U$ksI����\M��T
�H>���p*l*	���\��	�B0�n��� �"`J��yE�&���dq0��>�=�7�u��ՙ~ƨ+�w^L�%�,�����	 a��/�A2) ��{�I�A$A$RD2��i��J�D�@��d��*I&��('��پ���$Y���6��Ȍ"�>�ع�z��SXy����Ha$F���ڨ����f4���Y7 �Q�[��
�F���q������o�礻=w&���W����j�JF���<3z�|̫ԣu����L�޽�����y�2l��}%Z�Ti�t�T�8G�����L�.q#*p�����%0�Qp*�RF��d֡!�q����Ee[)�RL.�t�ʧ%��~U��Z�vg�����Z��W(�E�����ؽ~��63�x�}���C������7�J�7��m$��\mj4�F�]��+*5�����	 �TA$B�!��B	!Id���}P��7h*4�L(aT$�B	!R4��Y�2%^9l.!U�TZj��h*	$�H$�E@���ˑ�R�B��	 �	(I��4A$J!��Ja#TTZ���A$jME�TJ#PI�I�I �(��ĩ�*��$���%B�\���T�h)�@F�Urs~UuݧTcva�%y��D5{�jp���*T-ݙ�@�L۶/�^GL
�M�vՁED���A��E���Vk[5�roe���B��QDZ�%���*-B��S T�ܗ)#���0�̳xԙ�F�Ե��nB�Sm�ɬf�+e9TYU��Q�āP,j-���%B�ZT
*%B�[�/F^{���'�f��r��L�+aAe��Ori􌺣�3^{�e�<9
�2RD�K$*a!UDo�VJB�n%�^5W��	���}͖n�~zQ=�>�.�'��Y���I2��6�
fk!A��Mj�a�w��*�y4h���zk�$�2�&1�{w�]Y͕��#�͚��;40���W�kz��s��}��B����~���)����+���{ä�jn(�b���ٌJk�׫3lY�W�Q�ȵk�Lv��vB���EU�D�5��6.^^��G��`v�����r�IJ4���{����߻��k�������O���G�����;��ǿO�             ��                 ��  [@                 ��   �     8    >�         �    h                              ��                                                               ��Ţ��8       -� �vZ       m�m�� Φ��b޻kn$�5����m�m����-6   
��  �Bi@Z�Z;m& �$t�826ȳf���&I�Pl�l m�.��AÎ,q�$ � Hl�� �v��`t�km� ٶ-I�B;^�@	;%�Qm-�   I *m��!-R��U*�US� �hٲځt�6��  �ȡ�`*U�[���T k[@&�2m��끶��Ht�oV�v   $� x�Tӣ���pdpZv��]Tm��K����+xsZ˸ ��vj���R�U,�PT�R�@��c!m��     ���ք��m�m�6�:B�8    ݶӠ��nm�e���           �;��@
P`8 p (0 8��  �J  d ��   ����  �J  d ��|�� �p �@
P`8 p��        � (0 8��  �J  d �� 2 R���� )@A�����p            �  >�      m� 2 R���� )@A����� �p �@
�툓�p         R���� )@A����� �p �@   8�    �h  �aJ@           H           ��        �>               H                                  ��                                                     p       l     �  ��& 	�-��YZ�5зL+�Vʲ��J�A�-]U �\ [E�   ��춀    >m[|S[�    �.��+ax�K� j["@��  ��e�� ��  -��IZ�    �V�6��p�  [@ ְ j@�6ݭ��m[` *U�� -��U��Zt�h^���Z�-�m �i ���ʮ���`�P6j����m]J�b\��NO=�UuTʎ%�����M�N�kH�n���L,�:�J�i�` �j鰫a	���\U`���	]j�A����=T�]@� m��N��� 2 R����l R���� )Cm�)@A����� �p �@
P`8 p (0 8��  �J>��� )@A����� ��m왺�N])�m��
1�5#��4�[tm����ϳ��"�,�u�YNӲh%�v�8��T"�n�m�d6Yl��Q!�J�J�`�Vl��v��]��H����Z�k	s��ժ�ծ@��
B��ڐ8�����ZI0m�KM���a 4Q@m*ѡq��ڪ�m�5�6  �\6 �k#l���c6����$  �f�Y� KV�m�6Z�aa�i�� H��ۀ(�2�lհ6�3llXi     ��o:N]6$�~�|  �� � ΰ�M��d�m�6�M��D�m��Ձ�����m�kl�m�[�/-+�UQ��T�a\ �� l�rpm��ٺ�ڨj�av@�`�` [B�    ��Aa�Z�EU[N5+�+8U�i��$� l ��i�V��;m��m�m�c�ݯL� Pf�+r�T�
���f��X*59k��h��D�! �TYZ��X&XA�/�|�8Wo�ѪL�h�m�i��m�Kv��y�l @ �a&�=��`m�U'�� A����[��^�5O8����N�tt��&"����[:�U��leƄ�p�"Izd㦤x�v��E���Z�x%Vq�
�W��
����8��
��`*�Z¤.�*P*�=�`*���*���"Y$��� �]�*��CJ���7]+�'=��\Z��VR8�M�gm���Z�A6�/�]��`$ � ��:M��^`�I۵�Vm��jه.�m�
��ƃ�aV�!ж�5Kc-�;ms�z�AKWU@R�@6Z�Z��E�J�QeUuJ�l�*��*�˺tC���$�,KU�m�u�F��P;URp�Ҫ��]U�s[c�������p��J��C���\m�WN���̹%�jB���0Im ll>��m�vکI�56�,cj��xV�Bې"@l��h m� y�۳i0�.넭�i� *��@[V�c �g�� �Nɍn�udgh����b@m�l�RG� ��` p  ����{g����Z��6�M�6��(-�^�fə]�n����J�W��v���$��mv�*۷��۳���*��Vʜml���s.��V;�ݶ«�UU+���&8�WnmK�HRۚ'S�ۤt�@vu��r�'Y檧���ϔ�s�;#WUP��\��`͠�]�VU�������m�m� nӧo;SM&6[$� �'\��oIz���i2&�#T�lUX��cnXƫ�.���.f��"���G'I��L��Pݭ�籎wjÁ�6�kأv4���E9��W(|�P���~p�K+Fs������6��U�p�tJ�6�
���Z��]�{v�8U���]J�-�HD�T �i��m��% H'�IoW5�)P�k�����iUVT���l�Bp⹪�� ��   ��2H�$�M����W+e�P8lVQ�L��3���[�f�km� [@ ;ZŦi���7^�@H�Ͳ��-�m��I����4����H H��,oR��UP�j���M� $:t������k�@���F�o9uWT*�F�\����>*�]�m�4P��@��z�6�ʭlA�8m/. e�bE�y�ݷ`���    UUU�<���|~/��Ҳ��N� a�pp8qm-�FY�m�"nY&Ā6��l�����pr�1�E�S*9����F�V�s�n~|���8�7]r�u��LVT^6�2 ��&]�5�� �ԇ��-�ޱ�z!�]Y�Ѯzt9�H�Y�t��f�K���u�M�WfZ�� �m8�Z-�h�����׷aa�$�����U+�nO��V����X[*���T���V���y9�a�� �t���$B��c��m�í-�&��bP�c"ԫW@U���_e�x�Q�-�uL�B54��[�8����hWh��OUX63�"�ݱĻ8K�*6��8����=�F�_��O���]�'�j�*�P&+�".�h�7K�6mt���T�i���ڭ�m��iЫ~�o��_�m�f�U�u� d�H�"�Y��q/ �UV�h��xb��^����X�C��U���lt���kz����M-�R�[l p ��� 8����)��` �-6݀$nI ���l� 6��V�N	����$5��8X%�m���m���>�|�kXm �e�H��\-�� 5�lpm��M��5m ��l ,��ά�Qt�v���L[O�wNft*ʴ<��.�� m�H ml�Mp��m�ֵ�0�,�-�#��� �[J��UJ���f�Ue�&�Uۭ;[MJ�۬3��/�������������f� �?��>�VO���|TE��i�ADOF
!���w��?�L0�
����5� lD؃�EXA��_-=Q�EC���� h� Tt*Vg��,�� h<x����\�Si@��Sh%qt��&��W�E"�:��n���/�l5�v F1�X��t����� ���Ov�p�]qS@l��ƨޓB�M"��P��/���A5�����#�pP�m@2e�I���> �"��-Q�8�E_oB�⋁RQ=M`x
�銪QG�  @�+�����$`F0"ŌHF)� 0���	��BE�FUg����H� $HĄH,\E`�D�)*��!$��#	"��P�@`�9�@ ��B����`őX� E�B! �a$� @����>��fi�b��F$bA�) �$	�A�@�hn
D 8H���H(E4���
_QCj�(�� �q)�Q=6�=1JC�6��LTت>���!�!�%�� ^!�D���E� xY	-]�������Z�r�C�6�X��_P
�\T�C�E羪XmSa�X����6���@� vxw���'����  hH���O����!���AdP��I�I�IAQ� a�II EVAQ��I�I�I�IFTd	�I�I���D	�Y�I�I�@AQ�$D�I�I�HA$C�I��$A$A$A$A$���I��7��$�I�Q�I�I�I�Y�	$HdA$A$A!�V��A$A$A$A$A!�I ��  ������H1�	 �	 �!	 �	 �R$�H# �	 �	$�H$�H$�H��	 �	 �TI�I�I�I�I�A$A$A$A$A!�IA$A$I�I�I�I�I�A$A$A$A$A!�I�I�I�I�HA$A$A$"�$A$A$A$@��I�I�I���B	 �	 �	 �	 �	 ��H$�H$�H$�H$�H$ �	 �	 �	 �	 �	$�H$�H$�H$�H$�B	 �	 �	 �	 �	 ��H$�H$�H$�H$�H$ �	 �	 �	 �	 �	$�H$�H$�H�FDF��I�I
�����Y^�[�{�O�ߤ���zN�?���  � K( m��   ��@ �� 6�$      �`           � l
��n;���e��e݌�lZ]"�T�)��LvK��E� +�tY���5@f�m�j t:*��gj�F� l���ݳ$d� �`8 p (�� �J m� E�� �p �@
W  �  )@A��Α�  d �o
�-� �     �     �m�       h 8 HF�4�:����x�`�ظ,�`-��H0�t�-�J��U^z��QƳ]@��q�{{6��\���g��g<�6.���] m&��l )@A���� )EӶ�MV»::4eKf�w-�st���>�'m���b��Wi�ث��TGa"�U@YA���%�$� k��`Û��r�D8�}d�]�������Q�f�n[[ ��4��iHZ;d�
R�u'��s��^l��Ƿ;m[=ґ2��Ws�QAU�f���F�>�;nn����We�/�Ύ�k)��p�i�-�t��y���-�0�$�f�8LZAG'X�Uy��Ɛ���;n(Sˬ�(��3��.����`�s��ӓ�bպ��6����14s�k��;v��p�'\rn֥	n�]���ջ%��4���9hA���/\�� =��Z�*�Y�h��2F%�Wk�8螁-����\�g#մ�x�LF���:r�[qc�uX�T��qm�@7�e.q4���n�e0c��:�ev�a2�=�N����Þ`:���얛���Ԏ��s-e���Z�yb��.#�ꛒɤw8y.8�M��U[JP){,�I��@S"��3$˪��������_�@B�:��@q؉�+�\��J%JA�^z&h@���+k撵��V�_/Uo�muӒJTH�$�7� �6�[N���$���q�5ڛ[R m&A�۶R��6�u����5� [v[�[,�8՗^��غ �R���i��ca�]���踲Xp6Y��6�h�omӉ���kJ�Kƛ�o��=67��=i�LKGl�EX.�w�s��ڠ�a�z7��XƲR�:%�þ�����n�{���W�����{(=�����; ��v��^�i&:�������Z��� �;�mZW�{[��+�T�	�Mw8�J�.W�.V�*�8xwEZ�ҀJNB)�.����\�`]���j߮�����R�H�p�����\�(�� S�VL��^�����#D����8li]���.|�`I^ �Z0��!���L\�e��6y�����U͕��IٲAU��۲����.�0:]�Rh��\�}m���X �W��h��� #�R ��ʺ0���RNs��tq-\A m�0�9��U�����Q.($��JmS�M���́v����뷰���/�����椄N�8�J�$�0G���`�,��� �rM7"��v�U۹�/�Ŕv����F�m�r5)�q�:z�vȫV�4�)۝P�.�ֺ�뀎���i��ƒ��J)9�{ ����r��ۖ��]��}=SV�$!Ju)D����р%INʒ� I+�2U�]`r�%)4�Hpǖ��ݭ��Q|��UQU�u"]�l��6Q~�WM��RB�%9"�5�k`~��=w,�n�l^�h�mȚ�SM]U� $���� J���9RS�n�߭��}���2��-�I�W���3��Ssn ��x�5��k�ئq�𝧋��&�.&�*�� �F �%8*Jp��V��n��Pt7C��I[���ʒ� I+�9%��{��VT����nE�=n�l��lʤ��3u������GlUi�JTBr5[:��,�����ȮS�����>YIN}=SV�$F�JQ%$�������v��ݭ�E�����ƪ*H�m�l��+n��+-�ek#{9�ַ�:�+���T��F�JM8�NV��wk`r�� J�} �yH�T8��r(�"J�G�=n�l��l�J�3u�1fc�{Ţ��"j�)�F��I^�,�JJ� �IL`�P��IIʚmS�M���w�-\��=n�l��lv�m�Ct�椄RF �%Xr�� J�Id`@���{��_~���m�$�Ԓ�   6ٶ�zYպ�t:ܺ���껤��}��b҆�k (lD��Υ�l�   [v��s�gQmgYZGn�W/[dp �Β�J����T�}�4���'Wm�@t�E�Uɕ	,�bۃqm�δ�|&E���2D�����@��ݐ[VS����<�Ǒ't$;NY��޷73���gk���z��n��ww�+�i!�ֆ�=:vȪz�Mx~�E�i㛁�>����y�雜ɋ2��OI���w�� ]ݩ�=w{��k�o`{�V������G�.���ʨ�K# R���%=��|AvX�ʚꔐ��R�II6��r�����Q��	%xtt Ȓ�K�����&���� HK# J�Jрu�utڎE�IRH����[ I+�9+F �%X�R��&ja��.K��d������m�;X�WM�H�����U*i����]����`
RT�ﾈ��M��:��,�Rr�1�I6���V�
�QZ�#�0X�D�$�����B_��[��r縋I�Z��:��I�� R���YTȒW�r�F�xV=�� H�zNG��U*���lw�$��M��*\Ú&"f�蛻������%h��� J�u��X����5D$��㎝84��l�MchN�k'zZK���p�3Ϣ��7D�M�����f �%XId`Wn�z�V�GJQ&�@�6��b�%%��	%xJю>���&N�.�e6��IIRH�ff�`wsR�<Ry`b$9�榤��s��$9��`ۑ5R�Rn'+yZ�H33&�����`���9T
�TP]�Յ�U��ʒ�uZYZ�Y ��l��ƥ'oA�:�P6ES�v�g�R�{]V�Gi��㛙B�˨���t9�$MŰ-]����l��f�� �y�i#�b��G�r=�Id`I^ʒ�JJ��J�SB�R��i������v�Z���=w{��}=SV�$R�PII6}�舂�[s�29m� ��F{����J�����s�갺Dt�i���ĕ}1˹o�r��y,�oФ8��WsO�a��.Km�@e�i2�v�Kϭ��.�خ��t]HL]��ev�mY����N[ܳ�_ܼ�BU��G AUWsS�]M�|�W�/%���}˹dr�D�����4�rI�z�w���o^�z������ڶ��SR8���.����^�ww++U�/=���լij@q����^�z��ww5���]�����ֵ�j���INH޶�#olM�   
��KE��V]QK�Yd �\�6��� ���6텷mm�   -����$�i�yy'V��� ���n�/nli�pY�����]N���ՠ6�Jܱ+&R����v�r��:G�rZ��]��ay�F5���vۜ�������;�2��n��*�%�mֵ P���W^y*�w��;�����䝹ʠa���jZ��+9��5���;sW`xmKr�횮1���ǂ��Y�>ۼ#�%���S˹b򛉒&�	�����y,�D|Cr���O>I+�W���ҔI�G7��Z��׽]��z�w��_���j8I*$�9"��UQyi�ͷr�Y	JS��G AUWsS�]M�x��ܼ�t�w,�{�UWu7Rmhl����͎�k��M�	sjɬ���њ4�Z�O	/e��j���������Gt�w'}��_>n]T�PUE]�2��G�׼�x*�E[�|�h�woW����<\F��G��z��׺�wo^�����Z��Ui�IJ�RA�^F���#�%��'�L14�FC�E�Ԥ�Q���ū�n�]ּ/Zׯ�{�p����Xz�\RE�:zdq���N���;4���h���{-�l�e�y7b�Nh{u�;\Q7��]��wO)��%��J���er��N��Q�BTi�rE�_��\.����׼�k*��������mȚ�SN:�������T1OW���~}�*�	 ��
.�D2����e����.��f�^X�B��X��.�E:p����wD�Wt�	qh��XƂқX0!!с��ƥ�U�!�Vie��f6Ai�1�)H!+6Q{�^�K ��v��4�֠4@�Q�e�EeVă#QH��%{(�4DS�; ���wzT!� �QQ`��嗏�Z*2yEɫ����h��2^�XF��M�m��c���5
 1�R��%��AR��$��HGٴ��L�Mh1!#��Y�bi�) ! �B��c���qB�-��BV���P��0��J�3޳�*��׾z&}�TM������󈏭�9Z��R�{�> ���R���*y� "�mZ�1j)�^�ZRE$M��qI�l���\���Օy��$A�k����_;ZRE$Nw��qI �������H=�����MaY���zWY���E9��k@Ȥ��Q �����I����Ғ)"s���u������6bLnF�m7IE�SD�i��c#�:�q�z����˴=�]��Փ&�.Q�/.�1�̭�"�'~��hw�O+���I�9��{i��g 2)�_߯ED*"~;��G�MVr�2]fhw�O+����2E$N�]���$S���zR@dNw��p~���rt��ª�+$�������H�����]�$S��v�����# �$�}���p�~�����H����:T�+	yʓZ�X�)!� ����Ғ)"w����&�2)�w��)"��|�'�k�t��H��Q=��b� H1�����X�)"�#2��mG	%D���޵A�Pj�/3t�5 �i
S�~#����O�{ ��?ߩ굯{�5�׻�-�q��u"A6y��n��.�GZ6^�k�{[���+��v&������*��˫�褊{_}��I�9��{a�<�H�9�և�QI�w�;�H�~�}e|\���Բ^zR@dNv����'�Z�w��ZRE$N�߾��)"�W{�п�2'���}wY5�f��e�k3V;��'�}���I�>�w�;��5�s�Ғ)"w���X�) >zN��]T̗�y��^iI���N�߾��)"��}�iI�9��{k���P:�-}���$D��g�}W(�XfJ��u���RE'}�sJH�����@�u���>�dS��~֔�I��{��E8
�9ҵ}̫�UW��6�6�   m���s�i��(3�Z� �*�A9Am�R��Gݰ��Z����|  6[%q��G��We��e��kl�pX��gV�62ݰ�TqZ�Gi�qI�F���K��v�;\ݹfy�A�uӍ�!�B;c�:ƫ]; ��m`� h7U�v[v��m�s�q��z���4��Kָ)��������=�~l?)�<��fs�k�l
�u�Z'�678_K�������I!��U8n��㔩��A�&��"�'߫��X�)�Jv��ޔ�I��;��'��s�JH���NI�S,�&cyRkY��$S��v�� �?$$R�2'߾��C�������4��H�;\�lw� TSڟ|Y�wYy30ʫ�32���H���}��R@g}�sJH�@HAj'~�����)�w�^� �IӼ���.�2��1�����)"���h�9��{�;�H�k���I > ϻ���$S�Y>t��Sr�!�I7�"�Z ��W�c���?1 #~���Ғ)"w����qI����) 2''���Y�S܉�,�p��J��i2��L�m��앶y���*�a��yxi���W�V��&����p̼�fj�Ȥ�}]�ץ$RD�y��w�I�{�ҠJ�H=���ֻ�H��'��K���+,�Ư2���H��;��D=<)1v ��*�P`J�O��3JH���+���p�s��)�@���"�dO�>���W(�XfJ��u���RE'����RE$Nv����D ����z\�QI�p���)�N�P��U.�I�.�4���"�D��߾��R@~���)QI��{��R@K�]�{�E$N���:T�+	��T��j�qI�s��) 2
@;�~�C��QI�>�4�H��{���)"�흺��ѕ3:�Z<��pJۦ͕�j�9l[6*�&Õu��Aإ���������a�r���{ĀȜ�;��2);�{�R@���ܮw���qI��ޔ�R�'�Y_#�mȚ�4�NW5����G��٠>5�;�w�w��O������H<�;��)���\���T�u��RE$Nv����)"�����Iw�1[��D�2����DOV҉�b� ��i^!�_Q*'w�y��R@g��sJH���;���d��^�����X�'�����߷zRD��Q>�����$R}Ͼ� �"�n'߫�߬w�Nt��J�ʙ�+/+�2���H��;�� |����٥$@;�w�w�N�9�Ғ) ��g$�����]am���y�ӶER��	�6S�!����v��9d�yۈ�2����77F��+$̕���3C�RE'����RE$Nv����)"��s��_��! H�QI�w�;�H�ܝ1����fK�ʻ��)*����s���? ���B�\�~�߷zRE$O�}���qI����)�R?�#7�?|t�'�YXL��ֳV;�H���ץ$�	Q9��t��|��Ĩ���}�RA�%D�՟}c����S�/���fL�2���̽)"�?) ���>��hw�I�>�4��I�v����R@�ݠW4������ �5��vMɗu�fVI����qI����) 0��1;�w�|�H����zR@dNw��qI�y=�.���VYyw����d��zک�9��761��.���Nxk��f�w|@I�4n��rfxar��fmI�<���ֻ�H�k���;��'o���`}`2)>���	"
���|�mT7*J[�l�-�m:�j�Z�Wx�`?$�H�g��C���O��٤dRD�k���D��	����}+W*fL���j�/JH��߻���$Rw��4�*@�"}�����qI�_}����H�=�����+�Y�.�4;�H|F���٥$D��߾��RE;\�oJH'��#�\O�}���qI��>-�XQS
�%�J���
�H<�s���RD�,$1 �}���;�~�C���N��攑I�x2{]�eU����$�`  �����g�7aHւ榋X۫pj�pm��  qXI�ݫ���ͱ   �l�j˭�
�t�v�\�t�TQUV4���6��	�28 �3ۄ=:8[�1'f�
��i5��ݷs�nɛ��R/<d�9��ָ�n'�������ed��9[ݷBrN�������N�+�Jԛ9$�~s����߯wp�#�N��P[hl�d�	[u\�Yg%���$�������w.�2�Q���(EXR9f�eL����/*Mk5c�FE?W�~�)"�';��C���N����	"1 ���b!��D�H���;�w�w�O�3���*VL�Uxa���$D�y��w�+� ��B@b-E'���Ғ)"w���X�)"��s��~��$BDX�P�N�'�e�f^VI����qI�s�JH������pT�"1�TCQ��߯JH�߾���$S�t�p��3
�1����Ғ-�G��\N�]���$S��~�)"�;��C�����Eb$T���٥$RD�߾���ɬ3
��L��k5c���v��ޔ�I _�)߻ߦ���Ϲ�٠*5�9��{c�$�)�?����H}����N��*�kbhkÞV4���H�M�*�3��tVe��) ތ���ʙ�+/+��Ғ)"w����qI����"�';\�m,��CȤ�}]�ץ$RD��'�}WU*V��2]fhw�I�{����{��ҀD&�ኗ��|����=���O����I�9�w����'� �������U�.�U�f�������;�H�k���I~X�Ċ� �D�����"���Y�$RA�N�ҦYX]e�&����RME_��1R �F g{��I�<��}��RE��{�Ғ� � DJ�߫��c��z}�Wu�SɕW�fe�I�9�w��$W�,�5�>�4��H�����;�H���oG�E&�{~n�O�Op<��qr]�(u�e�/;v���8���e��%w32eL̼4*��"�	��FԎ)Dө�k��A�Q�?~��H���+�����;zUO���=��}��RE;G�~����*��0Ғ)"{��{c�~ �/��_}���H���~��)"�����$@>b�;�~���ɬ3
��L��kX�)"�W{��I�<�{����Xw΋a��?� \R~�ȵ�=�s���$S=���ܩ�3.��̽�"/�A�����K����5�~�iI�=�s��ɸ��������Hy��2���+�Y�K���) 3����$RC�?�_~�c�BBE?W�~�)"�'���ָkTZ�f���*IȩI5��ɶl���$��ͳ�g��.���[�T�����VMwXQS*�S%]�mI�v���;�H�k��)"���{��RA���w��dRD�y#޹EL.�ʓZ�X�)"��s��?�0n)"s�߿hw�B�w��Ғ"s��{o����6}�Uu�T�ɕW�fe�I�=��}��RE'}�sJH�W�py���X�)"��}����H��s�vL�����cfe�qI?AO���߳JH��߫�߬w�O;|;ZRA7]S)�FD�T	 �<���$wZ�C���{Gw��0������)"�'��w�;�H��ů~�٠dRD��}��M�$Rs�w4����O��j}we�yyvHd��=8��N��%�@i.���.#���jxne
7^�����u��2kµsS/+Z�X��I���4��Ȟs��qI����*!��*)"w�߾�٭PT5U�_�D�H�r�RM�T2'��;���� ���w��4��H��w�w�I�y�� ����""�"{�RE�ߧ�?U�*V��0����RD<�~���JH���W;��	�w��"�'s37Z�U�֪�eMb��4TDrmI�
E�!Q;���X�)"�߻�h}�Q$��]��)"��P J�;�iI�;�$~��*ar���&�Z��RE'��sJH���'� �~��C�RE'���h�9��{c���P�:i�{\��0����M��t`�ŕUD����f`��a@�_^U��1,ѫ3�,0�;<B���E������
�d%��Qf���e]����`ʽ]��Ku��矂i�hXRP�=��1)�s{�T�(��D�S
.�M�a��0}�"[��QWA"`����!��p)��� �r���g^lSnІ�KD=�Lh+]O2��yy�=��3��^K�	l�{���w�M��   � m�     ���  m�-�                 � aC �` K��m���Z�mZF��7��r�Z*�M�Q��f鰐�gI�6�,J�<i����JP�Nu�4k�:S^f�����L�7:` �@
P`8�l�  �[P [@���� �p      8���� �o86ش�m    p $   [@              m  �	f�h��$��m�i -�n�m�`�v���� ��h۴����R��,ڛ��-3��d�#4M�5���g[���(m6��|q� 2 R����S8��m�XZ[�Q�@�w݃Ƙ�h�g�����K�4Ɍ��f�R�UN�k4�U���/A%�i�E^�u��֬[��0��k�F����צn����82v0褙.�u��$ȳ��m�dk(����44�\K�����P<d��'�¦�n�Qc>z��CR���(@%���瞫b^y��vT���<�vפ�XG�X�T�$3em��a4�t>�v:ݶ{����]�1�&�tg��mQ�.l��.mY7Z�/=jF_A��Q�Q�s��>`�=��+��qUYV�d���j��[��*K��nnv����><���v�%��.��l�N�G`#CUW�S�>��������A;Z�,���ےP6�7q����ڵp�-�s���۷X!�㫮�nSa����M�l��ǧ��w&�q\^i��uXw�8l�vۙ�A& 9��:4��]�y�+a��r���LUu����eح�X���}�m�k��lH��~����/w�Tl'�)�Ё��!�OX&(�` `�bx�҆��
�@�=9��UUUffIT�am   ��O�Y-�� �Z��jU
9��6���8�%�ݸu-�knH  m���޷%�Ͳ���N��&H�o8���^��C�a���v�Ne�3�)2�;�]�v��^z��q8ڍ�l���<c����Ƽ�f�9�H�\QH�p7u�9�焧I�0��3�-��ndyƯ:�p�3A<К�2u��	Y/)����m�(� �&Wm�!��cy���n�.�֜P����b6^�l���ʅ�L��ˬ�Ғ)"w�����)"���$D�+��D<�Ȥ����RE$O{;��I�u�yXeB����)9�;��"���$��߿X�"�����RE$O{��C���PQӺ����*��3JH���W{�Ÿ��w��Ғ9~��}ߴ;�H����4��H���ѓXf���zkUy��$�	�y�Ғ) ����$S��w3JH H��s���$S�NWej�S2f]��YY��dD���t;�D#��E4��TӬ �j����߰r����{&[6�̱E͕��k��6��;m����̴�횮�w�r�1ue$bRmu��M�v�1��y>�Wki�`�b���bK����ɪ����v����u�y*S,B$���"��)��JCHB�P;�DƊA!M :(�>�y8��{��2e?��M�G�@���s\U\�\��yZ���{��kT��&��~�|��S)�ԈWq6U�M��}�Ot'y %\���h�^M��=��R8�IS��� \���DJS�׀;���6�8ڪ�f���Ԥԍ"pt�0��N�:���Aa�V�W [&��ש8�;�����[ܦ�IIʚm5$��|�P�+�%��Ȉ�����H��-�T��%-�ddܛ|�{2n�Z���e�� �7xU�����
Y9DIvU�faW���	�{��rB{�{��1dB�)U�'�0da�B	)���2#$	��B`�������� ���s���)*O�� �n�@l{��W(�X\��&flܟ�J��Db��+_�W@n��Հ�W��\�!�D �{��kP��N��XUC.ꌩ�wW��'�߼�r�~_hO�	 "�����<��ـn֫���?��*�w<.���Y��5���\'f��&ڃ;oa���X�+�操vM���"1�N*7&�@.��l'��;�r����	���!P�;���>���SM����$�M����p��C��9!��� J�:�y+�"��*�� ��|�#��s�g[�������#�4��@�z� *�
����	)5 T��¾�Z��Dp�M����}՘�F=*�X���}�@3���y���P�)m�#&���P�d�$��O�������{$�w���$�/׏�=����M��%�T�$�+��ҭÝ�䨵�v��m ܻ.���5{p8�ȑ�Ԓ��NP���>�@�|������p�G#� �n��h1�M�����w{�t�u�G� �t'ZOsw�s��ڪ��w�u5�RED�Q&�`��րw7y��{�t�u���e�����Q҈���
��ܼ��"7�t<�`}��@�ru�S'���-���RM�w2�|U��^�{*��@<Ӽ=q����/�ȩywUV�$m�6�   *��n=8#�OL�m�@2��6����@۶ж�  ~C�'Gf����Z�DW7]f��Mm��곒��sn��ob�����m�Ò��ݏk���$��!��3T0�v[z�<�M�g�6!��u�Y�A\s������W���=W)��k���6��E�)!�`�Vg�X;��x����;|W����zB;B۪������X)V�&ճ�ry^��+��.�Ҕţs���:[�XU�րy�y}���iA�WW��a%'*i�ԏ`]�^>��<Ӽ[OtS�� �����6��&s�//2��;�5��O��G�}IX�>{1�|��X>2�#Q�%+����>��m=�O'Y %<�ht�Z^ɓ`]w��&*Dd�I(�s�5\�lD|����ۼ[Otq���|>u���Q�l
�u�Pc'��nrs�:��P�.6*��î������t\�U�	W'S��w��Oc�@��ǰ��5"7�*77��;���q0z���o_orO��c�o׎����UH�}�O��ԉ))��ԓ`�~�>�
if<���Qv����ɰ;����#��78q@�"Uju��N�>Z���DD��|��+>��	)9SLm)��~�|�4� m=��u��G�2�u5Or'$�q��Y'`^�1�njNn��s7���Β�wM�j�~�-���>�h�w����
y:����1��
^�픉�I)E$�̼�?PZ	�@VW����Rﯿ~���W�̛�11R#$JID���z��I�_���R��"��)@hb�@=4�����(��o�ԓ��}�~2��JH�ƪ2$�{
�kZֿDs��_�?Հt���_@ϖ��6}����k3QR��Q����r�l�#�"#��<�:�t*��¦c�r������+�s��͜G��l�YqPD6m�*�g��9����A���������}}r)D����jI�>��~� ���[~����U� .���_��FԎ(DSDw�ϵWb9��� G5ΧY鐉i�t	�;���(�(���.�L²�+.�����Z��@���O'Xw1cj�R%��I�s{|UGr�l	�;��rNW�횓��
�$i7UFq���nŃ�(JF�RJQI6�Ot�S��ι:�4� �p:_ɺK�:���N�N���u����R��Fcum��qYߧu���O���hZn�H<�`듭��KN���{��WfT���*�j�"Mǰ=�ُ�j9�sj�]��Zy�l�UvG#��Cr�_}��D܎���|�k>���y���ǰb�c�WRz�eL��R$��RM�)e�������^�y��U_=;y��H��|�#��wy�}>�]��|���K0���"FY'�]��3.�ė�$�~~  ���.��N댜ݺ:�V�R����i2 dp�q m�8��ͱ � 6[%Ν]o<ͱn��yΜ��r�d�5��M���8�۬�de٣�%�cH%�4����:�����un5�V�Oe^��Z K����Ll�Xj��u�F�n��N��c�7nI�h�89C\��L��<u�0��o�o�ww���9��w�2��-�I�W���3�mѪ�����u.�NW�.�a��;��:�+�q;q)O���~u��Ii�@�f��
i:�;�6�� ���&���r�n�kUET�֞`
u:�U䫘�9�s�{Q,{e"F�RJQI63>�9�-z��c�c���&�x0��H��)$&�#��ju�5ַX��}�"V�����pLM�L]3Uu��s�ց�w�.i�
y:�=	��?�tvz��Y��<�깲�Ƭ-do<:v�$��W<,�J���o|�����0e�V�y�x��
y:�� �U������mH���mI7ċ�g&������B y�4"��<)�`|5I��4�>Q�FԎ(DSDs�V�x�qR�<�>�"*�4�ɧ��66�U�M�rn�n��w ۼ=2�{��3w�> �Z�� ���!6��J<Ӽ&��
y:���6�H���W�J�}����N��*�k����S��ţ-�xe�	8�nX��L�jV�a�A����y��ϵW@�O���������"2D��Ns�Z���Λu�i�@	6�@\8�a7��JPMǴ�Ǚ���ɳt������<a��P�xȐ�t5)i(��4�R��t�6FJID���#ES��t��TU����
BS)eABM!("H ;ҁ^ �uaj�H$HsHl��Oh�@$�#��a%�dI �$T d�B�%�E[�z�2J�2�� �Q)�e-�ʄR,˔���<��k+Jx�J���!�Ҷ/�f{��̬ד/��}�P(� �uh�ΝT��t-�1UCv>�b"��w�8��U�⦕(�A
Q$�����o�WU�=��fj*Q7#����`~�s�>i�@I���FϵW@�<�ǝA��y�M��6���ot���;��&�@<Ӽ�=�g}���y����`P���&W�m	O6���DvY�h�Nt�ʑ#jeE�����rju���� >Z��g�&_����egқa%'*i�ԏt��*�����0�j�������r��H-�7T��ۮP�Ϥ��[��&�@�I��܉ee%�]Qwq77w�.i����N�Aݬ��AF�0XP�U(*�ॅ�B�CQc���-i��R�M���Miv@&��lP��h���&�ʿ�&*Dd�I �� S��`�Q�A��	4�@�X�ʿ�v�VCR�\�Yz5bk���eA�{���gZNΩ1�<��v8�:�ɪ��9�N��;�&���H9O��ya���T�n(Q�6�ܼ���E�<��S��`*ԫ=2z6*�MTȢp"��$�ڭ%F_��8Pb���c�f> w/&�9g�0#jG")���C&ru�2'I:�i��|.i��]^F�II�SR6�{�;엛{�!����{��)�� ߭��D�D�B�!@M*��P��5B���v�O���ϟ� V����  �f�Y%�ۭu�[�&��fU�%X�Y� m�� ��8�n�:�ݳlH   ���4��Z�X�r��:W/[d �r�I#�|O��+�P1����g���n����p�,���:��œ<��\�ϴj�]��8Mv�FȪAڋ#��lu�y��Z�}�+�	
r]֛���^�%mp�X�^@c����r��$�f^ۭ�zqm�*��"Y��+=/�8+`R^+0�s���t|�|R��d�v^]�h-?׾�#���zB6v�~�G2�Mu����K+(�.ܦ�%(��/���5�����[�=�ُ��ɷ��WkZ�^��&*De����7{�)I�뛭 �N��� �R��R�㢜q�+Ty�7Q����{��m�`�>��T�n(Q�6��ɰV�����B�N���s�ր��˛�����0��b��^S�Hi���!���wC랛�C�u�)��96�D���mI7@_��t<�`뛯��;��Q�]5#��� ��ǺZ޴�UZ��0�� `$!� k`Di�� T��Q��J��5�p""#�Ŕ��=��Ѓ|�f7Ȫ1W���t�ԩ�R=�;�����}��<��O'Y铹�ک�6���K��w���Ds�G"�u���0^���<�~�|
>����D�6I)\�Y�.i���Vι��4���g�Lo#E1�M$�'	b��+Y(�E-�h]�5�����v�Wo·���AI�k׏t��1�
;��`_���eJ�R�JQR�q��%X�ʠ����<�gګ�
w,53QiD�P"��m��yS`_��{�6��������W|��I;����rC���mH��q�$��y�k׎:��Ug�;�#X0�����.$�����6}���':�|@zF��˼� [���Pj�Y�1��Ԥԍ���%6S���k�I=����3���Uʅړ���S�#l$�MJ���#�1{2M4� ֓�>���u����M��d�v^]�h�w�i=��Z����/Uh;굂�)8�%����x�՘�*�� #�ηXܼ��.���*2AH����Dp�[���:��@�;�>�G��A�����o�.M��pLM�L\U����	��:D�xi=��x��<�-Si�Z#��A���D���6Q��M�wm�m�c���+���m��t��\�\�[y: �w�&���Ns@^zf.�t�6�Dr�8ڒl�M'�t��	��: �w��<�a�R8�@��s�1�-�y阸�y6��s�yU��m����5 ۹�>DE�R{m� ��W�5n���i��n]T�qvNae�^N��6��4�hݧ9�	�{:n���/?cmm�F�؛\  
�UWvJз\-��kSWM��� p�Pmm�m��H�nKn�ے   [Ck�q��mJ��+�[�v�B� )N�kxѯt�+�[����ֹa�d��e�/����l][K�c�2E������O�>s�|6�9�[p��n��Mj����Ml�ƨv������>[0NnQ08�nD7[M|�0���;{$�G-&���q��Q+��Уp��Z��q��:���<�C۰�n8N�S.����@rO���s�'\�{�v� ���M$�Sq�H�����m�i�O���$��/�Vg�)h��nJ1T�"r.��s>�-/,ͽ�۵���Kv���8�.d���.L��o&)Z�X�n���S�q.�����y�&Ԉ�QR=�Vz�qrB��9��N�-:�7�����g��hl����W0,]�G8Y�Ln�s�c���x;q��iJc�nHo���� ��Zwy��=�����	)5*jA���ۼ���V��ÓⳜ�O":
o���՘U�zꪴ�����q�%)�Q$���8���`V�0|�7I�@s����Vl�(�$�ԏaՖ�9�3������F�e��Waf&�U�%ݗw�t��y�z��`&�@*��1���MJzdq��a`U�sPcC���w'W:T�zS��g|���|ؔ*Q��"F�U�1{3'I,�{ot�9�5p|��2YUsarm�e�Zu�4���Np<۽�ڑʊ�MH�]�s�f;ű��B�#�J�^y}��~�䜬�{]��DmH�SM	�p̙���%yS"����j�� م	�U�� Tcn-����'��/���g8/^=�WU^<��jISMSQ���嬓�/]��<]�Rs7I#s�V�]v�2���9)H=¤�S{���ũf �ک䃖���r��%�]Qwqu7u�M��u:�
V�yS&/^=�#+,6bi�qHI9��.N�-7z�N��{����	�&&蘸�����9�4��T�[���y��r{�S�H;��s��<��y��\��ʫ��*����Ut;.%��������o2p�������hl�g�+n�6V\T�ٶbk��!�Bm�/4Pc��6i�sOͷ�����O�W@S䕿��u�<Ġr]T���\_*I��O�W_.�s��������� ���	)TԦ%#�y�zt��&�@rӬ�n�q�%)
{�I7�8Y��l]�W4-:��6�@ơ�'h�.�n����� Ij��9�Xl˔�� �o��I?����3f�9�d,�T �JXJ@;�(��r*P�$D�*+
X"S
a)*��H%b�:J�
BR * ��
HD����!�2P��7�2�5�T��]ן�׷ޥ��)*��TN�    � m�p    p [@  �                   0`l �RY,��&)jV�P��87��z�VRZU��U;��$6�U��-p��3�������-f�5'�^nݨ�ݙz�X26��.  (0 8�4P8 p (k@  �J �    �g 2 R���  p �Am�����    � H   ��    m�        �  �8mqf�]��lk]�-�6�WU��m� -�l����Y[6䬢^0�6ԶLR5�v2�a;s��x]�iN�X�l���8 p (0 8��	Η1��1�:�����v�w��;�z^y�+�݈ƣ'h��q�l �]]6v�� m[W)9vͅM�I��u�l[M��-$S����v�VF%E�E�sն��M��5�+%U;����;&�q����6��vd��4�&L�VS�W1q�=���FW�k�psYְg`�V�0�n.g���T#!�^/iN:�%�.�$�ds��L��U�mn'�u��=�ƺ���|��Q���0g��ݳ��d�/\]����t���n;g*6�݆mŇ7c�$gY�f�Y�S��y�5�N�'��SS'Y��p���)�z:�V�nl��u�`E�4�]��I%���K7e듎 �$�:�q�q�����U���ix�	���]v3ܲV#�q�p���%j{u˭�<Z쬼򗑂������w�J(�)�/wc<n��.vxzn�u���]ҝ�c�t�s��V뚺Tmغ��v�[=�8���X�nU��ө��0�U�Rܪ��f�I�1��@���{��{��lZ��Ci���/�C�@�Ne�j	��8��-X�����_�@j�^Z�V��� �[���^��zsK��ꛮ[�kY'P�9@���2��$�aml��  	-���/X�-m���t��[ֶ� YVp��tk6ir�[�΁E�m�����Y�]�+�*ut����]b�I��ֹ��+c�q]%��n����`;d97jL��2�{g�GR;�m��\����<j��/Z�&�\J�׻�_W;+�7Is�Z<���"��6�u����R��Y3�6ֹ��j����Dc��Aɝ���y�8c�[/39�=fT�)B�PJR8���%xU�zԖ`
V���>H8�,������˾���9�T%�dɾ̆�q^Vd���y��R"9N%us�|�r'm����@S�+�<�ql�wF"6�qB!��p��68�DL��M��'MO@^If�L�~�{��f㇖�$�֊�3�m�ԝu��n��«�E��sԎ�5k�j��)7x�j����f@�+�QU�Lx�a�JA�&�M���w�m���R0�)�6&,J�U�G��$�y滽�I<�{����̜�u���S$j5$���`g�{����S�z:Ns�G
�4�Dc��BI����6/^d�E엋`e�3��eMb�-*�U)Dԋ��&�E2�<��6�@7x����?�u�=Y�3<�d;R�꺹Yn++Y�^��}�Q�s�����6�z�Ybړo3/@�I� ��� ����ݾ��t�6�DsQS�7��fg9�j"d�M��@r�w��j���n���Ԏ*�4��� /ٓ`b�̜�kV��X�_��	��}��$��y�:��u���H���ɰ��|�>�`�9��,��W�=�T���.&����3//@�I� ���dȹ��1f^N���Z^����jT����N=:vȪu��,�w򹯎�-lۗ����z�37Q<�De2D܊IQ7@���~� /ٓ`b�̜����Qaf&������� o����L�u�x�Nz�Y\��*k�iF*��jI�1{3'��S��/ɼ���@�x8�,����������9�s�&�=����ת�[a"�) �P�X�]�ܜ���6�Dr��n-��if o�����+�<�T���q�j7���Twi�f㋒�@B�#T�y������s��ˮ�Vn':�etXڙy�i��� �����n� �I� �ou��WY[�6�D��M�I�1{3' �S��9și7� ���G�iU[JRz�M�ss�{��.�;�䅭�G2Aζ�rCT7Rv����n�.j�p����� �w���v��^��HTD8��NpG�&�sͻ�9�s�4�݀'�[�G��菪��j�V�����G$H�T�ۀ  �6�^�'[7<It:"�Q�����հ��I�  ��A[�q��ٶ$  
��V1�PR�r����:W-�H)@K�;�<�f�=�*QIB�9��$���7�8U��W'vcn��n��=��6�s۸�3rzډ��x���G�7v�hۘ���7�c��#-�bf�p��^�|��w����~���D�oRkz�m�,vt�"�v����㧆�8��v�Ht��iF*��jI`|���pe'8I���ɑt7x�o�&.�.2�}�ʵOL�&� �}���2p�S�ڑʋN$�[.�� \��}2盬�����%&�������̓V�w��uz��>�j������U���i�$&�Drluͻ� �'XI��sw����_�.�+6y�ŶȪz��z�a���ݍdn¡�]F�e���+?=/ʼ�����������n�U�ѶS	"D��R=��y��⪭h�Qڭh�kU���6+�d|A��ǿ�>������#�)9�6�}8%�ށ��� �otË��̑7D���Q7w�9���<�a�-'��瓼A�@��AT��DrM�p/^>�-�7�5'}O�+�G#�	�}EG�������^S�HB���/=ѹ�>��n�=��.+��\�in9����� >�W��R���t�0�����JTIB4�� ;�ɿ�>V��S"�n�����66��M����F��[A�י8W�ɕ�4UWT���H��4BPE��1a	HB�(Z-�5x��F1� �&@ (]��w���V�I^}�����n0� ��$���8+O���� >�W�|�u�N���捲�HD��������B���}y8���ΖbLo#E1����s,Qsek#�uV�miv�3��2�t<�䒊HHD�8��Np�̝O��x�ک�"#$ȗ�O��b�򊐣JQ�I6.��p/^=����� ;�ɾy��
��A�G�fh<�`�Ot��Ჩէ��z��`&Ԉ��T�G�3��� ;�{��v�����H>�Ҡ�]��ޤ;��6��)Q�)9����s��jw�
u:��j�״UU�Sq)I����HJl
�6:��E��\�s��7N�GSuL٤�]͹��"��k��uJ�n��>�J��ڱ�P��`]����Rz�M�����ǿ�H��� {[����j�s&�n��Av\�]����@~�� >�W�̹��x�Ϟ��x0���#�)9��w�9�'zO'X�K�'��Т��!F*��b�l
��^N�k\�y��^}��}�6��by"I%$�����   �m��/S���z�q)˫;6xj���iCm5�6�I�^�:�ݳlH  m���޷%��h:��N�I��l� [���@���\����u�[=+ZL�n�*q���Ν�o;]�wnur�;v�v��m�Y<�p��q�n�6rTm�e�(����4��#k7^Cu��,�w	.�;��k��E�/6{����y��`���<��fs�hv��6Q����k.�[��,;q��L��
sPU�hQRnp/^=����@=�� �ܝ����	���#r�8���w�󜕤��̛��W���<�x�0�`F�r%*"%'9�!�t��&�@��� ~��@�
�4ډE�h�M��]���^�{;��p:��d���
Rz�M��������� �7x�rw����[�_ܛ��!4㇖�Wek��p�[U.�6٪�{9�yS�a�������rT�G�>��ܜ@wٓ`b��K�W1��x0�� ��%'8�w��@�p����w�u�<�7$�}��9��O2 Z8�9��&蘸������
~�W����Χ]�Nڮ��x*�*�9	J#�os�yz���OtO7X�sw�t8��j��K��
�����'����Ϲ�Щ�����y��R%P��ӨҊ�-��`��)0�PխM�lu�qǅ��*���m)2%*"%'8W����fN���[=��s-VVV�M��R��t��`9�7zO'X�O����_�Vܧ>q��JA�RI���p:�����^s��"�-��o��pJ��%�.�l�H����X$P���LP.�\�	U�(cb� )`P�F�kp�	�`6A���J,�&Y*��.�G�TN�S�x4Bl�
eUՖ�t�By63��%j�V]��a��yB@$A$A$f��R CHRR]$��y��Gzܕ)�=K�� ��yj��P�*��*ąS7�I�o5�n����v%��������/�{��/T{�p���qH���]z����(����7;��{z�y^������6�TQ�"���9�:��`}�ބ)��� ��sS$�%JQ���^�{(>�2t���=��p����jS� �t����Q�8�cG.�G��Nx����6���3N�o<��&���������7zܝ��>p�f=��x*�*�9	J#�os�z}����B�N3'$=:�t>�W�Qz���mH�R�)���>� ��u�L�����N�3��������˹���sw�z���zܩ���L�l�Y���'(�ӹuwYU2���K��2eϹ��.Rn��{��d�R���jISMSQ��*N��$��i3��]�G[������k��]v�7l���vV}ww������ ��� �7x.�2p^ٶS*(��`gr{�L�y���N�� O'y�:����I*�r�q�'8�������� �N�ܞ������$��.&�*n�YN�c� �(w�>��@�W7\�aWXATi�JQS{� ��&�q��O���u��� ڎ}9�������|�@j�_-l�UUUUUR����c#Y�b�*m3&�mt��4����86�8h�ݰ����  	'GE��u�P4E�nrv�v�ʵ�k��n�!�t�Q��n1��=�.�rR�+�Ұ,�]�[�Dh���k@�b�<���v�=��V�$.w@���[m��ݼ����UpBr���os�j�����;v�u�{���O{��|G䝬��:<��pJۦ͕�nlݩ��2��m�8Yyb�{r�
QHF����9�:���.�2}Z��Py���������T�DR�5'8���Ϲ���N��Ood:aE�F�Q"Bj:Qǰ9��2p(�����^s�u{1�>�V��k>q��JA�WwyY�z��V ������ �����1�l�"8��`{.� ��� �ͻ�:y:�=� ���\Is�Z<���"��\D���4ˈr���cF6��TmS��gBћ��o��7���O4�@��� ������u�T�!�]�Y��'+�󹿅L2¹r`�L+��|�w���>�$�|#�fR��F��)�qM�p�>��OtO7X�sw�2w�)�����R��&��{ל�^�{}�8����فQȔ���5'8������ �N�ܞ�72xd}��Op<�,�p�l�!MFWm�̝@��79|V{7m3rs�R)�u�W].�7s��w��՘��
����+H���뻼�̽ �N��Ds���O0N�]O�J��"d��Tm��ʊ9)�$�]���^�{;�^�������u/�נ�x�p1�JJ���I��UM�_�=���_}8<�x����p��!J*Rn���O���:y:�<�=�==����Ϥ$����ٙ�!ڕ�U͕��-@��6����r0.���&8�x��M\\U����<�`|���n�^���=���	�"�H(�{�x�BO7Q�)���<�`Ę]R�D�DT�)9��y�`r߳78����^g9䄪��#M��!*��`
y�zܝ��q���ޏ��"�Z�]j��y�����U�
Rz�M�^^�w'x4���zy���n�����CD�7��N�FFM�|uV_4��>�*Gc�&����3vg5��N�f��+�Zo0��U�6|�� �j����bi%QR�H�� ��c�H���z �w�sM��"&E���QPL�U`l�%x�mY�9�rg�R�η]��F���ɽ�p޼��o{�4�`8�J۽�qM��M����QSWU��{�GRn�>m��=�g;Z�c��1�0��X�UE0��BFQ#�"Q	J��]�2�ko`����l   �P�/gώ�[dn�OT`��4P@�LR��#�n�-�����F�d�$��b�ݳsCv�4�d�[l�p���7��q�vϬ���S�=e��دmp�<�w�l5�Ɨ�s<��)�x�p�E)��gH�7����mu�v���ɇ��m����[v�rO'�%���,u�/:�q��}��R'5�����3q��m�([dj�+�n�/=�:ö�h����Z�3vq[JMѺ������� ��w�t�u�y��@�
��Q"BTǰ-z�' ������� ��c���i#�u�̌
R�nooyz��V����� ��w�rf6m��ʊ9*E#�}Z�kT��}�xJ����O�<�`9������.��n��#����)���O�T���� �E���F���i!8�"kz�m�,Όr	"��us��-��h��ǌ��EHR�����{[��N�]�M�ܼ�p�f=�#��R�PUNT��7�ܒ{�;�֣��� i�j_y��rLWx���c�խj�I���_mH�N˻��������U�7թV {ڦ��W�̈́mG%% �H���^w���d|�����l�u�>Z�`��B�mD�	PtG �yx�o.^G�=�y���ǰ9�0��F�&�h!�zqm�*��"Y�-�g���G��-�x��.�SmS��
R�nM���/^=��Գ �|�<�S���51��(*����.���R�q'�[���Sw�yz���j�#��>M$�6�I�ܓ����jI����naW��I E���sh�(�=�o��I6w���$糮8��)EJM�R=�,w3' ����i��=<�`�8�sd���]�\�y�zO'X4���n�6Us{z������wȨ�-Ϙf㋒�`PyN�!�kA<��G�\-�g��޹��R�H���!��>���~�|�_�'��/^=��.�#j9�J�QI�����2)���:�t�Գ ���º��$%A�{׳2pz�<����������A:Dݙ�U^f^^���.��9��@��u��舏��
$As`��5��srO;�۹���xee�ŕvt-K0�V�X)�����6Y����4St�M�Rp���(����ںh�׮ؐƣN�A�]��٪���� �ڔI$Rp��f=�kٙ8}qb����"Fx�Mb���)7MH��i�zC�[0i��=<�`�|��1�
�I�#�{����6��9��^W�=������=����ӑJI�JN��9��@��u�)����l�9�x��H%R(�� ��������}�t-K3�L�����Ԟ0����B1�:�J%��H]S��(�.��!Q���,��E�
���G0�Y5a�T��U��,��H���aI��̠��C�(^!!�L��R1�1$�$a!J���*of�����f�H�B�H)B�}]�Z :��T$�a$�h*��I�T2��^�@$b B��uRvFV��p��!-�J DH�da�3��甄���@��,����0�RU&z�>!+{��~J	L�1!!S
}9~n��׵Y������^��i��    �h     8 H -�  m                   �  m�赸�9a�.��S`.����뫞�� "Z[��p��s	y��V��J���l�Hܧ� �7\l��śmF��dKA�v���   d �2 R����m�AJ  d �     6 V� @
Pampm��j�� �  �  h     6�         [@ � [@�mfh������"�� t�I�u��۶m�R�	�����3�n.s�ysI�pV����b4� p=�D��IS]�lH�h��� ��  �J*iq�&q\L�S�ƺ�@�8�d^���kk{/JW�j��#�ڗ�)m��眍�][0�R��t�V)j]��V����f���X�Aj�n��6�]f�����������kae@(Ʋ��c�1���#=n ��ue.pv�GkS@ �����'�����A{=��WA���lM�I�ڬܷe�q� [u��q�9�'PC���]v�V�1:��s���l@�5\��v�V�/5<�������������lct��qG6ӟ����%qm�����j2ry1d|V6lr;mZ��V0]�\[:��Ż �m$(-��s�-Ale x[t��m%�eEm�׭.Ո�)�^d�e�L�Te��nCb�����zx\� �Ѷ�q�<���q�;��η��9�2��L�g�4�J�(h�VF�H��(��Iӛy�7'�!ۂ�b燛�i�v�VR"=p;�iηN��Z�	�Y�J�ʝ��[*��	�p1��tg�.�iФ��K���%eU*�gk�jmXE���������T�!�)AX'����'���� <Uub�q�u^�-�В�RKh  *����[u�#��P�u�%X�Y� m�� ��8	2�Τ��lH  m�7Z�bmH4���v�]�%��GK��N]]gJ�ϐ��(��ێ��!V�=�Wg���:�T��\�öζ�����\uҜ䞻E��ў��ru�B�[��ʎ��)=i��Κ:[a������3]����wo{��_�ⴗ�Z<���I*�P-�]H7M`��GX�9��]ώy�jR��<���8}s
��ǹ��N��P�A:Dݙ�U^f^^��V��otO'X�i�h���e0r��MG!�//� �����V�I^<�>�\�`^U��ITmJ$�)9�:�x��/�>�\�a�j���w�w�jkT�(�I�jG�/�V�_{�3@O���������3��g~��Ǵ��Y��5���؇4�u�v�s�[.�H��4l�4�-q�c�ڮK�̮5�4���N�D}G��5��Ϟ������ND�nRy�RNw�����5�x59�@� ��#��x1Vc�}M*�>��:�u�QȔ�U"�Np�^=�x�1�����9�
��f4ڂԄ�:#�`j�J�����G@�Z�`~�Dr#����`Uۺ��Fe)��6�}s�M���� N�u�$P�sWv���N8yj%vV�i��d�j��,݇�sH�=N���WN�tMzk|�}�&�@��u�'I��=�َdu
A1��FԢI"���׎����;�l��� ���QR��&���Z�`z����"c��s�bi�������*��P�4��r�76�kQ��'�i�@M7���U�5V�X�<��F�$A$[��9�:�x����iw��l������F�!ԁֆ�6q��-�ՠ.dŵ�U����c���U\��ғAX:��~������X9�T���I� �otS���	PtG��w���j��ZH���l�y�}>�]s'۰�A8Dݝ�U]w���=���Z�`�gө�@N�u�z��Ͳ�TMɩ$[���}�}�Og;��n���ww�7�A���= �kU]���e.�3I%Q�(�H�� �}�������7_��jԳ~6��ɥ&��γ3�zv��*�v�N���u��@�Ku�^r7g:��3N�o<��WND�EM�`	�n�u'8i��=<���e^�JF��T��� ����2&��ө�jd�Z�g�O(�
�"Q�	I����� �����%�<���=o>[��ڎD�H�������t�7XޭS�r�o�%UXW��ӂԑtG�λ�|�I�)�ZotO(u�8��S���BK}D��  �U݃��uKt�D�3R�Yz@�����6��$H�ݸu-�knH  m��Ͷ��u��gY9'j���� �H巉�&�-�T���7F�9��m���{bIf���)�3��p��كl�)�/��v�W=�:�d��Y;7]�jm�;YN�r�����������M�.�®�3.f�wy�(&�U���Or�,�q��Y'a^�(1�x�qOpn�it�0��W]����t�~��y[������Nz@%�f��U~�2B������e:���RH���s�v}��3&­V� �ժz�9�L�`Bc��FԢI"����粂��f>ֵIy�Ű/ٙ��3SX��)EJM�M�`�7Z���sot?G�OR�`w+��|�
�JH�*sso�w��l�$�3����U�V ��]M;���ͬ[hl�d�	[tٲ��9��v��js�u=�/.�1����	[Q�G�h��r_�~�����yV�W�z�O@�]�F�r% "DI9�:�x��W��T$ I`%R�"��F!�m���>x���Y�	 D,��	h���߾$O���}X�IOC��If8�*�f(�U.NB*tG�����>�;ų�Ui/��q��S����J���"n�򪮻����O�Ӝ�otٟO'X�5���p��捲�TMɩ$[����\�`�7Z������uqu7��zt�T�Kr��k���EႹ����88�q�I��D�Np�^VΓu�>V�p\������ssM�U7u�<��V8�=��������ǹT�ˬ��)B�$C�9�����^v�$��w���P{BF$�D ��]�w�7]��;{���T����U�rw=�e-m� �O��;�|�w�`^���D�%*jn軽�=<�`Rn�u'89���8�ʶ�H�t��㔩Jm�� �&Wm�̜�67b�ӻK:ص]�M��<�6ZnTT�=���1���-��\����j�֏+Ϟ���W�#�n��Sz�^�{|�k��0D`����}���Y^���v�}Wme:���Wws�/ZK������U&� ���3(��t���CrNp�^=�w����$��gf��&�0P-B��w� �/SX��')R��5#�n� �Rs�>m���� �1�S����q�fy��v�m�see���)m�vsV3�8um���Rc��>��ƺ�s[����۷����otO'W��&�@]�mH�m�DE�3ٙ���ǲ�-�c��[�Fa/6��)SJFK��<�9��7Z�NpS-[{�����ӂҐ��5"�n� �;S��Y���Ӟ���n���"n���/+BԜ��{�y�s�5I��ѵ�����~w�ʥ@j�_-l�   moK/k��i�.�a��Pڪ(�g(���@�`�9��v���i�  Kn�2K�[��h�m]�zkֶ� YVp����~[�>��k�ƑY`���鸳�D{@�>���ܾ�ٮ��N�=�F�;i�m'��3܅t�<P5���⸇��t�˻c�i��.���;k�����pSmtN���w�ɲ�$f%�ֆ�=:vȪz��gû�ӯ��b��z�JHm�f��k�^dє�Q�&��w�-�����%��oُ�Am�-��E����FԢI	/t:NrfF�7Z�Npͽ���V���>���*B�T��&��R>ǟq��U)V9�6�@�� ��n	�%I�9��ͤ��^-����}����`}�>���S��M���H�H����t�� �&�@]I��G�~Qݧ�a��.Km�@B�#T�]�t�y�@�FӊGk��+�3�F��V-s��w��'8T��u'8���e{NJT#�M8-���1�_4��(��(eH�Ȁ5
����B!���Q	AUVc��C�WsY|�jI�}�w�;��l_�1���JCzm��;}I� ���t��s�5\�ށ�Ct���5*6�Ԓ-��y���x�[��}]X�����,�$"6�H]�`*�=�9�� �����Vs�}��U|�>I����i���T��ކ��f��9t]��S�xcZ]G�5F8ϞtڤJu)7I��i,�N~w�`e�{�y�s�j��7ėw%]�M�f����.ot:Np<ӽ�������6�J6�R �쿾� �_;Z�R�k=�y\��!5��SeY�����H�z	yXF]�����6_1߄���l�� �a Z��h𔄳B4zEBh`H!��=�4eW�ߵ�JpPЁ@(*z���:�Ch�^���GG`��@�H� [8�-<רyh(Ep	�U���ܓ��Ű2��M��JTґ�Np�[��Xz�N	s{��r:��'�.����p-��;��rA$���x�v�m�jRjF�8:u��ES���k�� 5��ZZv�a���s�]\�<Ψ'H��>���˭u'8I��<�b��-�;��h�)�R�5$�`6��Γ��j��r�tLt��ڌQ�I9�;��lY�����\�y���5)�ڤJu)7I��-��;��p�{�"#�舀".� H"�Ct�*�`Qc $D�Ш��uZ�l�ӏk	B%I��q��[�k3����řoU$v����-����t�3�������jM<���q�\��g��n.({\�@iȒ���
C`fg�s�{���-�v�����ڎD�M)$�@U�z㜉��j���O@�ֳ~t���h��ത#�MH����w֌%���I����.�t��3ꪜ���+f �ot:Np-��9ڻ�M����5������ �Rs��\�� \���z� "	��b�� ��J��]T��"@��$�l   6ٷ:�I8�o+���h�&@-���i7  A�H+v�:��6ĀUUT�챈6A�A�틻v�t�[,�R��:��n=\��vi2��[�����"P�����9�uŃ�2�nv�nN�N�Y���\��؂^Z�Z��w[z��N���~��t��}�틱2/2}��i6
i���̣�Ca@��j�M�\��]A����.e�.l�du::��݂;cQ�n-�X��W�c6x1�.�Z����~:�� r����G�G-����1�H��Rn�qo��!fm���v{�-�3������U��R���wZ�l�M��9��� އ�iȒ���E�.�3�<��Şǰ/�ֶ��Sj9�4�e�����[��ڼz�N����������_�p�I����HF��H	J���;è'�h�AfsI�V�œJ6ZR�b�lY���/�ֶ߳9��Z�����|�r��.��鶶�������B��T�5<��}��'y}Ű1f[�ڭj�;��N�$RjIs�M��S���9̪R��]}[��/�Yx:"6�HI9��UZ����-���{���By��}�/�&�*S�I�MŰ1g��w�́w��p�Y���[i�Z#��A�����T��s@!�ۭW=��ΰ&�c�6�T�9騥
��H�'��_�a�.����w����>__�`w)�`&ԈQ7�
�0���Γ���X{��V�IY��ڎD�JB��Np|��ԓ����+B��5D ׷�ɩ'�r�s��1�pZRӦ�[���/���X�l�_���I����.�t������'.��ـ$��Γ�`b�c�H�A��=17M(�b�娕�Z��6Kf��c��z5��9��n��c��M	�5����3����Ş��_�a�3�a��H��D��0�j��G#�����]}������3�jS1���%&�7�Şǰ;�h���@�� ��n	�*�ڻ�r� �7��'89�}A�	 H!*B$b(w�e�A&��/RO|/ӒU�fT���*�*��&�@�� r����`w�E��5D�*�N���n��-��N�����$�&7=U���&�J��%Np�[{��},�~�� ++��pZRӦ�[s��֌�k�t���ANK��"j�>�2�+@\��\�����՟-����{�;e�N�$Rj9�	w�lϝ'8��X�#�r�`�B3�Щ�(�BI��w�dK�O]`{mw�f-DA	s.]��m�%����  UJ�;�����lm��Wu� �����
 �#�볩m�6Ā  �۶��1�T��-�����muUU]@�luغr��=��\v��mt�5`��,I;�bP���S��.v9�w�n�+'���sq��\q]�ݬnW�nkp��:�;s��r+<���[���u�v������\
��s�{��w�M+�i.|�39�0�V��i�6s��5�qn�E�N]�v���ӥ��f��i�Rn�qX��?��a��Z�w�8fs�g����*��P�B1I�#��`	s{�L�s�9mV�+��Mܓu6U�Uـr{�y�s�9mVm#���a*���ڎD�JD��w���ۜe�X{��M����?B�>m8-'*:tӋ`qf[������9�;�1l�{�*��#�m�t�sq��Y'e^��c(�n�C���3���s�J�1y*D`�Rr�Lksq���l����ID�G#��[U���35�"��fB�0�̚�s����Ob��pa���7=�mW@��zw�L�`B�T]T�we���M�@R��G���ݴt���p���*B�JM�r-��1V�֌$���M� �t/��Sv]�w�WZJـ$��Λ�e�����N�U�J��[�m��2m�A����j8��d�<,�����hr!F��*�y��ǘ�1�/W��X]� W��ڎD�M)w{�zR�r���֌}��F{N$Rr�$���x���f���!���$ ~t�T��w�w��=���;wFb#����{������６`��ۜ�&��;�ZI��N�$)�����p�78�O(���UN���:���N�OQ�E���t]�"�1� ��3;��f�c�)v��}}m�_�s�k�� ��F���`|[��6�
J��\������,��+������W�R�I�	G8���h���f6�]>�@��s�>د�NDF�8��lw�g8q�-���;Z�>�y�"�HK(�x�4j�"�}���ԓ���'��e�R�4�d������ߦ|���6�ﳜ �e[Y$zIӧ�R�)�(@C�Rev�\���V��t�9li�H3�[6�$Sr$S��[������g �}��q���3�M�@����'���QQ=̝%l�;���t���9�=ۢ�4HSr����g8q�-��w�`{ޖlz���R#jTRB��;2���y�S�=�^��y���e�4V��(�7I�K`s���Z0�7��78� Q����+��=�=�#��}�%�#	Ѵ~� P)O1W[e^7%�G��UUJ�8H���	E��@�&�e$a!�R�� ���B��`X�=H�JJ4y��Q*��B�@=��dT��!!$a��G@b6i
��^�ه��E|�M��C�_��n���y]��㤝{�����e�   �  �     m� ��                    `��O+v1��k�#L�Ux���T�R'`��X)z�ں�V�A�M[Pt݄��3D�1)�[]�G���};�O��&��k$�U��u$� @
P`8>�H4R  d �� 	 8�� �  �   p (	e� � [\l-6�  �   [@  l     l         -� p ���ܱ��z�Vc� �� ��G[�-pH�}J�-�����PK�x��f�ں,�W�Z��K�k`�}��t�M�$ �c�� )@A���u�2'T�����N<��#`P�H�M��G��e��X�e��|ݍO�v(@�y�	��	��Z��@�M�rW$Y!���'6� �$�y�쵇��4��p�����wǾ�ܚS���VC4�d������TnC��c�8U��"��<��<���x2;k\��W��/<nڝ�<\��݌�6�[Z��ƵD�l	);.}q�4<�^[�e���۴^�:�۔"%U����v'�L�0�%2agv1��M�YfS��m��=8מʞ������*i؆�<n]��[l������M��
���(�`sݲ�܄�7X]��8Šc�Ur�l���)��.��E���89n�u�Mw$�λ��N,��!�ݝm�s���i1�[[v�F�v�C�9i�p:!�����m-&����g��+�����k��O�Hk��X�;��'���:s���wm�q����Fl6�U\ŀt�FJl��V����HR��m�u+%촨 �灪���lbEB\=����x�/�rz|�9���"���"�A���mD_E�@�h/�wZu�o�/T����I9 F�܃i�   ��t�����a�*Ň���USj�r��khl4Yn�[v�ܐ  im��r�7mP#HZ8�z�i&��곒�:�>+�0<��!��/%)�������0��@��z�����t����v��s�c]�wMn!m�7��֎�
 �|�s�˰��//T:����ϛ<�v�0ћ�vj������ ���J���ѕ%��[fg�l�jV�6l���5Y��$7nr�k�������)I	�	���g��9�7��78�Np(�5w%�U�Uـw���s'U78�Np�K6����ڎD�M)$� �<Ű1V����O�s%̭]y��HqLT�Hc�"RN-���������g'wb�5�Q����'+t�K{���t='�K0|��:nzΓ��G��ڿrFb_mhl�ӧl��Z�χw��[\�g��ˎٌݙ�p�@3۞M[��ݚ���n��M������Jـ+���t��6梒Np��[]�翄G�
����֤���vjI�����j�2����AiB�Ct��`w�-�{ק@��k0������B��q���-HH(�\]ֵ�V��o�`_��������U�^�g�`{)�`&Ԉ��T9����� �Ǳ�>䘦�sޖlV�`�ƲETGN�N9J���^f�/>�Iy���m��ʮ���gN�#��"R����s�u^c��x�}�c���}�� Wk��q!�D�B��t���֌|��ғ��DD����@���	�W�*'������{��s�4�B-Ah`����^�U��?���V���I��[������B���m s�^s@����+��Ӡsw��;��2�dDmJ�JNNp��{�w�`sޖn�#���+�Z,Ę�F���i!8�Rkz�m�f�s�$e�:.Ƹy��:>j�}�(-(Q(n�q�u�-��zY�9�Տ���Pl�u����7$�v]syW8۶���L���y�zRu�3�Էąu��6�DN���lw/9�=):�7Ԝ��h�:<�8�����SJJ�Np1y�m���/'�-�۹����ȀQ! b�@�P����h
T���{�$<����uyU.IJ�`s��lڪ�������8U�=��UUU{�|��5)5#A�=!dU:��V�k6��EN��m��q�.�S(�LJNV�S������9ܼ� �ǝ����iK�ulz�$��M܈������G��{��x�=�f����x:HDt9Q�I���I����U^J��7�=͐\S��AiB�%I#���[���`s�y��w�cK:z�X�$!�F(�Z%l�#|��ғ�}I�삯�ON�~>Mm�^��m�  �[���[:s�3vmd�8�jՒ�`�Al��6�828�6�B��i�l $l�M�z��P+7D�e�x���@8ʳ�*k���l�H�U�$�76�2�;p<�sS��i%���zZ�I�'I��MOj��ؗ9�A��&�h��FT�m?��R��
|���vdǀ��Tu�
fl�+֝����ޝ��QQ�[�0�盙��K�vi�ړMڮ5��.��<�.({]s��Q��T9�����s�	]��s������6׳���QȔ��%G'8e'Y�&����Z0�Ow>��B>\b1��C$�%
G�;��[��ݜ�i��I�栗#�	�&�2(��̝�[0�OtJN���}�C��ϖ���$���B��p���~����uW@q�Z�8۶����)���&�+�c���+\ʱ���KE��Ɨ�S�Fre�3۳U��͞�st�n�3�I���� ��Dl��/���/��+�* rT�=�޻Ž���T)���}���ߎ��'�Ӻ��/�F�)Ir�G� ���`s�����/,��[�y����Xn�R"'PqQWf����A�M��Rs���֌�.�xM��JjiIQ���y�`}Z����=�h��K0Z����L\��kCg�����d���[�-rܗ.��ۘ�e�.N9y4�uX�a��o���l�=�h�;ͽ�=)���9PN�5q�EMNa�rV����қ�������ZI��N�$)�I!�=���$��ާ���O ��]k�ύ�ys�}���t*Dc����0?O�7]�m��{�� �=Y�_��V(-(Q(rT�=����`}^��0�o0�R���@�T����fs��N�J8�&�u`�۳�^����a��d�p�j)Ir�D�pz�a�=�K0�R��r#'fu�gё!�0�&�CN��*���}���W��w=�6=�f��V�2�QȔ��*��tJn����f��F�m�wPt�6�q!�A�a�Uj�T��s_MMU{�gf�'=��������� )"ĂZ����Wߵ�ԓ��}����I��1����z�a�=������6��
?V���dNH�ļ�ӎZ�]�z�Q�\s]�J�c�v��sL�� '��I�E:h���$����tɻ�<�ف����䱘��
�!����o0�����,��fs�_��V(-(Q(rB9x�[0ɟwZ0�=�&� ~:�X�$Rr�D�빆��s3� ��M���lߪ�t����8����{�`"'ɻ�<���>��N����r�Uͼ�����I)$���   6ٶ������t�WUc4v��V�
ѳ m�� ��8	2�Τ��lH UT���zآ^�o\%�v��r��B-e�;Go<�BF48^֋c�lh�bn��i��8�T��lu�p�׍��rrצ�sm�箽����|_��0�S��5iq�ўÑ�șsA&��ȁ��C��%a��뼪<D⽖|��.�YteKɒ��M�l�8%m��"ŵh�l� ���m�pO�j��26�Qȓ�T���g��`w:ـ{�рw�{��#������$����<�ـ{�рw�{�M��Fe�YLq9[�4��\�s���� �N��?}��ߕ�3�H�Nfr�E6�Hlw��p��M����`sޖl�^�H�(����� �N�>�`�h�;ͽ�2?$d�ڿ�����瞨öZ���X��;�̽��]j�Yv�8���:Xt�K�0.����# ��F��f2Or�t�^�R�I�6)�8m.��6�k\5��<��"�9�������u�8��;��o��T�;Yu��MH�SVE\�Wg@ߛy�n��/Z:{���"��a�ڎD����$��{3/ ��f�֌��� ���MZC$� )&��za�>�Wn�� �}���n�V��Omd��$�Ӎ�)Ryn�Nʽm(�r�v*]�n���rk���]���ڔ�0uƤj�M���p��6��Y� v�&��ze����F�	
�wf�m�y'x�[0��F}���ЩD��JNNp�y6s����(W2Uw��� �h�6hMw���!
�%JIA+����RB� �tm7�x/���I\2T������%%0���> ��4����
Ƥ���w�*�o�E��b����D�WCE1���aE��!&���Ֆ�00#�i�ȉ��$�h�o%1�������o�d
℩@�zx�(%�a�yY�Y�!*ƪ4U%�=G�,�>��9�-+E$�Cׄ+{�D��-���\���� ��e"�ڄ��B����KCTګ�>l='�Ї��h�\
CI �@�7(8�.���&g�3�v�=���P=F�؊<U�v������i����8~>Ñ�Y����o2 ZV�
l�M�\we���v��֌�i�y��:z�X�$Rr�7'6p��6>�O�ͻ�7�ـ%J�������<�'�V�W6V]ubk#v��؎ҡ̝g���T�v�[\%��1�[����,�����~�Dd��mX����9EINI� w/&��ra�=�K6{���H++��q!�A&��|��z���}�a�&�w��8�M\dUI5�h����|�/�$��}��6<�I@�.�"I(��׫UZ�U]r~Λ�}��j��B.���� =�����w�o��0�]���USUZ�~��r9�L�N�N��*��Jۅ�%t=����9���\����f�����GQ�I�� _����L0�Z� =�h�pC�'���컻�|+GY!��G@��� >Z�`gOVk��NA:QG�p��6_'����hݐ�Ѓ"jn䨛���*���RO3t�;�L��l�����`{�M��JJ	)�9��w�F��0�\# ��{�T�j�������m	-�:�   m����z�o������6���v�� �ILmmlD�ۇR۶��  ��c]*�[�[M������l�\[� d$r��׋7NY��8��Մv��@Q++Vwcr���۳θ��6�h�K��'�'�ogv�w�ûm4U��g'n�tp��oAgmX�F�a����f6��g&]�+κ��ݶ�>��=������I�S�<�7\��$��N���ۮd�F�C�֎�kJ�v�7n8��`$I8fO��"�sf��^s���s��Pi�@�P'₣�j�U$�a�1%��;�{�i��v�s��BG}x�ڃ�����RC`]��s�Z������}����}
Q9Q3]\�WQ5w����v��֌ɝ�����X���
%HI&��rـw�р�^�i��l��rv�5��3�6C�-z�l��I��k�r�7r8�mՆk�T��}c�Xxd~�����l�7�=�4� �+f�:dI%'� r�G;���~�Z��~�Mw���"@y�o�'���=��N��f�M�ND�FI9�1y^M�Wnfѵ���K�����s�:�<�q�T��IE�Ėwx�jp�Z0sOt=3-;��8�M\dML�fN��[0��4�@<ӼU58�UJ�f_mhl�ӧl��Z�χ-7�.g��l�v�q���8�2�%,�^պ��}~�r���@<ӼU5/d+f�,��*DqS�Np�y7j������},��^rs�G�?����(�9!$��z}�`_�Y���*���W(Ѫ�W">;��� &��>��qM�1%]�D���N��[0i=��4�������1le]`n�%'
q����9�v'��*Jz>���@w�C�twi�f㋒�`PxA�L�ݬ���[q�0u�Znl2�u���;j�Zt�q /ߝ��)ݐ�F�'�����j�&�'&ë�/k`{ޖli=�6����\PTi5q�53Y�:JـsI�y�x�Jp�ֶڃ��$*I��A��p���I7��+R8+�@���7�t�%* N����UN���+�*e�2��꫽�6� �IN�֌�Oy@bLo#TSm4��J��J���l�4s��9�i4��p���c;l�pl=�,}6ApUݗWx�Jp�`�{�@{3s`gOVk�R#���jَdT�� 6��IN�7H���q���j���$���g��]��-�ws�ϋ�M��JJ	qww��8�U��@�S�>�^��us����Ӊ5R��I�� �;��]h�9��@S�� ���#��ҭ����ݽ�&�   T��m�v��� :\�i���Jr�[[hd��,��l-�m8  F��٫e�0I4Ů,<&��6�����9��]5�����Si��`v��WK6yn���ts�I��Īv�]ѣ]�>�#���2�:ݸr����ϐ�HvC�FL��v0��b�q��]v6��>@��5u�^���9�η�?^�������TkF���yӭ������N�F��͎�k�n�L��/k`Mv�%���A���b�)�����&���������/2�8��f<���{=x�ڃ��$*I�`	��`<�`W*�<�рoG��T��R8�ܜ����+����֌6���pC�'���˛��K��K�����:��0q�[���l>9�&$����&�Xym��&��O7X�ʰ�ʣ.n�~'ϝfg<ևl
Sc;4��jLT�K��ԙ�1qC�띮4����o�o����� �<���X�S֌X���r(�"J�Np�ُ��V��z�֨?)�E�$	H�$Y$BE�EB	�TQ$BD$ *���S'U'8��� ��T������W3WX�ʰ��p�{�9�ǳ�fQ2�S\��MI�����' M���n�6]+U�/r���*
�.Ȼ�.��jZ� ���k�`r��������E���4St�M�pښ%b��V2(��sv�,��	re�=�5^)�(ҤF�B�i99�����~U�B��8m=���6O�`\M]�7u�9\� ]\� M��I�� Ξ��)B�Jn���n�l
����n�T@�E)����$�s��w^��#D��N*$�a���>� s��@R���|��9��O@��P8�Qȣ��)�9�H�s�Ş��?�Z˙�qg��8Pv����U�D�;<�v��$�zR`+Y���8ѹ�g�r�6�M�FӉ5R��8�,���~v� I����`@�K�
�*�2*��3+@j����"M��Su�yӸ��U�V�3׋m�:��I�[3�����`_*�-u��{�҉t�"S�rM7'8{UUZL�o`|��{�s��+RV�wH�
G�H�[�,iH�4�^h@X���p���J)9�{z��ȶ������z�`Su�3Cgjk�=��:��y�����D�dz��\yΔ�����������^��ƹm�}��s2���r��Su�9榰���t��)=&�n-�w���ԑ>y�χ�������;��9��)��9H�w{�29M� �X�Jp�{�ux�U*iĜ{�����^=�������f�Dr"6�sm�@j�\PVUqت��{���S�""93U�O��s`�z��?���p"9�nG#� �"
������?��_��kB �6�isx��\� ��,  	P� E�TD�PތD4�@ �H�EBPF�A�҆h�Xh"�$H@E��Ȫ����(e�&�I E$EV�.�A7 PP�X*�(!"��"��
iC%*
:��A4� $�����*$@W*�DCg����'�d
�n���Dd dQB@Q��ò������?�������/����?���ݣ��_����������?�eW��̱@ �_��G���������?�O�� ��TA�@TQ���������	?���'�g ������A����������t?���������y��jB$%2C�������|��؇L���?���#�w�������(/�AТH�H"�H�"
@�H���)"
E�� 
A�����(�X"�H�*$b�E �B �H���X��*$ �)�)F
$ �F �Q�)D�) R*$AH��X�� 
D�)�����)�)"�E"�E 
D �DX��"�E ��)���) 
DX��`�D`
A��V*$T"
@X���H"�TH�� 
@�) ��� 
D �)B �A(�Ab�@U�)T�)  �@`
EP"�D"
EA�� *$"
E��*$ �� 
@H����"�E� ��)H��`�@A 
E`
Eb
D�) ����F �A����`
H�� �) 
DH��$(E`�! �	`�!H$P�Ab� �H� �U�H$T`��ER)"P�@�H��EX	"T�E(DX� �$�A`�) $ �DH�"BAH$A"$$U`$ `�@�F	 $! � ��(B!!�!"@�@�"�� X�H� �RD $D���,�����EE�� ��� H�� B D���*�LIRQ$I RAQ$I �ED��H��H� RR���_��h�������O DU\E�@P�P�����!� a?�������?���Q����A (?�?���6o�������?�����g����C?��A 9�����|p�����@�A ?�ȋ����.��� �cg�Z�  z���~�D�cL<-�1�
��<�G������l@�A !�m�O�����g�PD ���AZ�}�_�� ��6�������a�/��-"" ��'����@ ��� �/���8;	��a���3<OO�4����s�z�ρI�?�j���T�����@����o����$L3�����o��?̇��U���H�a�* ����F�����������?����g����PVI��@�!��P`�` ������\��QB�  @     (  
( �  y(      )!D(�B RR��*�PR�*�E	%E@(A%P(
�$@A (�S    � �(�  �Q�ϥ2t�|�}n�2j���,g����q�wh�&� ��(�`b5�  Yq�vne� ���<Q�c�0�gJQ�� �P`�z�v�;�]� �� *(P  �m �p�=��SM� 14 <8 �Jq)�Ί � L@Ҕp�����ce   R�h� ����()� iLl�bh�Y()n@Ps�)KJbi@�t��PÈ$    )+ Δ��4�ǚ�N,��>�]��犳}�u�y�9���K}nON�*��Q�����Ͼ ����g�g���@��.�z��ζ�ۗ��ܳ�� �>3��{�y��>���祿�K� ��  
  2O>�����O'\�>��1�N� -����|�=�u���ʩ�қ���Yq|�y�cx�����=��}g W=I�����ɯ^[ŕ������������μ�]�/ ���  � (�Y@#�2}'qw>��\����/� �����w����M��=�w���)\�u��� .�ϱ���ʗ�
�Q�{�_O�,�rk�O�[��μ��w��'^�>Ou�[����    ��jF�J�4 2
�������Rh 0�<z�T5  ��UI�J� �?�%�)R� D�5%@� x�R������J��������W���fO�J�U*�~���(���@AU?�EU�EU�QU�������p�X*��$�5bP"!	���$���P�`�		KD F�!H��D�0�U�c������g�����Ns�^���;v�^����y�b��@4x��
$�H,Bឞ��)���8�0�P��A�`��q`��@A*�
���<k��/3<^���磿W�fx�
j�o��[\U�vr�y�_�'�ը���.!2��Ex�����W���rb�m�xg���HƤ�¬.<H0H�[8�����٣�L3NÆ�%4kg �q�o���p�i����4az��jH�"��_}ֽ�4�(f�kz�bU�熷���)IxL0�H���Ħr5#����1ƙ��:"�4T���
c$+�@b$0�ΈNM^kI�R�:���}�^@���"�^J��sڨsA��<!����߸�	�`K<�O�9��,H`A�M%b���/�`,1�lJ��\ug�
�l�1XP¦2!	 �瀪ه��������jB��ݢ� SI	&��}�Z-v�]�o��;,BB���`��@!��Sq��P����i���o�Á��Z�!�x\�4k���z0�!7���C�]i$R��4XVīE1>��FG ��MŀC0��"�N Cg�2IS4h&��c5�Z!�ω��./{(��T5v��!��s#K��w͞�`{&��W��M��3	G{K��}BP��!$��l �bB�H�����4M$�t��A�#���0�"�{�.x{�ʤR�ܔL��k��8�$&���r���ŋ��G���\4�p���]o��<��=|�0���0�^{Bj��A{�W}�Z=O���HEv��$@��E��0���6(,��_�����������75��3�8xa��]��ō04�Y\��,iq�nk3�n�9n�.k�R���=C�i��)�(a��%#}LF׌
�h6q��#L&�O�]�!LtȅpѳK8iѳ�湰�ȪG��"��Ir2�fg���a]��0�Rl���=f��xy�@�"�I��B"��ka�H�
��W�P�k����z&�$`D"]z|CY&�4x��z���`@�PH���
�M;x	f����i����@$�N�6M �j͓�������/��\��S6�!�3Fr]����� � i6 U�y��P)��P6��� U�R)@�)DH��6s羚/�S�sd��ןx�0x���"p�pw�5�y�_t]^pLcH�1����Ѡ���<RI����㥅�Z���!L16���V4��縧�Jr��'%��J��:�!ں��3����3[y�_&���%1��5�^�B�����S0�{�X�`¤+�B�B�}�<� G���5���������� �
a��K��96A��C0��F�		���b\���Յ3[H�v:=aq�6�p�4-'��{ٚ xs���g	甅=��HĀF	���X�'G�M@�ѧA�!$ �ۦ53s[	�@`ā
q�B �7"W#\��{�3����)���������%7$l#������GN�<|	44���Ē��0��M�9��0.:�<>ύ�M�>����LM&�P���	e.k���0=}	L�3�Cs@b]�9�C��p��.�����H��Q��f�H��kg2/�3Þ�qb@��%���S4�V%�q"Q����q��}�s�'=��k{ݒ;v���!SH�,��[�j�3P���W^y�zqk�p�����K$1�{$���S���*�ٮ|��<�5!
c��l᷇��z@����<�I�4l�a��< �Lt;? �l��1d�S�%����Cf�{�}�g�Y��xg%��!�8����
�jk4�%3Z]�V�ōV@�)��
"�!	 �B@�@��H1��HA,��Q�`PƱ+�E�F� h�+���dq�i�.aZ�,��0����6�I�h�N�H�ɱ�\+h��h��
jK)%��
�ڄ��C~�#�ԍ3���߷3o�����f�@�g�.�D�0��*+�k�\�?HF��%qw �D�8��vh�|$)�Ӵ�C d"�"G��N��)��5��o�xp#7F��|��O~�*J�v'�xN��ҵ���"� ��JD�M����p��a!S5q��xdu�m�6sV{)���`H��zf�����D�
av��H�ޡ���z��L�Û�^l�V�*Y��|���ѨCHXzS�1&�B��.]�ؽ�����3�_M�JR$|}=w}��B�*dJ�(m�$c��[9��OCD6��ka�g�!F$H5�=�����B-LX�8P�_��nza�K.h���p5�� ��
a���x�_9���p���ӛ�O}%�K���{��w�^.l#H�,�#B�V%IA���X��D�"�ap���{��9��z���r��laaa�,M (eP'�aM�@��(l|.+�g�<a��;�P�!�$`R#V*l�l�ղ
�.��p�W0֣@�Қ�0�rB����� �,�����a$7$��Ah�$U��q%q�ˇ�����bsx|[>Zc�=)�F%!R��+��)ű+��K��x��B,A���5o&C`P�;M�@
AZ��r5��;A A���� ��CJA(�h��+C�p5��kY�ڈ����H7u�9N}YBV��o=�	C��4�8n��q�~<x�d+�F�
I���=ȗ�Gv��$k�h`�"xE.�ia��C09��C^�7�l�//��ǟ<	0lT����y����֮��[����b����	#H�!���<!I} ��N����0��g/��֍��{���_Bd�.�b�n��*Ji&�%!�)9��{VJ��75���Bf�p�{�6�2+���<#H�#E����h��X����K� Ț�{�6O.��w����Q��.{���+H^�t�1�$�� �х��h����C�z.�$��Ձ��2E��=����d���aP�E=b@ap�n�\��Xo�p<�g�@��
U��GL
e5�l�Y2��X���H@�7����za�J�p<	sDa0׼��,k��H�H��$��˭���I�+���peL�ӲS4H�5��J�p�y�l�L��Vx��	�S	BY��_���|[����f�`��0\�Xl��
I	���"�F��%#V$$=���ys�N{�&H�e��уHzh�j]2$���)�D���M1�n]o���6p=�za�zk��WG�sF����v�ﯺ{�s��o�ߟ�                   l                                	                          mf�j���[�G��6���X;l#m� m����5�`    -��kX�]��i $2�f�6�d�� m q�� H �[�6��-�Н49�/kqa�7mF�G\�F��r6� �$��J�"]0���l����7m��櫃���^Z�jU���(�ન	g,�kM&�m� ���m�8H�ͪ���ٶ�mr��J���P�   m�dU�v  ��4RںM��q IJ t�8xId���,�HK(sZݹ-'��                                  [@                                m�                    ?�                 Uv�                       ��         �                                �-�                  ���π                        	                                         � -�                     �|    ��#�k���׮��FX��,���jU������]� *md���ɺ�l��  	hI�@UT�v�RB-�ݶB�)�lU�mNP��5Յ��f�m   �l�`�����[��N�k�Ä�n�m�ͪ�a���� �Ue9t/N�v��fBP�Xaa& lYפkX  i$s�u$l(  Smulŗ���G6��"^T#���mSR�c��;2�q2�ɮ�ں�U�r�+�\��rd���m^�8ڱ6�6 ��F�����ʀ�R�����(.]�����N깕U^^@�*��U��%�l�  [[-��y�YUZ��3ª)����� �U*�HMU� VQ��� R�km��oP��%M�p�o/�59�IP�,5T���\��5*�P��幪U�`b��� ���VʵJ��0U��@P �m�`[@�M�zp��m��7l�Im�����b[@S�m���m�@�u�ɉ kk�9�`�k��$� ����`��66�I��v�:kr[M�m��q!�6��  $4i�ٶ[d��@I�Xն����b��{!��J�`Imԯ�'I$���V�nl�l���l	sAt���UҭXv�*�U�9]<y��мP;K;&�ٶ���>m�wu�U�]l�
vA	:�;�-��.�P4��U�XI�v�]U��& ���؛Y۱ �0,״�oZ� �m�l[]����8*6�V�)-UJ��@uR����YM�ip�C�N����6�ci�@p��69m �-��oE2��6����-��  ��H%UP)]��jU����y��m��.î�
*�d���m#�^�B�n��yjU��;m���bB�8{j��An�jjwq�@Uen��rö��=mm��@��ʢU�n�S�Yy+` �3��j��C4�@uj��̄<Ocb�L�W/l��sWU m�K��]ߪWΐ:���$�&�]b�%$٢���m��8�`L�*��A0�jU�a�UF�Z�����m���"O:��9��k-[�	 $���{հHm� ^luUև��Ғ��+�vmp �4�%�֜���d��BiUV�Z:�m�@-���A��g��X�`+�� �/F�	}��m� mU*=6$:�p�;;@L6��[��l�R� �i���5�-���@ m"���Z6���OHi�Xv�·)-��m��$8�x8H 3��ai�H�vm& �l��9:87m�lp  v�%�m��
�y�H�ϟ_�7@ p$�so��� V�p8	e'M���g���(t[[����[`  6�@ѓa��H��8�`X`&�m�	86VTHz�+�T�] ��[�n�����K$��������Uy
%�:݉�-`;�v[R�ml�����c���a�66��%�v8.͑��y����%�`�1s�vt�F{Fz�#ź܌�t��=j�T��l=h�;Zzxʹ���Ŷ����w�o� ְ ln�#�}z���6݀k�������U]R�:��P��9�B۶jٶ���Wb��.� ����Msu�,ր[d$ 
�U;75UUm*� 	Ym��M[R촸�mSe�-�ٶ �m�-���[%8Ѷ�l �N�hm�	9�M&�d���ձ�I��Ipmm��m���l�K)MsfKh ��&����   �i$ �m�n�-@ut�]�[��؝-�-�U�U�h�*��M�86�-�q7k�ѭ� mXe�ֳm������|��� 2�A�-P�@UÞ@����j۶�F�X�p �m t��H�[K�����@H�e�Z8 ���)�5�K��R��7�J��r� ��j���� s�	-2:�[��l۶�[h��$ન����2�R 
�$�vv�z�\�y�-�(8  �۶�[��VW�]�j�ɀj�Ȓ�[@ Hdm���]6�����#���6Λ]���M\��s�FJ����Bn�t�a�:�_2b�[[.�Q����wf��p�r��u=#��T�'�;��nuk�����܋*�·Rc�qus�s��If�ܠ�W,�� ����FE����]U^v{i.�1���j�pKq.�ڃ���@��&�m��=UT��k%M#@��{vH!�Ul�=D$�S����V�����vG�xtv�Ԫ3J��mUU�U>'tU[�
܇Q  �6� -��m�7t��z'j�g@���8 -� [Am ��n�e�r�`	�pzk�F��-�3��m�@��H��=�U2�Ҡ@U�U�h�e   ݰ-�6��$I�:���\R;v���J���۶�	 6Z�uUT�R]�MȷXl��Ѷ�  �����m�m���m��> � ,�� m�n 6}�����n���I�� �@ k��$-���u��۫g6�ɕ�z�y��'�X���v��tݕ�Yy&�"��.���@�].�m �88<[��[@����h�m�HmU��`��ÜN�5��^q�n�s��6ݒ [$����$�4Plej�W�x-�6����n�uY�{��m��@ r��R�g�+�X&�X�Ҁ���ԒG��*m�����ul��H,s���H��{\�`8,��|OM��hd�I�{t�N�@ kX����^��jL�	:�l��H����cZ�z���a٭۳L�+UR��ت���<%��u�"ҝ���+�{O��l�$7m���n����$q���V�l�SĀ[@�j;]���ul ���~�|:��m� 6�q��0N� �6�0zt�8�-�j�V6���.�a�]����&����GUQ�0�������@٤�f�$d�H[@`n�   �[���cm� ��m&Ŵm� [V�hҰ%%��    mU��u���Ŧm�cax)W@�]T�-��c"��\v�4� ڮ���XP��e��V����wπl�
�*��1P��nq���UJ���X�hmڪ�mJ��K��a����[!o@�ްn� �J�m�! �`�a@if��n�6�L��׳Y��im6�0�m��(��׮ٶ%�       (6Zh�mq ���T�m[[[l&�@  �`  m���JUV�*cR��6�[e�=mh� ,0[@ /Z��  lm�  �(f�]j�2�#٪��', !+R�Z���
Z�`-�� 9�l�   �j��� 8    �pm���Ͱ  �m&p �jYm�e�%^�]�:������4���l�I͖�F�%H��$S^�A �����*���!�����q��1x ����	�*��>�A��"�OTP�_P`��� lTM)� ���Q�OS�Q�a2db�H���X,�H�PD�v��0}D��ȣ�/�@��v(	�(�@��S�*D$&�T|@��$�"(x��DHz!����)LU}�1��� t���Q����b��Ox
�(�� �	�� "��P�D��P� ⫐@X��ڕ}DH�z�Ą�$)X$(� E D�$!$b���I�A�<RHDX� � D�#��M"1	+�@aH��R� �B�q|J���H�X0�",���D��`!���$ؤdEX'�,$ ��I�$��D
�A,A� ����S�%�GK$�O~6����pT�ҁS� ��
z!�U<T�>C�=U�U���O@9V���Qb!���E�b|,ؾ�lSk@0Wh�����EhU <D4�ч�����?
���F(������^�ֵ�              lӖ��kM�-����#L�����{��3٬��ʩ�! qs`�P�d�Lۋ՛D���`            �   �   �h    �:6���     ��  �    �6�      $�   ��г��t�G8HK6,��"�HS�X��+:MY8yCv�n(�K{&f̓��;�(ae�n����N�T�9^���5�[N�$��� ������"�KUWmK+<]�\�9@y]����X��
d����ݪ�Z��rnK��X�v�5��6�����!v���\F;V�.��R���+maFОݵ͜v8"�lH���;M���ĉ����F��Y`�G�,�E�!��͡�W<@l�H�nΝ�nn(u]�ڧ9���mm�B �S�������״�h� r>�[U�\k��Hc��ӣ%���&"o]�ˇ��y7%Sw<9�n����d��h6[����r�[���V;lt�ģ�s�6��"t�"m�-�v�Y9[�.(0�T�8�ւ�	U�;xV8�U�m�ۮ�BV�j���t��W]V��B�:��kʓ�i�sv�]gN9����
n�������g�q؍��b㠎��\�Z�`MO��g��]��m�2n6�r��4l���\檕y�v�TyY�C�AV�^���4�g)*���Mˑ�	5��2��*ط:{�����hy�)�޽�]��zzT��]�[7<��Ǡ9sm��סV5c�E�G���)��tc���u8N��l�Su��[vTh�[ͪz��
k(�q�YH'R����Q�j5�!;\�;4�=�x�N�M����Y#������œT��E�Zmjj����ƥUU*��uC\�ĠX6�d��޶���M#8I�Z�T(QCI��T�:��>�C�	�6���{����{���>ߢ@ �[���N�t�Z`i  m��g�V�m��p _Z�w�bM��;�vdLO�x����w`�iη���{aM��K��i�,0w=P�u9ϴp�	�-�R���d.��l��n�S��L�"ħg$I4���6�v$W�]V֑��nA�v�n'S��^��a�<��WF�r���9`�,���'kSZ�]a�շjd��⁥�(�?8;� �p<��v��E{)�Ô���yPp�������n<���M�|@=��ހw�f��|�
��)�5!�2bh����4�@�%#�,F�`H�uv���f�岚��=Ş�w$�_��'蜻��4�@d��#kw�{�Y�L���%�4��<�S@�ҚWkz}�h׋����%PK�U탵n�z�뗷�ut�[�M�tl�sP��q�����B�4�)�uv���f�岚��p���,�E�k33SrO~Ͼ������D�s�@�Y��<���^�M�\w�q�L��$o@/���e4��_[>4����nW�c�	����$�<�S@������އ٘��~��:��8XFF�4�Jh]�����<�S@<��tocQ1��9�Z�s��/]�&[nH�^����iN�6fX�=@�,n$�FF�Wkz}�4-��/�)�{��,w�ca?D��@�h.&����#kw�g�,�&Dc"�dM94-��/�)��R�T����;�y�| ��' 3:��AD�Pn���T��9� ͽ�z}�4-��<��6�1d�(�]]�F��@�h.&��������׷ޞ�K*�-f���ݙ0E��9�B)�k3tВ�Z%+�����<�fwY�½Y�w�G4�@zbh���^�_�L&�Q6����hLM6�z �s@��W⚫��a��/���:�[����u�h����<�!A֖#��iŠF��@�>\M߷ߩ�Z�'��㱯�q�����@��M��ZWkzW��D����]�M��E�si*��f賻Y�uz�4�t��v��2�$�1ɑȢYNM�e4�h_V����~����9��{aUxhZց�ހ29�|̦��w\1���&E��"�:���#������T}o����_�2q� ��h^��/�ՠu}[�/�+����j&ԓ@������h���G4Lp3332�j�qZ{W=�+eN���Āh 6�6 )D�8 ^�Ѻb��U�.�h�q����Akq���w	�qtۨ�x�;�b��܏e������5�v�P㲤�q��<��g����p���s:�6��#����vi��N�XY��Ʊ�����õ���m��(#��ۄ��d����w����U�R�	�{�����w��_�]*�8})k����E���mϞ�nob�:���x�4��qC؁��Gi���m�~��Zmn������>�EakK�d`4��:�[��f�岚�ڷ�#���?�_��	�'���������6�z����L�fEȚrh[)�_]�@��o@/u�o,t�!�2L�A'�Z�#kw��h.&�+�^�zL++.1�Z�����l�j���Oj���1�9��l��D�ˣ���]�]�:iH�����Y�yl�߳�g�}�U�؇���,RF��Y�(@�Q!Jڱ'�C2��g��?��[<4�ՠuv��_nW�c�	� 86����h�j�:�[��f��|�
��L����p6��f����w��rp3&΢��20qh]���@��M��Z��KBR76��[��N;V�#���U���r�x�[�I�9�'�F�1��N7��������6�z����V{(��D�&����h��h]����9�UISa����\��"��w�����̻�U+^�*$3���<��hgu�[��E��&h]���������@�\}yE���V{
�feހ=�>\M鉠E��~m�?���9{V��C�М�<�]e
7fF�������%������ݮ���$�<�S@�������߿fg���4~u�_$�L����hLM6�z �s@�q4�Q��F�0S#���� �����hޔ�=�^��~c�'�oCUS{���=ݚp���UR������ ?����FwD�� ��i�%y�-I%l�?<I%zX�$�߿�>�L+$@s9aqjM�$D�8���I��� 9@�'��W<\<�ۚ���dp�Ē�����[�$��,Z�K�v�x�G����dXE���$�����$��bԒ^[��Ē�����\d����$I#�ĒW��RIyn��J�Z�J�l~x�U\˦����v䏍�I*W~����6����m�ə/�{UI+��l|m��ҧ��'�`E�dnC�J�RI[-��I^�-I%�O<I.���3-�]UU*�Jˋ��Ny�ڭ�����Z��   
Ut�i���U@�V��,vQ�.	6as���rm�������ÉlxD�i��o�eĜ���)���-V]�v�q��{��rƴr`ݿ�/_��ޞ�g�� 
�.�@��S��KW%{�+;&^�Č�gB�i��-�ιi#�t��kb�?n�w?8�X����YK�V��z�2��+^;���>>'?K&f
���s�<�=�:6�\RI{�?���ĒW��RIyn��J�RI{��1v;��L�r?<I%zX����Wv߻���or����d̗獤�w+�ȆdQ,��"Ԓ^[��Ē���ԒU�;<�$��bԒK˜��HʑAA���6����ɾ'��{v���$��,Z�K�n��H�9\1�̋��4�ũ$��vy�I+�ũ$���7Ē�.�RIs��cy��1:��5;�����Z�d{e�'H�+fuKiv+��7I���S_������6����x�yٜf�U��oo2�y�m��ۦ����v�'m��s<�*Y���zH��j5$�����$^���K�g'��<�,# ��<I+��5$�w��x�E�I�$��|�<I/z���~S"I�$����Ē/JMI%���y�I^�Q�$�Θb�v5�5LjG'�$�zRjI/o_3�J��� >��������w�\�$J��Y��3��^�,v��ۉ�c9k�j��K���#�̊dC2(�DӄԒ^޾g�$��u�J���<I"��ԒK��X�H��d2��x�W��jI*�;<�$���q�߹��y��T�]�}X�
�F���4�F����_��H�)5/�ĀH�;>�%h�`�)��E��˓ c&S1
����$I3(k1�%�eƫ��BI�\6!��1��0R�"��&�؆<��75�X�!��3V),v\bG�$��B'Ƽ<�`R��BT<י�q%�m#^XR��$��$�D��z0��TԎ,4jfJa��@�t0�,�I1 m<���"x�J0 �"bB�(Ƥ)����x��T!JĩHFh�
y���	�2�JM8��e�CBr�nc�˚�K��
��J1�#@�Ԃ:��Rl9�G�̀h&��Bf�2,�p����0�\�V"b �.�O"����@M��5�P�C�� (�h>P<�_W�#�������kw�9m�w]ݛ���:�q�1L�Q�'�$�k�[m�s|^x�yٜgz�����獷��n��j&��v�'m��g��oUv}���$�����Ē;�&��^���,)eS���;<^��:�7:�ZZL�Z��\˥�w7S�z[�vPz�[���������m����O<m���O�R_$����o�/<m�߆KW����	.K8�J���<��mω�$�����%��ߛi{�a���E��LjG'�$��|MI%���x�m��j5$�����Ē9�W2)��dQ,��	�/����$�]wvn�o������n�7?p]'`��UUUI_�o����j��Hʸ�./<m�{3��m���$���_z�fl���K���Ԓ��GdƔ�%J%�[�oM����n�B�5�v�r����g�]TDW������
�ģAn5	r3��^��<��{0�m�﹞/ʪ�|��BK3���~�8�?���y�7I���&�? 7��}�>��%$o3�^x�y�s���y}���ͤ�ȥII_��L�Ƣi�.nBq��g�x����s����U*�}{�����3��MI%��I�C�ә�/�|�3~���m��v��x�g��N6���w�s�K��#ǣ_���a�5$�}��獷�*��%y�|O[m�}���o��9'��~�w�ӽ����m�cf�]�$��l�R�[X l ��   �@�&�J��Nʮ�wWU��	Ȉ:Cg�ay��Il�ʹ����8��ڰW�.R��7�:ϭ6�^#�w4v��M�7�3��` �C��u\I���\�6�o`�h�vx$9g<���8渟O8��;Z�Ȗ#e����L�n�m�M�X,�������w|��GǾ\/�X�U�w,����˟�r���:�i�0u�-��dx�0�\��ws͡8��:������lߧ��m�}��y�m���i/.�{y���l��mŗDѐ�պ�sS[���}Ü�UO�����m�{�����=��sR��m�����&C ���%���ԒU�^O<z�%wgri8�o���y�m�W^![�Ȱ�!�ԗٙ��-O<I#��q�߾�x�񷪒��7�q��{�6�r1Kbq@�\�x�g��N6��U|��,Ͼ��[o6}�q��_{y<���yh�=��U^Z���mu#�ɕ�Zp��,ݖI7W/gS5ny����w�9�'ã�lٵ!<I%���g�$��.�RIW���?fg��֒:ω�$��ؾ��M�a#�3G9m�{��f�D�@"@҉�*��T�9�w��~�9m���������p�?�O� �"U.s�~�2Z��m�DK�3���^���6��f��$�_P�T�3~�y�m�ϸ�6��{�U㎬r�(�\�x����~O��w���[�������[o���q��J���ܽ�x�f^#n+qX���n�8�o��<^x��U/��,�>��������y�m��a8�o����W��!d�j^�6�ЯS�d�R���҈V	��[-�l�L���ݛ������99���sy��m��r�y�m��a6�^]����/<m���k�
�Ĉ��$�<m��ݽ�y�Uݳ�4�m����y�m�ٜf�����}�ߦ)���7'�$��������p�/��@��`C��Ah}E�A�R�Q��a�&�|z����vn�o��s��o�Ŋ�-��!n;�!8���$�~I��s~��/<m��~�8�o/ܼ�x����WߊK�~��8�ov}���n�D��������8�6��K�}�����m���&������x�G��toi���pە���+�M۟&��H�nmK��ۣ���눚��BUW83�������rFz�o�ϯ�獶{ل�m�{��m$�H����U$}�V߻�۳v�};��~�ՎXE˓�l��	��$����"��UU�q����/<m��~�8�o/ܼ�y��~�E� ����?g�f��5fB8�v�����x�����3��J�ʕ"�	*TREI>����x�fl����L��j�55MfhܝD�$@bU}�oπ|���p=�Á�J�R��)UU7~�ӀX�
��pP�#�?r�p����.�����O���6���׃��U^Z�n�tv�m<��b1[��cujM�9��W���{��ߧ{���~��FG�S Hܞ����h��{}��$���������i�����[���p��|�W���^��^}N罘s�~��~�ݿ��Rh�7p�����<~��������W�&o���3����=�̵ȭ�ۈ��$|��O��{8�ɧ �;0�~��*��o�~|�֧���۫��;�' ���8�%_w����;��>��o' U������(�һ_n�uM�Ą��pm p�`�� � �h��j9-HY٦��sl�5�u���V"�85�w8��vxE;7R�۱ܝƴ��]�t�'/hv�:��H���08˪܆X�m�t������
1�uv��+��ŷQ�;e���gc���%rt��&�%�N��zR�3ʶ�O|����pW�q ��*��Ù��{���{��绻ߟ?8��t0\��vQ7k�u�sb)��U��%�7@+ū�]���՗�����ݻݽ�䊵~x�.[�2�n;w@�׿� ���>��o'�T�T*���J��w6|p�-j��D�Q���<����R���]��o��;�>8�ه>��|�ë�]������ ǻN罘p�*I|���ώܽ��;�eD�bpc��rp>J�|���ޮ߯~|�o��$���n�Ӏc�|�2���q����<��8Ԫ�Y�ߟ�cݿ� ��w4
��m�m��i,O�mB{I��K�܏X���u�e�PoK�a�gb�����_��m'�XF�!�������vh{���R��{a߯~|3F}k��M�a	�ֵw$���}���Ո�h ������9�}��7v|p}��檪��I]������m��wdQܹ8s︸�ه��QJ���2���1��Ӏx�}F\�e�8�w..�_*�����|p�ߟ ������*_RJ�����z�ߖ�
�"W(˸���q�UUIv�/g�{��.�_q�3��k� ����3�^ͮS4�2����ڣ�&6����Ma��]f�Lɮ�?� ��!���B.
�~��v���s8��}Ǫ�/�E$��̽�����"����	.��{����_UR_�QT��~��>�~|���Nm$��T*����i����n㻻��w�ߟ ���>RI4��T��"�W���ܓ߿~ٹ'��l��vݩ4Ke��I|�
��9�>�v���s8�J�����������K6�D�#����p�_*���z��^����q�}�s#�nܗr��XE�qY��&�����%\�7<��DmɆ�ѡ������q9��N�C5��ﾟ��Zs�h��f��s�+�⌱G�Ày��|��Wʪ�ݿ�|��8��mRl=Ս^��"W(˸�e���o'�I���8�y��]x�w�pP���6�$�y���wvi�<��>$�\��
I�e�6�� �{�;w$����F���ۊ�rps&R�Kݙ��-|�Ws�@��v1�2@j&��8}�<\����YB׷31�{����p��m��?�@�ٳ3�Jj�L���jy$�׿>��c����}UJ��UE
��T���g�O��{e�n�ݒjk,�j�I���}A�!�H,ZH�J�TR���1��Ӏg�O��_r�����#bH(b�J��7~��En��D�#����4m��<���;��@�Y�%q�k�Y�h˚�kr~S�B)AU$RI
�^}���l����>�
�"@�1b>�{���'�s��帣����p�gf��RT�P�U����}� �2a���̈́�9��ǔH�۲I"H7�a�5o}o\ T�4lN+
�`˜e��A�kz.��������@uc$�R-ͻ�{K����Js^s�,rW3bȒ)�H0I�B��I�S�Gqd]��C`�aIt��\�I��Ԣ���P�J`h� ���*C@eə� @���p��� �}������� 2�eo��b�N)�) ���j'u�W'=��I            ��� �EclT�GYb	yo8�vPy��=�&n�7[A�\_�|;i,��D�J���q�]�t��#ol�            	        �P   �$m�       �l        6ۛl      �m     :n�u�{;E�9U��5�74�m���Z>|��f��t�l���Zr�	/Q4r푫���ʛv7b�]�kӢ����m<Q.��Q�<8�d�u�d�ٶM"�t�hۋ�\�l�{l�qj��tv@��$����k7:nkv��j��T�3/,�C��6;v,��8xñ�g/m�@�:�7 ��0�ы�D�[����9��ǗƗɺx�թ��d;��t9V�n�պ)w�d��-h14���x��R�1YL�7��3ubx�Y�L�8�A�t�H�;U溶̨L4�OeuȠ�$mA@�ge6�h�j�^E�&�}��W� lp�\�����/��r��kϝ�Mn��+Y{Yl�[��Gi�4�:���IV�����C�T�P%g�7=7Ap	���,½mVӅ�Fgu��uF5����w5S�ږ9u�=�
v�v�=��eҎz8R�ۨڤ��ݞ�h˜��v��UG.�w�y�z�g��A인)�_6���!�����G�|�|�a�M�����<�V�ͪ�"R�\n)V�Ѡi��[<p:����v��u�£�F��틜��#�'d��O=n":�ph�z��}���vkuY�v�60�6Ѻ�����z���>|~dD�ny��uƩ����YZ�Yxl�H�eK5�H��<�����b�;�����4ni87]�	�C]@ -�Mm��Pj�^�V�(���JBJ��Z�Q��Z�`�j��3�&��]�h�՚ҩ�?t�> 	�"�: �T(D��G��t(���w��{����w�ߟ�$ m�h�˛g��a%ϩ����� �t �  h�ܔ1�hc��V�[C�q��-R�窤}��Wv�8�z8۝�&�����$���K��8չJl��*[b�ll�趶ɶ	�&����E�Ժ�'/ND��r5���S�7	�;4l8�_��m��f�< Y��n�B�[�Nڃn��]�G�ҘVH��r��I�R�㇫�d6l\�m�.g��us��=�%_�)$9�Ư�\�J��v��������ɇ�RK��M8��]�D@\.Hp_{y9�*��K�UR���p���p�&���h�K1dIL�#rh�)�yzSO�~����O����z��rb$kJD���jK�$
��o�w���=}���mR���i�;��/mݷj@��$8{���v�/g)xRe&Re'�ݜ��,K��o�iȖ%�b_�/��bpRʧe.�n�zw0�5����G��=:v%3:)Cg���c|{�〝���֦ӑ,K��>�;��"X�%�}�{��"X�%��~�fӑ,K����iȖ%�b|a�oL�ˬ�4e�f���Kı/��u��>oD�A
ҩp%!!3�H"W!B!��)�%S4� mC�L4,B:�4���o���B�H(	����9�,O�9��iȖ%�b{���M�"X�%��}�w[NE$��J�L�ճQ��qF+#������Kı=����ND�,K﻾ͧ"X�ؖ'��{��r%�bX�����r%�bX��>�v�M�5e�M�"X� 6'�w}�ND�,K���m9ı,K�{�m9İS�2'�����Kı/N��3?����R��L��]ٻ/��)8�%�}�{��"X�%����ͧ"X�%����fӑ,K����߳,��F�ȁ�U��4ny.����P�+���^;�3:��������w/����E�5�s5�f�ؖ%�b^�kiȖ%�bw�o�iȖ%�b}�wٰ�F�=���%���k6��bY�7����{��I�H������7��bw�o�iȨ~��dL�bw���m9ı,O�k��fӑ,Kľ�����I��I��ٖ^ۻnԁ%�MM�"X�%����fӑ,K����u�ND��`��#@T<L�آ@a" ED�*�D���U� +D�K����iȖ%�b~����ND�,JR�ћkȭ��a.�r��&Rg�H �	,UX]D��?���ND�,K����[ND�,K��ݻND�,��Vȝ���M�$S�>-�g�k�˙t��flI�<�ﴛ�H��HO߷��i�ı,O߿����Kı;���ͧ"X�%���/�O�QX�U�sO3y�4��:�$�M��\ls��+����rsԴ:Yͭ�"X�%����ݧ"X�%����6��bX�'~�{����&D�,K��ߵ��Kı/��i�����a�SVfj�9ı,O��y��D?���,O���ٛND�,K����m9ı,N�_v�9?S"X�;��3?�$�SS5��r%�bX���߳6��bX�%���c�
�ș��w��r%�bX�����r%�bX�w�)0�d)�n�j�f����K��?�"`j&������"X�%������iȖ%�b}�{ͧ"X��@$�	�1Ut+�Oʑ"~��y���Kı>Ͽ�&Im8�-�.�NR��L��[�5�9ı,?� ��� 	߿���ObX�%���_�ٛND�,K���[ND�,K������k3Y���Z��׻mp��P�3.ОB�YL�2L1�̈.dQum��=ߛ�oq���}�~��9ı,N���3iȖ%�b_{��b?�X)	�L�bX��k��ӑL��L���ϭy,i�,"%�)xQbX�'~�{��� ? �$r&D�/߿~�ӑ,K���]�v��bX�'�k��ND�ș���3�e&�5r�\�fӑ,KĿ~��[ND�,K��ݻND�,K��ݧ"X�%�ߵ��m9ı,O�|wY�շ!��eɚ�kiȖ%������ݧ"X�%����nӑ,K����s6��bX ؗ����r%�bX��>�v�M�5ff�ӑ,K��>�siȖ%�b/~�{���Kı/��u��Kı;�}۴�Kı?}��w?���H��Ҹ��κۥ�v�Ύ���8m 5�     ��з+5�s��V���p��:N3
�%�Y�
��}n8�	'� �{�^ɺ�t��-����ū�8[�ܦH�����C�+�@�M��Le魱�	��r��؄۩[c�n7���W�1=���g����]O\^;Hq����[/f��i�Xx�&���@�$:珽���)��)�B�[��t���ճ��vzr��q��g/JTۗt���MɩsZ�ؖ%�b~�_�fm9ı,K�{�m9ı,N�_v��Kı>ϻ��r%�bX�w�)0�d)�u�Z���fm9ı,K�{�m9Kı;�}۴�Kı>ϻ��r%�bX��]�fӑ,K��=��E��R��L����kiȖ%�bw���iȖ%�b}�w���K���Dȟ��߳6��bX�%�����r%�bX���/mݻ�@ Ke��K)1$�O���6��bX�'~�{���Kı/��u��K�K��ݻND�,��Y�3my,i�,"$�_)xRe&%�ߵ��m9ı,K�{�m9ı,N�_v�9ı,O���6��b]�7�����߷ҘX�K��R��|����N��9��y��<Z�����rg���\�s&�5r�\�f�Ȗ%�b_�~���"X�%����ݧ"X�%��}���9ı,N���3iȖ%�bxa��̈́mإܷe˓��)2�)2���|���낣���2%���|ͧ"X�%��u��m9ı,K�{�m9�R(�L�b_ߎ�?C5���Z�����r%�bX��߿fӑ,K����s6��c��9"^���[ND�,K��w��r%�bX�����aP��_)xRe&|�������KȖ%�b^���[ND�,K��ݻND�,�>�����Kı<�zRZ�,MF吗nK�R��L��O7vm9ı,A;�}۴�Kı>�����Kı;���ͧ"X�%��}������)eU嬡�:6�-M7nc:�&gf��*�ٓ����y�#�^�X���35��"X�%����ͧ"X�%��w�ͧ"X�%�ߵ��l�K��I���R��L��^��/mݻ�I&��Y�jm9ı,O���m9�12&D�?w_�fm9ı,K�߿kiȖ%�bw�o�iȖ%�b}�e6��m���"K��K)2�)nM�ͧ"X�%�~�{��"X�G�@$"���^D�;��iȖ%�bw=�siȖ%�b|}��/rN�sN�k3iȖ%��>������bX�'�����Kı>ϻ��r%�bX��]�fӑ,K���ӹ��շ!��eɚ�kiȖ%�bw�o�iȖ%�`�}�w���Kı;���ͧ"X�%�}�{��"2�)2��J�>�{�[���XӒR��mYFˣk�!R�`R����]��VV�S_���7L�3Z�5�j˚�O"X�%����ٴ�Kı;���ͧ"X�%�}�{����DȖ%���w�m9ı,Kӷ��̚,�jj\�fӑ,K����s6���@��L�b_~���"X�%���w�m9ı,O���6���!�2%���ߊe�̖M[���̺�fӑ,KĿ~��[ND�,K��}�ND�,K���ͧ"X�%�ߵ��m9ı,Osޝ4�Յ5u�uu���ӑ,K,N���m9ı,O�ﻛND�,K�k���r%�`b�XA���;ڂ`��2&}����r%�bX�~�rg칖��IR��L��Yy�|��I��K�k���r%�bX�����r%�bX�����r%�bX�}�^��fQ!�=emt)����gɪSi��\6f���ڸ1��qk�w�.��;[T��w�Kı;���ͧ"X�%�}�{��"X�%����̀r%�bX�g��m9ı,O��|e�Bi�W.i��fm9ı,K�{�m9�ș�����6��bX�'s��fӑ,K����s6���X�DȖ'��>�n�ܷe˓��)2�)2��o>9K�,K��>�siȖ%�bw�w��ND�,K���[ND�,K�����D�H�c�r��&RbT�Yy�|ND�,K�k���r%�bX�����r%�`~H�D����6��bX�)�����0�;��K)2�(���s6��bX�%���bX�'{�xm9ı,O���6��bX�'�H +H�pm �߻�~�@ �5is��6����%��� 8�l �d�8 /�$�e�7g����5�c)n����v�@�ãod�[/hh��w>4�O��A�i�79��g��[��ˠ֞z���1�F�l����k�4#�W<v��F�T;GA�c��WC�v���Ո=�qќk�&�ˮm���۞]�Geۗ���M�D�<�t���{����~:�)e�9k,p:��/'U9����a�v����B�����L~����|�?�6�u\�ֳ8��bX�%����m9ı,N����r%�bX�g��m9ı,��7n�K)2�)w&j��r��r���35��"X�%����NC�E�@�MD�?g����r%�bX�ߵ�����Kı/��u��O�F!�j��2�~�Yl��"�K���)2�(�?g����r%�bX��]�fӑ,Kľ���ӑ,K��~��"X�Re,��חm6�D�K�/
L����?w�fm9ı,K��ߵ��Kı;߻�iȖ%��H��;����ND�,K�tt��!4᫗4��6��bX�%���bX�'{�xm9ı,O���6��bX�'rn��&Re&R�����nK��m���<��u�ub"�K��v����Jت��t�u��!��榭�u���3Y�m<�bX�'�����Kı>ϻ��r%�bX��]�f��'�2%�b_�~�9K)2�)?�Z��+��Z���rm9ı,O��{v��@x����~V(� 8����_Q?�`���'9�}��r%�bX���~�ӑ,K��~�fӑT? C"dK���C3�&�&�����r%�bX���߳6��bX�%���c�(ș�����r%�bR�����^�I��K��M[/�F��j�f����K�C� "	�3�߿kiȖ%�b~����ND�,K��ݧ"X�%�ߵ��m9ı,O~�j��r��nY��9K)2�)n��ͧ"X�%��F =��~�O"X�%�����3iȖ%�b_{��i��7���{��o�����P��w�����=c�]���[�B]�+u�91��,[$�)xRe&Re,ɺ�KȖ%�bw�w��ND�,K���[@� Așı?~��M�"X�)��~���Cq�	r��/
L��,N���3i�?� DȖ%�����r%�bX��w�ӑ,K���w�iȖ%�b|}��-�4᫗4��6��bX�%���bX�'{��6��c҄	"F{ߐ�&��HB&���5r
XHB(}u4t&�1�JK`Ē�KBX�ĥ�R@u�E�0!��Đ �y�*�����BH%+HBBE�EB#��P�%"�A�V�&�R� A5��	
$# A"D�*F�@�7=$)��ꐄ!�a��! ������e'���+�� E��*8�#�{F�#UsH��"��2�2���u+�HsQ� x<���8�� '�|��$UG���U��pЯ�b�4P *���Ȝ�����r%�bX�}����r%�bX�zw3���0Ժˢf�Z�r%�g�"~����ND�,K��]�"X�%�ߵ��m9İ���J���NR��L��O
�"V������r%�bX�}��v��bX�'~�{���Kı/��u��K�e-ٚ�K)2�)w���������vmt�ղG�[��&z�r�����Y��u���ۻ���/綸�ec�yı,O���ٛND�,K���[ND�,K��ݻ�'�bj%�J_}>��K)2�)g�ߓV����sZ���fm9ı,K�{�m9ı,N�_v�9ı,O��ݻND�,K�k���r�!�2%��u��h�5����M]ff���Kı?~�]�"X�%�����iȖ%�bw�w��ND�,K���[ND�,K���e�v�@�ˑ�&Re}E%e-�o�iȖ%�b~�~��r%�bX�����r%�`(�u��ZJ[-amW��Q2��1\Z�h�bK0��Z�5I!;&�/��(�y"k����/
L��L��tg�חn���v��bX�'~�{���Kı�����[O"X�%������9ıL��3_)xRe&Re.���.ݹ.��XA��X��Dz#�\�p:�A�=���l�f�Z&�͂C6lɶiѫ�4��6��bX�%��bX�'{��v��bX�'�k�ݧ"X�%�ߵ��m9ı,OL=;��M[�j]e�3Y�m9ı,N�_v�9Aș��u��iȖ%�b~�~��r%�bX�����r%�bX��>�v�M�5ff�ӑ,K���}۴�Kı;���ͧ"X ~H��2%�����r%�bX��k��ӑ,KĿ^���&�0�������Kı;���ͧ"X�%�|�{��"X�%����ͧ"X�"� �D�w���r%�bX������ܲGwr]�&Re&R}����Kı;߷ٴ�Kı>�]��r%�bX��]�fӑ,K���"��Y��;��ֵ�kZ�feS�7kf���{Z2�nA�@�� �6�6 )D�8 ^���2WE<�Pܮ�rkGp�D��w����`���K:w`�yq���ƧGL�li�"v��1ۧ" v����9����#��Y�ҕ�����3��=9^�[q�:.�7aQ�3��db9Ys�ɎZ����_�{�V���6v��nW�jiGe��X�J���q��,�B�-��p��x/V,֐�����^^.��Za���{������ߟ��fw蕯��ؖ%�bw�iȖ%�b}����r%�bX��]�f��D'�2%�b_~���^�I��K�M��ϝ�`�ֵ��ND�,K��nӐ���"X��_�fm9ı,K��ߵ��Kı>�_v�9?Er&D�;�����n��䏔�)2�)2�v}��(�Kı/��u��Kı>�_v�9ı,O��ݻND�,K�tt��iѫ�4��Y�ND�,�Tș��ߵ��Kı>�]�v��bX�'�k�ݧ"X�%������ND�,K��V��#wj[��rr��&Re&R���iȖ%�`���{�6�D�,K�뿳6��bX�%��bY�7����>�\+$@s9g�ѹ(2*Q�f���m\qm��E�u=.��<\<�\�t3T�3Z�ND�,K����ӑ,K���}�ͧ"X�%�|�{���%�bX����v��bX�%���gIauu.f�iȖ%�by���fӐ�+�B
ł�	���H- �� �P:�D�+Uh2�@" �v�4iCm��,K�;�m9ı,O��{v��bX�'���ͧ"�ʙ���ߊarp���Mj�]]m9ı,K��ߵ��Kı=�_v�9ı,O�ﻛND�,KϾ��ӑI��Kܙ��e�Q�dq����(�,�
	G"}�i7�O��fĐI����n	"~�{߻��"X���^��L�jX"�%��^�E�bw;�siȖ%�a�I��~���=�bX�%������"X�%����i�����oq����������YH�+{���̡�U�c����|���z�!PT$S�j�n��I/�^��I��Ks~�8��bX�%�~�bX�'���ݧ"X�%����ͧ"X�%�Ӻ:d�4��˚55��ӑ,KĽ���ӑ,K���}۴�Kı;�����Kı>���6��X�%�釧r�F˵-�G$�/
L��L������Kı;�����K� >Q
h�MD׺��ͧ"X�%�{�{���&Re&R}�خKr�\j"�|�Ȗ%�X�����r%�bX�{����r%�bX�����r%�bX����v��bX�%����$4Y���ff�iȖ%�b}��iȖ%�b�����r%�bX����v��bX�'s�w6��bX�&�|�{�e�5��ˑ6tCnY�9��^�t{WD���N��a��5.��<:�A�P+O�����,K����r%�bX����6��bX�'s�w6*�%�bX�{����r%)2�){�5\L��h�28���^�K��߷ٴ�Kı;�����Kı>�_wY��Kı/{�u��A_䂄2�D�=���d�~�k$&�����r%�bX���fӑ,K���}�fӑ,KĽ���ӑ,K��߷ٴ�Kı;��;p���udԚֵ��r%�` �BdN����m9ı,K��kiȖ%�b{����r%�`l � �TM
ȯ����K)2�)|���`J�8�-K�k6��bX�%�~�bX� �G���i�Kı?~�]�"X�%�����ͧ"X�%���>˙��˙�D��垊<<�ny�ς��8��CM��=��j�y�ݸ�j�bK�U�����K��߷ٴ�Kı;�}۴�JRe&R���|T�=)YI��I���9K)2�)<�־��*Ƣ$�)yı,N�_v�9ı,O����m9ı,K���m9ı,O}�}�OK�t���O���
��
&Z�����r%�bX��_�k6��bX�%�~�bX�'���ͧ"X�%����ݧ"X�%��zS�����5�Z�3Z�m9ĳ�BD�߻�[ND�,K��fӑ,K��u�nӑ,K�]�͗�^�I��Kܙ��d��Q��WV浴�Kı=���m9ı,�_v�9ı,O}���m9ıL��sg)xRe&Re.�f��I$�v�,�.��<�t��8,��Z��   h�mi���:W�Vk��B��sێ,[o[[��	��u�w!��X�j��ș$�v�g�r�ۋm��X���u�=��d �+ˬ�{>���������k�ֻ+>�]Sm�<n��ѵ��{j�h�9k���H/M;:�b�g������T��V�Ɲ:���u����Rʧe,�����{-��n�5'k�k'8��Gfy�1F�ȃ˱��۵��V��7���x�?~�]�"X�%����ͧ"X�%�{߻��"X�%���o�iȖ%��KwFk����� K�>R��LK�u�u�ND�,K��w[ND�,K߾�fӑ,K��u�nӐK��KE���*(㸠�K�/
L�bX�����r%�bX����6��bX�'{��v��bX�'����6��b�I���um��5w.Ȉ䜥�I�b؞���6��bX�'{��v��bX�'����6��bX��L���w��/
L��L���Z�+��PjF�ND�,K��ݻND�,K��}�fӑ,KĽ���ӑ,K��߹�)xRe&Re.�8�٬��%��2V⇷mQ�'&ճĎ.��jq�N�\��5uQK���k�z�=ߛ�oq��O����m9ı,K���m9ı,O}�}�ND�,K��ݻND�,K�~)֙�I�u�Z�3Z�m9ı,K���m9��t���nD�K����ND�,K��ݻND�,K�u�u�ND��eL�b{�w�,ֲ�պɫ�sZ�r%�bX�}���ND�,K��ݻND����;���Y��Kı/�����"X�%��u�v�jX"�9R��L��[�;v��bX�'����6��bX�%�~�bX�'���ͧ"X�%���f�g�PH��#�/
L��L���wY��Kı/{�u��Kı=���m9ı,N�_v�9ı,O����~�/Jab�/3���}�����s{L��ӱh^SXG��Z��N���^�!���ͧ"X�%�{߻��"X�%��o�iȖ%�bw���iȖ%�by��)2�)2�U��������ֵ��Kı=���m9ı,N�_v�9ı,O3�siȖ%�b��l�/
L��L��Lkb�	�kV�SiȖ%�bw;�siȖ%�by�}ۛND��p �j'e�ȗ����r%�bX����m9ı,Kӽ�C3��-�Yrff�iȖ%�by�}ۛND�,K��w[ND�,K�~�fӑ,K��w�ͧ"X�%���L�&��ɭ\��\�r%�bX���u��Kı=���m9ı,N�{��r%�bX�g��ͧ"X�{���?�?^߼[,����5�S�;34�5�)щZ8ͧu/K���G<ѩ���Қ�̺��5��"X�%���o�iȖ%�bw;�siȖ%�by�w�6��bX�%�~�bX�'��L�,�,Y�)xRe&Re-�;R�Kı<ϻۛND�,K��w[ND�,K�~�fӐı;��;q�YDq2�K�/
L��L����QȖ%�b^���iȖ%�by���r%�bX�����r%�bX���5�*F�D��)xRe&|������m9ı,O~�]�"X�%����ͧ"X��	�$��Țֻ˛ND�,K�N�wZ���k2h��ֶ��bX�'���ݧ"X�%��~���ͧ�,K��?w�ͧ"X���Ow6r��&Re&R͉��mے�5�qPR��Dq�;^BuKL���a#�z�Y[�y�tu:��#��>{�7�ı,N�~�m9ı,K߻{��"X�%�{߻��"X�%����nӑ,KĽ;܄3:I��5�&fk6��bX�%�ݽ�Ӑ�T��,K��kiȖ%�b}�~�v��bX�&���)xRe&Re.�55i��dl�Ie���ӑ,KĽ���ӑ,K���w�iȖbX�����r%�bR��׳��)2�)2��3U�r6��̚��5��"X�%����nӑ,K��w��ӑ,KĽ����r%�bX�����r%�bX����N�5�Rk55��ND�,K�߻�ND�,KʨG?w�����,KĿ�w����bX�'�k��ND�,K��G���@�� H�"6 @�E�h�U���� �+T*F#�@�B0�*���m�I
��rY BQ���
�JB%�������@              @�$�KsN���M�9���be�%=t7W3�4����G��`�Q��W"0���%�Y�����    �      �       �`   �d�l       &�   6�    l�`      �h    ��[�6��E�$VŪUۯppt�I�6K�s\�ɠp�R��45R���	{z��E�s%���^D��%V�$���ْ,��b����q��U6P�q����$6�@��ĳV��tm�Wn�0�;m�,Bk���ٶ�Y�i�&x:���PV��e:��&�pv�.�r�b6�mԠ�!��ް#���v1K������:�Þ�\�d:����xG��J]���z�c��x:\¶�S�XW4���j�|����햠71���&7+�{P���M�ꍗjցW�kj�����ڮӲps�;)�����Xv����	���۳.�:�L�K�yűڳf�h�hీ� ^��\�籙}l�r��Ѱ� 7W ��b��1WO:�8�ئ�h��.iuH�nG#�;�h�\��b��·]sTf��U�n� ɻz2�<��ٌkOp�Y�;j��k�9���Z6^SsHz�rF3��V1�.�hU�'����B��\�]�,����n�N)ŉ�+�*���	��h݋�l�QtU*������]n<@����f��\�/��9��٬ݱ�ș��v�F�g�-θ�"��	�k:�vZѣ���Q��A�n#8
�43��n�e^^/N�Cd"-F���5v
����I�H$	�e��la��Z�h�F�5u0^�Z7#RE���J�эѧi�%�R�ۖ�� �7U�M4!*�8��qu��t+��,6�-�6�v�$�ЛWV�ˬEq�(�
h� >�@J�(�����>��M � |(n��jMkZֵ*�F�����<�ķ����m���   h�6ؒ^�;K��ZnbMn�u�����&�Y�;@��ZgZ��ݎ�&�
w�;�2��Rn�al-�Ō<m�Wt0�@^�6N�����qulx�ccң]�^��vG(u�\�96w���e�g]s��b6]��*-ɚqXnG6��l��e��|�|o�?2�($9�Җ��st�f�9��6��\�P�vCM��Ku�8Țw���ڪ}���7��,K�^�iȖ%�b^���iȖ%�b{��۱�Kı;�����K�L��[�v���W��$�NR��V%�{߻��"X�%����nӑ,K��w��ӑ,KĽ����r'�J�L���/���i��vDG$�/
,K������9ı,N�~�m9ı,K߻{��"X�%�{߻��%&Re&R~�ƶY!,Pj��KȖ%��D�����ND�,K����[ND�,K��w[ND�,Kܛ���)2�)2�չz�$A��nk6��bX�%�ݽ�ӑ,KĽ���ӑ,K���w�iȖ%�bw;�siȖ%�b}��eΙ�[������89��f^KUg\	r����m��ˑ�z\��L��ݴu"�{�7���Ľ���ӑ,K���w�iȖ%�bw;�siȖ%�b^���m9Ǎ�7������Ƥ㠝5�����K���w�i�sH�E�"�+� �=�AF&I�V�z���\��,N�y�ND�,K����iȖ%�b^���iȖ%�bw�S���i��K���)2�)2��~�m9ı,K߻{��"X�%�{߻��"X�%����nӑ,K�[�3n���	(��I|��I��I�^���m9ı,K���m9ı,O~�{v��bX�'s�w6��bX�R�-�۶�m\n[����^�I��I���R��ܽ��7o5�;�'}�x���L'v�]%���;c��݄�ur��WbX[�,�n��j�tL�I�w;V���Z�U�x��_��{r��2B3 (�`�Z+���I$�fk�����;ܘp�;x��`Dby"Ĝz�U�׬��ςH���� *�C�i_��@:���ۋ,{���!���jI����36i��rp>��_��@���9���Y��	ɠwYM ��huVh^�@�����-�?�.�8#8P���>N�:�鹮�����-ɶ-��X�<�����p�t<]�k��C���huVh^����-�|h�3n��d�N2I$�{�'>�T����36i��rs�l�nڍ�q(�$�M �_���e4�ċ��h�/���,�+vAb�dL�I��O3y� 3����<�U%U�R�U���G:� ���X�̀�Ʉ��	˚#Nh1�G@�{������yW
�1��f������pe���9ՃON�HܨbM����7f���eH���}������4z�h{l�<��<x���,S$BQI�޳���gsf�>ISf��N nk��<�����"X�%�@����w�� �U���4}wĲ��`a2()�RM�wg 75���ܜ���@�DV��~doD�I���@=����& ﹓�J����U�;�ڪ�U�4�N�����]�` 6��om�l� ցu5MR&�1���/ih��юv��v��[����r�,�V�.�ݜh�lA�I�u��.`ݝ�q�m�6��-���ݴ6�*˱Gm��k^^���{�vq�h^��o ���<wn�N�̚�Y:�u5´�C�뗬�/b���`��.j�Y��5��3Y���!�S��7����K*��+t�'7�n�NMdc��6�z�v�EG�a���w\�p�%��O 3wg ��� ;�d���`gq����۽�i��j ���y�s��%���ﾚz���{z� �X�"k (�$�� �m���N��#�p=빠�.��������U&��^N w3g ����I*o;�8�~Ǐ=���2D%���4��^�7��wvp��������t��(qϣ/�p\뵰R%�n��p���s�e���T�"x)1��D�D�"�rh{�s@'.h�Nh1���U���_�=!4j�]jnI=�ﵿ�����.�:UI-�I;�~� f��罘p�"�-g�D�#�h{�� ���6�&��M8�ݜ�U���1��Wu�fVf�s��9��4w+4Ş�n�,R,��I4�z���U{��= ����s�8�J��O��ߪaY"��<7F3Z�Vm�ɛgZn���:�&��ɬtݯ�$�Ѷ���~���@:���f�v^w�aHy"B�h{���?�]���N�|���N��j��m�i���N w;��{��|R�ﴆ�[ �BT� 0BR��҅`��1����BF1*>
|,�P��� SI��(�Ȯ�d�$#FHIr��Kڤ�3��8�q��s�~R%�"Q�A94?�Y��@/����@:������YS�02#+�� �s@Ӛ��ַm��x�������YK�������X��Kk�Rߞ���[�%ER=N1����$�O 75��s�8����U^0/��u`�c>Ė8�jE&�u�NjT�gr�_ 3sg 3��pS^�ݐX�Y&�h�h^�@/Uf�u�4��Yc$#2� 9 ;����<� �w'ڤRIR*�J�*Uo�1��;x�$Dm�ԍ
I���@�3�_��u|��[�����Slt*�::�u��&v�����h��\�+p5:���\�� Ab�	�E&�u�4yڴ�Y�$�^075���櫔�m5�Grp{y��M�n��潜 �fN��x�V�02"(G�u�h�����v��[��"b�����4�Es@�kZ��`�6��KJE&�u�h~���}�����@/Uf��u�I$�Z�E#��v�'gǁ H ��i6 /H  6���T�3(�y}���Y�tn0�%�ɍ+v�G�����y���X�1c��v:�#�ގ�F�gYא�i<S�������nG)�78�s�:�v�g�����;#��˄e�N���7N5m�r���N��[�k�=����www�|zE�����3�z(��{s��|�;���8L���M����F�����0$��<�j��� �U��٠vr�!1�++��Z�1�41���he�p�&X��
I���@#�:ZրF9�}����ܺ����@:���j��f�^�hs�~Y!�D�"�rh��@:��z٠z���b���x"�U8+)խ�}��煝�Ѻ��J�i���ָ�َl�Q�2 ��t<]�F�L~m���� b�F9�2ִ���c*;d�I��d�*��"����L^*�,�����$���rI��f��0K�Yq%�$$�h^�@e�hc� ���^�7na^��(���M�/�������� ��h��Yc$'���E�y� b�F9�2ִ�=w���0HY+���^�Q�[<I�r3�ɓ3��ss���aUsnl�â^���Q��b�F9�2ִ1��>�]DHS$BRM ��h��@:��z٠yϮ9�$0ȔdPNM;y�����ڮ$�!%k�:}���[�jL��bh���hB Em�Pq�� @r ��Ze�1J�Pv��#�+%�
���k@� ���l2�b�f�� ��!e��V1Nh��6	 �(x��7a�K��/�/��JR0 p�0	r4�ԉ^
A��aq���bZј�Yi"�_H���1�ȧ���R�� �"�����]�O�D���C��*��x���Qj�H9�M �h.�q,���DE�� �s@���hq4	h�ص��D�I�m�׬�:�M ��h��17��&�R�u���>7����ɹ킶���:�^<�a3pg�$	6�LIc		$� _��@�e4�Y�m���ܭ��O�5I' ��0�ʪ�a��8�ݜ �u��VX�	�D�Y2) ��hE� �s@��h�-����P_�*��� 蹠�hMς"hT�J�'���nI�|S,޲��MǠz�����f�WZ�W���—���o�r6k4^�0-�k)ъ��b]��y����X)��	 �Ƞ���)�z����^�@�{��,���DE����4�ހF9�1��#��Z�~��"I$�*�^�u�4�S@;�f�Ղ\�ˉ,cS���mU7�͜sf� ﹓�c�e����n�,rb#sI4�S@���W�g�k����ܜ�EBHBT�:�߿�ڪ�UP����n�[�k -���  $  �Ut�kȁyUp"�-�yla�� z�-�.�vS��n:]\5�#��W&٤�=u�Q�۝�nyn�!.��y;z��Zv�:�����r��q�\���6�7[�\ksu�l�n�k�W���g*��z��5�m����z�u������f�0�4�]��X�5��{����o{���{�����Ą�ƶC�����Xk�&��N�b��U��,s��v��R�d��uk�IE�"���l�*�^�{zϳ?~��͚p���l-H�.N �[�c�M ���N_W���"$)��n= ����)��@��z���� ����	ɠ1��	˚Qo@9�hWz��ʟ��2,$��w��������/YM�|�ѷ�����%���Z����m�����k��]sPܼm��(��8�&�Q��&8��@=�� ���{��Ix�����`�]�����	��ֵ�$��~���SkG�t�P7c�O� ���h�l�;{�� �Ɉ˼�ffhM ���4�f�y�U�2B~�%L�C@;�f�t\�c�G@'��|{/��eQ���4�����	�����u������,nA��7�<;2�Zh��[���!�s����=.f��1�&�	�
d�JI�޳@����w�Ͽx����@����"2('&��ra�I$����� w7g =���I����kn�հ�(�$8�ݜ �.h~�������4�M>Jn�����.I�ڪT�svp��8�e4��hX%ͬ����L!$���4�&�N\���Ϫ���$��.��t�V"���W=��g=��*hu�P�gn���9̈́��������tq4r�t\�c��VX�"2dȤ4��h�l�=W��=�)����28�J�/3@:.hLo@��h�������"m��cw'RI$�{�|��N w���ʫ�Kj���EK��UZ�K�T���g �/��&
4�d~ʼ�����4����������brFp���G��];6.z�[\�\iQ[�G��a���a�Fܛz��Xh�� 蹠u1��������/������&8��@=�f�꽗�=�L8�s'2��:�X�t��z�|��HjJ��l﹓��٠v,�+vAc���#�=�)��4��������3��2����4r�t\�9�ց��ܓ�#M� Z	R a	XF,B	�$8�d0�( �)��{�jMkZֵ�Z����7gl�X �� �� ����H�ol��N�o;���nU���<>��6�\�[�=h�������qN��<Fszc/q�h'T@h�h4�ѶcWv�s�	96�I���z콊#pVCa����v����n�Sv�[�ۖ^_-ٜ�ٛ�f��<�έcC+�=<�9^��ROc#;���y�q|r�VH��g�Gkf�p�q�냖6��8Ї�p;OE�����<s�LC�#��<�@��ZG@'.h|�轲�
�eW��u1�����4�d�T�=�櫉���2Y�����8�s'���ݜ�so�y�ck�V���$�j������ w7f��^��YM�[��#�h}��u��w���z�h{m�m������Q)eS����5����Iɤ�k���m�6�a�M1��u�*u�z�<fff��ƴ�&�N\����g�[�$7F��Z�e6	D �SJ6O|��nI9��krO>����T�&ër�Y$ddj(�8 ������7�:8�<�[�#���D���z٠{_U�{�S@;�f�qn\�q�`$BNM��hM ���4�ێ^�t��D8����.����s={v�m�p�xa㑽6�wJvu�<�cE���M ���4n5�}<5YS�b�C@;�f��u��wo5�{�mR�����c�Pv\d�$�svpr���^IH�Ud)4����j{��ɹ$�Ͼ��:�K�YpK�&�h��h�)��@;��b�r�dHn�Y�+2�\M ���.h�kC~?�^���%^g,����l�6����,6+�n���nmd�;v�4r,��{+0�	˚"��ƴ\M ��� &"d�4���l߿~M���|��N w���:�"+q2b	� NM����e4��hu�@����~�Š{l� ;�d�{�8UT�r�Uk�;��{��k�V���$� ;�d�T�����ߖ����ciH�j�����'��=zn�uq<j�>��������d��#bb2	�"G$�߾���Z��h{l�:�K�%�)�g����9�ցˉ��4E��g�[��91��)��9s@$\�9�րw��噙G����{+0�	˚"��ƴ\M ��� &"d�4���l�=��>�dÀ�2pHUD�T���U��i��M��� � @��2\0&`�
���B�
��ԛ. �@Z�F$!թ!�bF�!K(J�ᴔ!Ysfʋ͂ �bA�9��
�U"Mp���$�FBd�)�6�"a�����e&"Pn���JQ����l4xm�X`@�$��*���%ȱ�ԅ��t�O530lD���N�A"M�/Ȟ�cE� �"E�BP%�B	$R"Bp�\�#I!�	 I�����bK���Uz{����߮�����               [j�{-K�C��y֝@T��ܬ9+���Y$�kz�	�#�f6�nDJՒY�m�:qtݒ`                   mp   ��6        �m�  6�     6�      ��@    ����2m^$�U@�g�1����$l�n��c�v8���]�����Ͱ���t��W�L ۭ���dWm�k�Kƌ��,���wd� ������ S�PHF�9�G*��}%Q*qpph�d�l���#�a�[N�ȶ{HG�By'%]�	�dX�{m�d���0axI!��0�f���v�H��"��ϮQ��u���:�6/a��x�rn˙w8�s�AO$i䛎&��m��IyWr�)e�(ָ��F����q�s�:���j���>y�u�ۅ��tu��$����C��Q��mppOvJ�G���ی˺M�T���=+8�C[����%�n5�9�mr��͸��IP��9jY�q�r��hfx�Z��Jx{AG�Vy�OD&��R�YJC��`]�u�ۨñT����-휡E���[�/P���]���ٶ��)�q��e���n|i:Bc��p`�ԻY�-����.�s��'[n6][]���3�9xmeD_J��2�K��a^�Ƴ�ظ��g�l��yU 
��B�n-�=���	/k��4h쓉��sm3�;hȂ*�ch�)׶�um�i`4��V�mv��lM�ya�x�Z7H�m�kn�K/=���m�٢{v]�oci�3�uv��Ԅ�֑f�'Rqh۬h�����2�g%+Z�\�-�m�pI�iB�M���L[@�r�[3UF��r;S@ ���ݳ��$�EH6�"[��o[I�%隔�j�.��|��==X��.*>,@} O�P����{�����@����&u��.��n��8 ��8�J$���]\�Zv��-�Mغ5�28ѭdF�={#��;Y@�.WA���>�iӓ�D���z�Z]�4��ny8�.��s����v�*a�3uN5�M��u�/&���h��ƌm�8���|�ԅ�4c<�ix:#>W�s��k��眧R2mft�zN7[�~w{�{������7�D�
�Ύ�.�U���C]��O;:�Ci��(�n6��Gj�& �"��-}V����4�٠y��b?D�����=�S@'.hE���hOW��=x,�2,$��w�� �����Z�e4�B�-b!��"G$�z��sq�����4ߪ�.��%�9��I$�=���=�)�z� ���������Zo�&�F����kr�{s��|�[:���T61Ob�����ݱdnB$�FF��^���z� ���iRIx�6�_ :�+e�FT��h�֦�߽�[�H:����}�����|�ց���	�81$Q���z٠u}V��YM �m�+r�1����d���=����� w���ԩUS������q�@�葊dXG����4]k�=����xX�JF�m�JYN+qs��<�tDI����y1��m�\�6�fL�idN�Y�dXI �m�.����h�)�u�ikLq������sq��@'.h^��~$��ԑ���h�)�j�R��������ݾ�׫.����]ʎG��I$���8�ݜ�Z�k��s�X�	� E�%h���-��k@�kZs�~ݝp�$��*�ۋѪ;=�,�rG!9
��ٌ���Au\ە�BIV�^f���n5�t�� �������ȘE��r�����RI_�- ���@�u�@����~���%��=��> w���j�o�7o�wo5�1��|���Iq�5$����כ��=��>��J�*��$��j�'�>��ǖ�,d��$�' ��2��J��3_�w/u���_6�������&HrK��V����Ż>{�vuNV�]����X9�k�6plu�x�Ƥ��;�~Z��Z��4WZ�Ş�n�$�K#s�R-�v����^��r�|�k����&302��/2�r���n5�tv� ��� &(�i94WZ��}��=��>�o;�8^��Enb& �	Ǡ{_U�{�ՠ�@�u�@1���g�Զ��I$��$�Eҙn����b�|UW@�@	� )D� ���X{TZ`2�uX��ôfE�8�c���5���!�6��;{c����'����]�Q�vM�{��w�?>|�Մ�b�pm��s�;�Gk/�yݭv��Hm�p�h�����ƺ��<L �z�6�w�S[�stv��u;s�K���w/k����çY����wt|�����K*�-f�&tv�i�%cg�����Z�fB����DH�9��1L���;���@;�d���_Լaݼ��=�kk]�V�?)�d�- �m���z��Z���ͥT�l�яl|��'e�IrN)�����h-k@'.h�U���R`LjH�k�yڴ�̜�T�����MumީwR�~�̭��h���-��k@��x��l���qPR�j+���]��]KOΫ��;��l�p�gf�,���^��Z9s@�z7�:Z� ���p	�"ENM�ֽx�ϡ��b�D0��Z�hd Hɲ���A�������:��$LT� "T B)A
�ON���Ͼ|��u���NjI��ujV�dL"����;�o1��I&������=�_\s9�$b�D��=�Z�	˚T[�:�ށ���W��,F)�d�- �m���z��Z��Z���6�6�Q1��?ѵE۵�A:d�d�tu:�9�nN6�p#s�81��#�h�����h�h{l�=�����N1�#�9�ց�ִr���	��y�� ��dn~�E�{�ՠ�G��?@@и� H!E(('�\��@��V�{��c$�fHd���T����כ��=��>�o1���1�	�$�Q���=]k�=���=�j��٠Uثʈ�JF�b�-e�����3�[���vq��ˑ�z\�m2M<�@jb& ��#�@���@��c�}̚��R�^n� ����&
�Q�\|��c�-T�/RB���8_w�@��(��rzcň�25%����8����R�o�y��w/�P�KX�!�#�h����� �����J���t��s' �<VV�bp	�I��}V��;V�w���ֽ�qK#I)J5�K�����!դ�����sۘ��.�88ϣ�TsŞ!�&F�H&Ƞ��ԋ@���@;�f���^��}V�{��c$ȏ�Y�/2�	\��uE���h-k@;*�'�ґF��@�u�@���@���@;�f��.1����e�2��n5�t�� ���uE��_\sHd�2,#�@���@;�f���^��}V����s��MݒHժ�3v�=<���
.@p��k�  � �*���zv��gyۙ��sG8�1������rlhB3�v�<=Ouѹ�6��ƹ;Z�vn����[��9����6�cK�rvE�wb�Ӟ��9�M&���`�5;���.{t��<�^��ݪݔT�p�q�]gRm%�[�Ԗ�$��lCd�ow��i��ђ�Bs��'V2h�.m��-i\�Fꇞ�7�����4�#ȲG�[��=]k�=���=�j�:�
����sՙY��uE���h-k@'.o�U$�6wm2Ͷ�w �ܒ�v�k@�kZ9s@�z�{�ۆaM�A9����;V���^���^��}V�{��c$ȏ�Y0r-��ށ��n5�t����W�.��,c��e���ap�a냮cr��t �v����N�೛�פ(�3�m�"ށ�ƴ���J��|��z�4Y4d&�Y�'�g�]�#��C�Ɣm$P+A�
�:����������ۼ��^f_ ��2��R��r�U��AAӊ4K��w/���	Lo@�zn5�|���1��ddY#�@�z��ֽ��yڴ�B�-b"XӘ��=����UU�3_�w/u���_ ڪK�������JYT�ac����swRs�#c����v���[,�i�K��ˤ;���ԑ��ߖ��;V���z��z��ܮ�A6E��Z��Z+�����_U�~���e��d�Rj"�|�� ��2�5���ܹ�HS����3W	�*f���T��9��BЄv�@��	"0"��dd�!��!"�� B0 ��aᡵ���#|`�!��*��(A#= H�AE=S�.׀> 	�C�;4 �ް�U�Q_�y�J�PO �@��)!$�]R��﯀g��| �7���	�4�PmǠz�נugW�{�ՠr�^�{n\1�S1�azVF����JczT[�%Fܲ�Ѥ�r!�W�����k�\Y����k�<�Y�e㑽���wJvu������3}$��Z�%1��-��7�|��zcň�ȲG���z��zVuz��ZZ!V����4�'#�@�zl��-k@���o��[Y�L	�I�՝^��;V���߳r|
E�h� P�(�H����y��rN��3�4\���$z��Z��~~˯�@�ί@�{fXЛq��m�n<N����e	�a3]��\g��ή�V�sh;&�۶�Dȏ�Y0r-���W�^�՝^��ՠR���iH�ۏ@��ܾm%M��f� �ou���_ ��2����&3#�:���=�ڴW��=^��9��1�A~S"���;�k@����[�#do@*zcň�ȡZ+���n_ �Yܾ緘�����SJ���C
(�!�
�)߹y'�9�@�`��Z\�}�]��H:�8 �`�l �d�8 /�v�Tu'Y��w6��&��rK���ܻqd��vy�
�7u�,t��!c��5fy��s�m��;{'7v֜��Q������wV°�=�e˼��87G���182o �8�v����/���:�b�_6
���r���ؠx�`؉�RO��K]������|���>p�,�u�ںٻ=Ӭ#�����b��?�-�>:����d������D��19|V�����=v����k�c����#=uY��F�ށ�Zց)��]�=Ş�vbl�	��=�]�@�czWF������Y���`e{<^eh�ށ�ѽ6F��ڴ�U!�~�)q��z��:��]�@�z��n6�"Q,�QgE��I��TJ�s��h��R�9����A�������:��:c}$�~iܾ緘�^w/�T��};�^j�Mj��5I����9�}��*� �$(;DԞ߹�nI��߯�w,�_5UU6fj`��i�)dje�h?נuto@���Z!V���!�19zg����.}~z���y�h�W�{^�:�̒�ґ�Y��z�Z+���z��fY��6��R(�x��"�3պn<�Zí;�m�
�
;Z��=;�-͉��'?4H�=v����W�_�J��3l; z��e�(���E��^w/��g_so�fٛ|�o1�U*��n��f���#����};{�O~���W�2����rOo����ňQ[��0��\���UI<�f� ��Ӏu�r��S��m�r��q�A~S �AǠ_zS@�z��z��:� ��W��	H�m��YC7���ڷ�z��m�9�x]�@t����k��x�"pǋ����9^�@�ޯ@�ί���gƁ~�B��m"n�w%����_6���6fٛ|{�M���^�:�̒�ґ������7�5ѽ�^�7n9��q~h��ޔ�9^�@���7 ��`�B"Ȱ�E� ��H�H, &���ُ�:� ��匓"2d���%1�����7�=14�=n֌�$��*�=�]I���gVH��&h��E����ꄆXĚ�k�YZ��7�F�ހ���%1��ˆLjb& ���&�՝^��)�r�^�y�@�\qE_��,X^^��14c��.hdo@���Sg�����z� ��g ̳�|�J��s�p���.� ���rh��4Y��s�޳@?}���l	$�H�rHȉ	:on��En���e� � H�M��  � K�\��e���]n>u�l��+g@ݶ�}��������)�����Xѓ�9�v^���ޗX��;sq/Kv�j�s��2n9�g"8��4֚�k�������{gun����v�PtogviAK�[g"���F�r]���4Og���]��V���ۻ�����ͅ�Iy���_�tu���Ϟ�o7X�{.��f셃���3g2g�3$�&�p��3��=�}V�[�h��h��s�������~h��s�h�4���ހ}���32#!K&
E�[Қ�u����9�Z�
�Xa?F��$�4���ށ��ր�@�_>0���&0qɠZί@�U�[Қ�u���\�	H�m��ۦ���ʛ$����L�$�0�[����ر�P��L����>�@��8�{����3o�n�u�_i�ɪkY��'�{����l1}Uf���4�>�@�U�u�kSA4�$Ԇ�y�f�n>�O�fg佮�����@����5�#I4qƴ�ƴ���h��z[��&�50��)��>�@��4��4q�Z���������$JF��zla�
�jچ;�f3�y��Օ���n��I��Y0R-ޔ�;��-W�x��%�v��{l�"T��q$���ݏ�Z���Z���nS&51L`�@�U�w�ks@��`$���B)�*��,}V�w����㈊(b��Ab������-}V�yz��b����7u:ֹ*�LR��;��f_q��m���� �޳@�7Fؔcj@����м��(�6��y�k��]r�]�n�p#s�8�t��Ͷ����|}q� �G4�ց͔J/�]{$b&�h����4_U�wY�{�=�vbo�S	�b�h��p��>�l�3g �W����,�I�ȢYRM��h���-���rq葂@H�H�W@�*T(��
��ϻ��'ݲ��wS	�H�MŠ^�@�U��Y�Z���b�*#�)��M�I��0�,t�և�i��N;gg����f�����ژ��&0qɠ[������-���Ix��sg �o5Yq�:qA�켭 ���Z����-��U�?<X������-�M ������ ����Z��4�$Ԇ�y�f�n>�@;޳C������h]LX�|���0$�@�U����M ��hz~���w�{ǔ�")",� a�E�!a[m��`��� F0���@�UN j�X���C7����$.��c�J�z�"�i������#��=a}OI0	@�h����b���3$�F!#��zAC�����7w���;�����;����   �`         T�hQ�R���P$įgX`��q�͛iNѩ�s[����P*f�I�#�8
�*��(��w&X��     �      �       d�   ��m�       	�m�        l      ��     $�h�&�Kz�V��8$�4�&��m![ӯTݮ�`��	P��a�S%�8`,��b�l�9{Wmòq���ێYv�y�\���Ơ�8�5���u.6�u��C�����VR�f�
�J�q��݁��cM�X��v��v�gps.,Eɓ��kU�8���M�i8^x�N(G���V��Z�
wI286DF��[v���n�մ��2��>s��s���OnzTpɷ3�;�o�\| B���;0X�P�m�Ռ��.�<G87Nv�����n9��N����7�<W9���]pu��Ms���Cm�ʖ�dpA�n{v�*����<#�����v��nُ�ci�5�VMr��/χ����wl=E��C,c���z����^Q+�im�U���UWj��g��쬲tG2���U`T��j2�(v�cv��˲ގz��<į%�9�<|�Wǫ����Z��{p8�Ղ��i��s��`��J�vQ���ڳm6�;�cfQ��K4Ѭ ���ላo<�Q�Z����  G' r�F�.Ұ��W'd@�m�NnÚ�N��m�s�}�J'l&�J�"u"[;N̚{H�Kmn�[N�$�]/(8Ӳ�v�n���C�Ѯ��W�i��񇎍�]r!Z�J��Q�/"�����!������.-�*ݱ�6M�F��i��s`��3�iף���ۢ�j�����pR�4�T�i��a�k��DS��qUUV�t��n�C�j�9����|�{���E�� >~Q( >���֗��^��T�p�@����[UU*�@�]�#���I/m���@  $   *��.�	�U�XI�F�Dc���M�ag��]�-Z!j�9ݼnSb(㲷c��Ղ�x��q&�d�E��G�>Zn�23)���ll��F]�99/e�ڶ��Ƕz�<m�n������܃�Gs�ml������nΈ�tv3Ga�ɡ�ZP�	����������
`������\\�����=z�������[�,�n��X_3��b�|���[Қ��4q�Z�u�&�"�dII4zS@<�f�n>�@;޳@:�V���2��� ��h�h�怳@�r፩���c���� ��bh�s@�����VV�Ab������-�M �������|�cxB!��x�K�X���ö�aͬ������s�;7����p�����(���NMޔ�/Y�[������:�
���ȓNbMHh���I6f+�> y�rp��9�;�'�#2<iL	$�>��h{�h���yz��Y�s��I��	�'#�jUUI�s6pܚp��'URI���[,�)ڌrN �@>��}q� �G4�VU��aY"���#���m�����7i�]�v��S\�vI�toN�� �G4�ƴ��bhy�p���LXL`��@�U�wY�fva�;ܜڤ�g�y�Ȥ��MK���l���p�T%\I&&$Qa�AH�x�T����N���>���5�V�q�qٗ��,���s@_\k@>�����h2$Ә�R�u���� ��ޔ�;�*�6����N
�u8���k��n%�L�I���3�F��!8F8��<�̏SI4q�Z�{��fva����l�Mue�$�\������'56n�Ӏ�l�-��h��,d��B%�
I�,���s@_\k@>�� ��,2b22D�N�u���� �����6R�"��D��$ 
�5�As>�M�'�{.ژ��	�rh����c�3g�n�Ӏw�8�UIm���.�i!�q��G�lj�7\Y���ŝ�<�e$べ�%R�]��5%����1��r�f��@>��}q�_W�f��(�����)�{�h���z����h2$Ә�R�G4�ƴ�h14fS'���J`9&�n>�@<���-�M�z��Y�s��I��	�b̭ z9�,���ހ��ց'��H����K.��ϡ6��.�-�� 6� l @ �rK�i�٧I�,�m�$���것���5�݃��c��gd�w!�pK(���ZH�I6�/Z1��%�����9� A�9)1$�w%����Cf�a;c��+�j�e9ܬ�Щ���A�n#Z�n֮�͖l��:�!6+/���)g�e�7wq.t�$J��Y�nu�ہ���<<�϶zuU�\�2d�;v�htwo,��!��N y�rp�}��UW�{�8���>�LF)�,i' ��f�n>�@=���-�M �-�cjb	�)�*�3@_\k@;���M ��4+댙#Pa�d,�- �޳@�� y�d�mUUS�S5�j�)�X�L�Mޔ�=�h���z� 늼eƛR7mbR��ؽ˺���g�AR������/���.��N-\��,��dI��5!����@�U���h������<��PiL��O�3߮�5	"4�I<�ߵ�'����y�@�{��$��A?LR. {�rp��8|�6{���7U� {�ܱ�a2K"�@��4�m���� �޳@-a��d�[n��=̜j�[�f� ;���2����Eq(�M���A8�m���k��s��+h����N��[ևV%��I������@�U���h���y�@��$j�)�X�8��9�,���s@_\k@y�y=2b�5#�@��4�m�<E]R��EP��t���}��}�N��
�F�"M̉� ��f�n>�@=���-�M��1�yQ��1L��-��hfb�O ��>4�m����������(�y���kp�;�۟gV��Ts��"d�r2l0ꮜ���t֬X	Q9 =��8gf ��ɵJ��>��hg}�FI��dQ,�RM���>�7�/�5��� �%�1�H���4+�q�Z����)��O�&2(�Z*�IS�S5�;�8gf�UR)TQ") �Q �����7w$�~�L��c��Ab������-�M̾������m%O�O-���.�U嬡�]��y8�i���*e�m��c������u�mlq��ͷ����|���ր��� ��#r���Vx1&�D�@�@��ހw�f�}v���0x���?$��-v����ֵ�|�k@�W���fau�8�~�����4�hW�h�[��nX�0��%�
I�_]��5*�fk��ݻ�}�N�]+�oϒ 6�{}�Ʃ+���wM	1�M� �� �7��(� ցu&R	j$�ν�^���c<KmE&ݣzK���:�ڒ'��o3�>t�<[GIn��6���v�b4�� �N*ܓ��`9���by�TX@u˛����iz�x�<�`�zpmv�{0&�e�q�8�[v�ڻ��b7/'����
�sn)).���49�y���^�w|�<��ul�$��*���ԝ\�玒��QቧqLc,^�4U�J��gW��yP	��hkw���ֵ�v[p`��A0���qh�[����/�ՠy_U�y_\d�����˽ ������Z����ŔX�E�D���/�ՠy_U�Z�o@;޳@�LTx�I��U��h7���@'G4�k@Y�v�cȚ��F��cnL�:���l��u�wM6.��oD!�����s�
9�x�iO�8���@|���޾ ��z����rH5���o@;޳|���i:�V�J�)Y�� ������wϪ�&�ul�EmF9' ����hS���@'G4�c����#Www'j�~�wo�n��� =����@�-�0k �H�Bq��[�>�^��x�}��<^�z������U^Z�/gͻ;c9j�Np���&i&$���W�ņvu-�ޮ��˽ ����&��Hހ��z�QcذY��drh�)�x���-v��wY�y_&*<P2;���r�����̻��W��II���!���>	b�XB����G1P�n\%p.�b�t��|�.\T�T�Eb�F�ڤ��[t�J�I���0��EH��J������6�יL +i�#��_	h>$#�$	�l!��Lڄ�*��B��Bh�	���O8�`���@�Łc)�Ͼ���ƅ�+��
�x�.��(p�.m �L���a\H0!L_���	">�0װ$�.��W��L"σ���$�Eb$Q��Z�@a? ? ����<�C�4�=⇈�¯�� v��I$�����;��ps��l�-�#���fe�kw�H���}R/@����rL��8�~�����4�)�x���;���׋�"JG\��vQ�k��sb)��jڇrul+����\7a�m��vI���yeI?��)�x���;����3���4�1Q�C&a2E�p�<]�������4�)�{��5��L$j!��	-n��s@���>��>���'���,RF���4�)�9|��ܜ� ���WqZ�,B%���
EZ��}��'|�~1cذY��drhzS@�{������z����zV�dm��O p�R�m/��1���>z��7a�Ln43��4��))�A⁑%1�����:Z����3@�9V]�_�2����^�%�ހ=�#14�^�qg����q�����@y���mn��Ϝ�3�FK"iɠ_l��W���kz{��鋆Xd�&H���4�hkw��h8��߽�uE����Y�u��Y-f�&�ˮ�h � �@�>�UYF�Q@�M�L��.'t��K]u(�Z�h����6����anw���uoh�=���^:&�͎��[f @��&����:�z�M/�ɤ���#U�ר�]���b��W^8^{A�]V���9M�+N��	�Ϟzn�@{]MoV�փw���^�&�\c��I�ɖ�M�=�t���d�l�N�dv��3[L��)x��I�~m�_�����N����J����_ ך�RfA�S �9��f�}���� ̼˾j�l��z&����m]�mI4���_]�@��ހ^�4+��Tx�A
cQHh�j�-v�����e4:�X����P=uyZ���#��&���i���������N
�,m��tAJr�����@��=/K��g:�ꝝ9�4���N7����e4�}��<A������>��"!�D�&�����q� �DUQ���>�ܓ����Y���ɘL�cI8h��>�y�|5U6nf���Ӏx����œ	Ȓ�h]���@��M��Z.��!�d�2+3.��������6�z�����ڶH�Bs��s������q�-��V�A��x���7�;'-Wu��ˉ�=kZ�j�����<(B��R��h����@��M΢)D�"&�Awp�y�����J�+�T����S@��Z���+�$g���N7����e4�h}��}�z��g��̊%�4��<�S@��V��ڞ�^�4{OVЛq���r��I��ˑve��WgF;^@:�G��uU�ČPd�L�d����}v���= ��h[)�y��mnbɄ��m��r�.���6���{�4��j�9u�'���,RF�����hZց[��Ԟ�^�F���RM�e4�h]���`z�Z��6�����{�����(B��R�ڴ����Y�yl��ｊX�i�*������\bת�"���y��q�3�F��6��V�dc������� ds@�q4�k@�u��o�2����N7����e4�h]�����&DC"�dM94-�p��I��ݻ��l�z'�̂�HՍ�8�O{7_ ͽ۾ ^�4-��<��6�1d�(�4�+@��ހ29�|����'�{����?	 6��nܲn���m:g[m` m�@  @ �J�	K�K�K�{i˧l�2�DVS5	���zyp����e�z��&G���룙㣎f���n��[	������f�ml*��Ȝ۔�w�\cj��;ۄx�6��𵏊|�n#�{��
��'Bcv�y�7k:�v-�)<���t��n֫$�c��_���I�C���=�:<n�.���o3u�l��wHp78fuKix�on�r��Hހ}��yl��}�M�����LX�ɋ#X�M�&�岚�@��ހ=�>nU���VD����/�w4�����hfL8���9�i��8�䋁򪧛7n��͜�ɇ �{�\�׫� ���	�'��Y�yl��}빠uv��_{e����QF����^��a!�a���-b֌n\cN&�5��g��O$�&D3"�dM94-��/�w4�����h���,2f$X幩�'�{��� &�E?�WY>�n��w6p3&�����MDG+�uy��#kw�G4�@z;���W��,P�qA�r;�}J�����h����/�w4V���1c�DԶ��rN�dÀjJ�{���
������h�<�6$�n6��VR��^��Z�<E\�n��~[��$�<K�����Țx(<P �1Ƥ<��@�mO@/�f�岚�D,R�b2&����4������������ܮ䑥���~�����h[>��U >=� ����ٹ%���z�{r�rdC2(�Dӓ@�ه �{�\�y�|ʕ*o{�8��>�L�d����}빠uv��޳@��M�q�VL�8�Q���%.�'	x�����K�#�#�k�3i4��z��d�ڙ�&E��&h]�����<�S@����9u�q3 �)�^�feh��.&��w�}k[�J�$ٹ�n��
0���wnI�3vi�=��Zր=�#r��%��A
c�Hhy�?f+��hqڴ���ܗ�s�L7VP�J��$X�Qe�*0�f��t�b�# �H$��@C3_{�u�B��K�b�8hq�Z ��@d��>\󞫿Ugab�W��=�=;����պ76�C�4q��a�*�͓�7U��m�C/Ͷ������h��mn��G�z�=YK"iɠyl��{�4���=̜����l��F��À.mn������>�v��Qƥ��8�O6n��{�8���U$�{��8<�z�r��rK� g���Ҥ��IW��i�'~��I<�=�3rO�QEW��QEW��QU��QU�����"�*��(���(���"�)��(E"�*
� �E
�T`*A"�EU��T��A`�DA* B
�PX��*E �E@��A
�U �A ��@R
�T �D�X*D�� b*A��H
�D �E �A
� �� *F
�A��D*��ER
�
�`�@ ��D@����
�B�����@"�E *H
�X*
�H��R
�B� ��  *F"�`�@T��A��DT��AR
�@��@ *X
�R*�`*H
�X
�
���E
� *Q��AR"�*�`*B"� *��B�"
�`*��A��D�P��EQ��AH��
�H
� * �D��B� ���
�`* *X�,
�X�"
�@_�E_��E_�EUz�(��QEW�(�������"�*���(���(���H�����(���(���b��L����*�
�-� � ���fO� ��   P (     $T�    ���       (� ���$�H��*ET$� ((@R�
��T��QD@� �ID�� �    �    Y���Rž�w�w������<K�������om9t�A���@9��8�)��   ׉�ێ��><�����Qvj���{�(�z�F d^���� � "K� �  ��� ��xn0�j7>�O9��� )���0��^�۽4v�gv6�s�� �=����W�����U\{���_G����>����NZ�<v����@����^�y5�\�r�^;v�|=� ����@�`
���m��i��4QE1 3��J8(��Q�((,��M�Ҕ�� ��Ҕ� ��P ��Ҕ�JR��F�)Jce M��QK,�s�r��1���,��R�YJR�YJR� n !@ E In�(Ҕ���JR�)J_q}�g>�R��'���mžoi�׶]���k�Ix�
7{jr|�x���9�Z���>�|��｝o��w���z�� o*gn�Ҽ��}��ܯ����x��
   (�s���Ҙ��m͏�\�^�3�>8 ����Z��vU2��W9ʞp�򼸺�95� i�#����_{Ҟ]��=�u_o�}������th������j�w{��x�<�U� a$�)IQ�O�M�I*�� hh"x�T�)��  Ob�P�D�d ����j�*� �jJ���0 ��?�����u_��������Ǚ*�c��
 
UO����Ut(
���B ���b ����*�PN'�,~H��Lf���5���ה��1��ro����e1���F�L��-\@�\8$R�: ٣Z�S�e���Q�
]Ѓ�W���� x�B��5��<���7��G!HL������c����AG��O_$�= B��C##!)�<�����p����|>!�h�ڃ�=+�Fk�ivG���D��hF�"��� "H!B7B�kGX�\� P 4rF�AkGؒ��T�$M`U�HI�L*�0r�l�cs
9�I��0e,i�J�p�BY̡ytL݁���\5��M��-tR�L���֩f�]�@�	! Hb�I��S��h�#��"8�@��yu��/ɛ9?�<=����۪��]�#qѲ�!L��=�����Q���(�6}�1"Ů.��텀f�#�e���P�#�I A�0bR߾�r���=��yO����xD��f�y���)��>}q,.��s�S|�$��a�X� EThМ�߇�y�6��oT���r瞴`c�B2��T��=ja�P�X�]a�BGy��3A�� 6v�Ȕ��7`$����ĉ\�U2P!$!Ro7�����tI�=)�̻׌�kZM1�f����"1 \���)(�4���d04��$(�$���Y�
�&��H�3���y�4]�P,X�O`V4	c\�v[a���|���􁠒�!3 B�oY��2o�Y�H����Y%XS�@�H\�[�����"R�1��a,�!���f�a0�֋�\)�a�������� �*�&�p��*�D��:�"M2�W����P"�� @�A�
1$I� R�7��XK�p��ݬ�8��bS�2/4�:ǐ��Cd)w�&\	i)Y�ɐ�NR��*)��vP Б��`Ih#���Y���0dv�z&
��bQ"݃V��$B���H����,�B�<$��CA$`!k��`��>�@Dt@���I	E$ �CCD�F��@�"F�,J��C�*A
0$"�z���͘oǇ�|!��| B���ec�s/��@@S�E�|2�l�iHZ1�T`$G�\����!EĒ$HC8l�4���#�bk�������������«0�"�/'9N2����*J{�5�8�)���+�B����A�#q���H,�]5p`�Ǝ`U��C�������&4R1��s�E=��	Le�>����I���g�|R%BB6{��4l��2��[I�<�f��M�x|0&��L���<��n� ����hb% Ra!���c�h�=�)㬍��1�8jF�Hs49�vBB��J�:��o7O.�|Yp��L4��h��1���I�c��o��ɚ�j��C��<h��[-��H`���P�i*F�"�WN�y4�h
������1�1��i@��h�
�kep�4�0%�拠�}@�4�D��S
c�!�绿��<��ǜ������1���!�Ga���@(`1����H����A�@�
F-W ׼|��r�y*SF�ro��s�l��<sbz@�@ R�<<&i���]�{�{�s.�O�-5���h���aL)�d$� ���B/#� �0ӆ�xh�,hH9�6pׁ�2$$�35��8�a�����e1ӳ���$���x¤+�'����0!�C�j�(B:���{)�0,��$u%�1�L4�$Jc��b�d� ��@�C�"�J�i�0�<���My�I�k�^K��y.CÃ���(����J�=u)!kWe�A-���	���=!6�zx�D��BF��X�!q��X�)��b�.�\5s@D�J拚]L0��;J`i�a"B\�a�Y4���=#�b9���Ab�|9Tن����ĺ� �
5L�@�.;qo���?N&�'�����57��9
��Z�z�"WN�fx0�SFW�J��bU�B�Z��5��ɳs�ڛN%0�q!O8���ƹ�r�5�E*<�.�$a �J`�djb���zf�$��q��ĉ4bA����D$�!���1<cp�3fd��(a;ɜ� ��X͗9�=�����xbD�!� D��>�ޛ\�B�-�~�8yZ�E�>�q0!�)��`/�� +�*�H 5U\���2��Œ8r�1�y�k7�1�t��!��'���i<q�T���,rQ�V� R@o�B>���',�}����Pb0x�X� �
}��IĒ$=�!"D r��N��<������.sQ��y�}�m��D�O��F<J%(��
r����珞{�P�35��B�|8K���OC�5"���H�O�,BJc���G�;ǆ�S4q�h�Jc�ٮpq�3HY �$ y�� ��hdX,� X�5d|�qM:20�i��4�k��� �"�A�@b�@=��x�R���@"@§�X�H�&�"1b2	Y���#~8%Yl�1J��K$H�
�cX�
bbJ�M�.t�Hz(������aך'=�g���߮��<�p��@����cO6��S����)��T���4B�H�FB%L������n���a)HD��]0�yy��0�	p�v��lxzG&SRЉIR4�.���a�6M��Ls�_a�\5�T�#N$K�ă�#�x�B�w/1c\)����
`i�T1Ip��H!!s)&V!!`߁�����L�z���}����P��nkg�,OM��[=%3?c�(B�i�pѾ_=�o�|n&z�D�$b�EX1O�!�f�[���$��
��F��Ml��l�6�I��o�	��ߥi3L��
�B��槾��,by/����K�rpɻ�u�Z�E�� `��C�sz�#6��v`E���I�d�\��fd�L�l���8��R�6���5$�f���7S�)�炨�Ņ$dH�p�]��(B��:-�:ɸw!�R��Q\�����L1�@"�A,caF4|u7�=��&�zz=#)$  D�!$D&.�)��уWS|�T���}���}�QFj��z����{�YEg���$O_	LH	H�d!�N}N����2��I���tZ��c�YPtQR�j4ĕ"-�t�!#\p4�㧃��A٣�#\4l8i8>2�i�aLM;Rq�yv9d3|���l!#&�X@�N	�G�b���䎍0��p��9�P�FM0�������1���N�,�3M1t����a��� ֘j<���<ߞm���ye���sD.��3�ۙ�4}�<'�	�Ð�0K���}B@IG�'�
8̑%j�u�u�qG��1�K�� ��l� �[G��g �h]�h��Ԓ$$� �Fu�pj��h	 �m�                          �                                                 6�                     ��                     �               >�          	    �                                                   p                �a� �  �(                                                          	�        `|                  �                          -� �`��H  �[� {l5� m�� m�'@��Z�a&A#��� $� ݶ� � 5� m&˦�l�ʠ %�� �u�]Fԯ]v؜c���36t���JHm�����6�]]@l��)�WURДԤ4�M@m&��m�n `-F;YCt:Y`%Z�H/7�ԫ��V�.�R�WWA�TpU�����/-iU��H� j�-bm��[xrڗK�( �f��fnm�` h 7mm�i�Wi3�Z���0��m��\�   ���K,�֭��[d��Q�À      $��� 'X�` ���e���^&�mu�t��4\���i;I$ Hm���i�V�6� <�Ͷ-�H��m   �>�`6� ���nm؁,�*Q_+��|��'d��XY�� H�n�H ����q�iU�{J;zP`t]��UGg��8��t��Z�[vk4�[x
�Z��e���Ɯ��ꔶ'�,�-��K'қ:r[m��S٥� 6���S���T�fl�u�� ���-2-�/N�5�Ɗt�	�kY�5�m�+�� ��ܮ5��U<���Ih���+�ڕ@6Zm�m���ug.ˀ   l��q3J�]�:��v͚��U���������nیK�/@��cr /[m�l�f��m�L�0�j�Xsj���6�UR�+h��ꪕg����k�sm�M���}��pthS)�ν%��6 ��(�m���ճI$6[�Y��e�݆�;J�4v�-��	UӍͶ�g:9!�mg1���նBv�U@P@���UUUJ�l�61J��0Qt��@\��UR��euY;`�m��i�l9�[m������T�$�36�䝵�$�v�ejU���ـ�et]��-��U�-�8$+��U)l�+UP$ M�
ڪ�yY"h
����U�̒ʽS��s��oN�v+"ےm�� Ȗ�!������askml �؆ÙjP���mX)�k3 m&���[�{m���U���X6�۫��UU���j��������׬`-����'�+l�C�k� ��� ����-��}��}�Uu  @�WUl��.�ְq�ěl�d�2�l�rNjU�� d���^��pl�-fEܴ�R��v��6�����<Z݌s����=�:�]��Ҏڎr�gN�&�R�n��cb�X�[�A&�Y:W��i9�� �I����FcZݱS]$oA�ϕ��U�*�kivZ�8*U3펻R��im�M�6݃�WM���fB�I�I�ڶ��T��o�Z�޼�p�-�qÁJ�A"j���l6݅��R���֛`	d�j�f�6�	H״�m���@��-  �M�l ڴ�@dm��U�h� �Nݛl� �cm�	1j���iS� �f݌��-H[v��l  #m� �YE��ڶ�����vXq:Yeeh�8��   [�� sm��   �F^6輫V�� m�K� /[��   C�p�V���X���ڨ�e 6�[A�K!Q�2"��m�����pm�cm�,��@m�sm�icm&$A�u�o]�VI�d0s�����I;[&�-��ק�}�|���m�-���Hݱm�J[�H�-�콰CV����P���S4u[)E*�*[2����c��
��@W.��n�V�(/*�W�}��བ٪��S�X�Ì����%t�m���$n�*�ϒ��<�WM�zj���3�ӓ��1nk����Qd��:������q��l��6H�㾏��;e��<p�,\�p�Tmv��+,����P�;u C�ycb܏OeJ���+V;x�j�)�,U��	�mӥ�,ʼ��,�08[�g.�$.������]���U=�Yg,�hG���Dk�̮F�m���@���h�
��!̷�筕�T�Z�4^p��  ��Z��@��Ց0
��`*�Ie媞L�qBN� �f���`9�����"��J��vǬ��nY���A���p5�:5���8	�b�k�&ۣOk�-�  m���ۃ0�U\�7�A�ݶp��i�j�MY!c��˶�}7ޕ`+U-�ղ����:ک	��\s���PJ�mT�U�5��Y��k�;�U�]Kt�8/h��qKʀ�c\��ܵTnv����Ivi0�J�
^�
5�
����UmX@�T;n{%�@u@A��j�vA�	@ ���UJ��m��W7�x8��[�kX,�F�ePUe�YW�j�ΐ6Yғ���+[�YFٶ$�`pH�d�l�W�VV���Hr��T� 6ۭ�l�`qz�m�8	�\� ��i1%���l��6�Zl8��  �il�����;��X\f�Wkv���,63Pn�U�8[nA���V��m�k5��M��"�$��[d��m�p�F�7W=@��K�.�v�­�8)����n���À��g�kM�\���B����J�\�=/l�iWj�*��d�Z����U�e%��$l�$������-���A! �ؐh-��l� 9$�ldt2�R�󴫵Z����H�[�V  �f�Q��V;R�fjW���m�m�����-�"d`�fmrY��	V�[^�am 8גi��
]�����YW�����T٣�ت�W&Uͦ��%�2T��UR���h � ���m	[v�I(IoY$$  �[pmm���  � ��  Zf� �N�����6ձ�p ����v��` � Ą���$ -��� �)2��Tkivs�� j1�m��s���.V�  ?�Δ 6� ���l�A�����f��w��E���I& |�x�+`:*�Z�j�^T@m�ml+��  �.�ZL,�@49j�N����U!6���MVF���6l  �Q�m��`i6�V��\6�mݱmm���� m�� %���cͻa�յ�Ld��  �on�[F�KNm���m �i-�Ү�PZ,H���,��eI$i8խ��M��N -�=���;mo�m[ $��D�m�[F�f/[n��Zf�8�V�mp�W�t[���#�sp�6ȁ�u�c�b�Q;�6硷h��M�,
�����m�F�����I Q��[7m�~�t�|�� hH��%$����[~ N�����m�m:�VUU���*{<i��k�m( Ŏ���m�N  h�:�k]�k��p.�«����-v���@I��\6�`�d���[�m��m8-:�m�m�6Ȑ�3Uyj�X�U��]��F��Z� \m���.�eU�r^�:� 2m��mk%B��*�*��i".�k�&|�jL�h�A�lX`�@  ö�Hj���f�VY�4Fy���Nמ�j��
�E8���=%�ql1�G    @ p �m�%� m���e�e�U�`   ��]��Zl� m�m�;m��bl�MH����m�m�����7m��  �v �h� 6�m	 ZĀ}��}�4V�IÁ��p 	4�����7�������_��j��U~~��P�����R!∭7�j��G��~Q@���P5ňD�$�11���x+������AO�4����@�"- �~}���
B,"����=�
�e򂡋DV��@�CtP	�������|�?����qB�(" �� ��٠@��5D0�sBO E�
��I�E� @�$D�A� @�a#� �B0B,0!4�)�b�q � <QB�(D�H�	���j�T"
��a�@���<_x��`�@b��A�B,�# �H,�}���� F$ �@T�T�b�@<0"Ea0 @a��� A
��:Q��� �QN
��Ă� �(AX�  �
F�_N)��Q6 �G��AU@�T�D=��<T}Z��+���*+E*�
@*>���IAU�4 �T�Ȋ�60 �Uz��(/�� `*(��gsZ�$��l֛mh��5�5�    @    	    �   �       l m��         �  �H      �`    � 6�   ��    H1,�8�X�����y:b�#	��5r���*�c���G��v�k,��Fiz+�d��w�����5�� ) ���=�*�h&E�U���=�4Ṅ�/sH�`�랹��m���GRf�l'v���g�y�c<b�UWa����:��ْ��S���h�������!���Mf��n�3�!^s��ݺz�t���70��K�vҔ�d����	��p�F��Į6�A�nDسE%�a�6��ΜէnE�2N������2�t)b=�m&���2���V,���#9n�	Eϣ�6^wg���c��B��n�nF2�lGU���0�N�j3�;Y4;�r���uj�����̼\njS\����H��^��������7"C�v�Z.V�l��z�����s8�ے�v�)��ZWE�m:�+��U��K�;��\�U���	v��롧g�]vú÷:�a,1�r���mm�&J�NO66�n�gz��=1��c�N-#�l���"^�sHt�#%;sc7\[���vC��ܧM��Gkj�5�]rm�Z髱�m:�	�+��G2	i��d� :��g�]��dY6�v-�m��cq�V�l�UEl蕁4M�nɯ^�%���@HM���U���T���eAˢ�b7kg�s�=T��wQk��	�`H�2t����9�+�;m=w�k�]I�.$0�Nvm��c�4���	�e�v��<���.�B�D���F�w�z� {�Ε�a����i��ݸ��i�k�*��[vmgLI:$����6�V�`K�[����ܱ�A�(C �{� x�ȴ =T�	�PڬTj�=��K�H@8hmͰH�:@ ձ�U�\ۢ��l;t�@��nfx,:�УGkk�:�v�695k�yޭn�i��LUyxcw!��#���(m�6�ka�c��7lr������]�Kn�oT
I�����AԆ�=vV�ut6����9%�[�
��X�#�7��$���`]S�h�����v	M:�Sj9���̳$�f%3��g;�d�󓳌�e����윹2��v�NȞ�~%=㘀t�wk䘀u+!t�Ɏ&�b�$�@���wJh��@�[^�s�HY��D��	�@m�䘀��1!"�9�6a���B6�8�r���mz���wJhW�*27�8э�$�@�jBEH�� �I�9��B����:��(n���GZ:h���9���Tk��z��������������ܓ����c����CA9�wJl��̡C*�P�����'�ݖI�9�,�α��I�L�&!Hh��@>��?%�����m�� �a�,l$�i����@�jBEH�� �I�ˎ��1��XI�Z[��wt������٠�U�8��۩�j�<�INn�+=�a�'Yh7i3�I��t� ���Ȇ,��d"Nc&h�S@�mz}l�--���cl�+��������zנZ[��^�M���md�"q�jI�W�z����UU�����M{�I��_,�p�`F&��;B����N�OƁ���
�k�=����LRb�
0��i� �1/������?9�~(�0�@5���UϐP�4ۀ�b�W\#6 ���#YM�ܼ�P=�1
C@�mz^����h�S@/u�<��s�9�W�������̒��d.�a�"j,�H�Kw4�)���į纬�w���9_v"�JbNK�Y�� �Iht����C"� ���a���
1c�Wj�*��@��s@�Қ�:���"Ƣ�6cv.�j��/hY�	�6�l';��BbƋ�Vt��ؑ����rE�N��$�T����̒�{�VJ�7�Dܒ=�[��^�M��hzנ{�Սܘ�`���h�S@��Z^��r�hW��0S&1��4�ՠU�^�in�{�4�X���2F����Z^���@V����'s&�$�b�O�ܰ[^`$�p�  � l.� ����km���/4լGMָCI��������S]�-��eU+�g@�6_[2񇌔2�`$n����GY�q��]���l;�'2I�9n��h���vɮ#&ix�N.^�k:���mq%��3��ɬl�GDu��ҽp��Uc[�8��C)�#�u+>"*�"	;Uu�$p�^����.�w�"�	F࣒J��g������"�d{uYW�N�{Ku��H횗�9z4qu�E�����ʐ��̒��5?��W�2%&0rf�{�7���?ߖ�~�ߦ�in�w�f\M((ǎ8h]�@/�������>�-y"j%���@/�������̒�{�VJ�7	���$������:�V�_[4q�BR'R&�Cp|�ؔ�]+�Fxi|*6)�g^ �v:^���9��L"��Nf�{�4�ՠ���UU�N�ݱd���%lI����`EMM�=�>���ׄ�U*
HAi(A�F�$H�
E7�>޾��}N�����b��#o�y�ht����R7�@9�Z�Ǖa\D��`�E$�--��/t���ڴ�٠_�tCĔ�4��ݤo`�s$�:M@HH�m�������K�^�8��<j���q����Ol�Ҹ���U��wn+eA�<q�@��Z��h��h�)�}^\���5��rE�[u!"�o`�s$�^��U��Lfbq�%�se�$���l�;UA%]�@>��ݎ�n�C��E�!{���@9�Z ��P`���PV$�Hd�)�k���@�YM��4��R���"Q2(|V�=��x���(�d�ȧ+�뵞���e霑�I7��x�6�z��h�fK$���t
�N��vI���GY�D�2b�9&�ʫf��ҚVנ[f����*�HcJLi'&���	rL@�jܹ5 Nu��d%�Z��6N���w]�Oۻ,��կCٟ����ϟm4W�F�E�"ƛ�G�|��@�կ@��M�k�;��P���6�p���}��W�[������6����Q��9)�fs����Ӧ"&�������@�빠Umz���\ucw"�,"q��w4
��@�[^�ի^��<�\��`'3@������Z���w4�X��$ȓ�ԏC�������d�ַ]�{��'EP^���x~�̙"S!1)#�:�k�<�T��$��Ɉ����gI������ 	  v� �UWW�d�q[��d�BdM���4��)�d�i�vW{N5�<q��@�\c���m)z�d�XrO<�p�[9�v�Ht�X�F؋��fБ;��eލ���<�Е%��Hq�v9	�r� t��ڻĭ��hd�s�����V�ܳ�gn�[���j.3;%���*]�[45�Ϯ�ߧ��[����˘K�Ț�Ň/����b��4�G�;Me���?�hb�D�4��$��:�ۚVנ|�נujנ�f\E�Z��$Iř�� ��f�Nk_�=��s@���[X���4ܒ4�Ɉ2��7 %�1 W��eb.�DD�r;'EK6-�d��~��*���ֽ�X�ȇ2D��=�w4
��@�u�@�կ�m�����!jH�����9^.ȯ�F�×(8�ݹΰW[]�^�C����d�c�	��*���ֽ�V���s@�a�qcxI�&9�����1W���[U�]�eɈ�*@K�b��yr���"�=�V���s@����Z���D1\IHcJLe�n 9��.I�[�eɈ��l�+�j4�,rL�*���ֽ�V���s@�e�JD�Q�t]�okc+`�����x���S���m���sjs	�#k�	�nI���^�ի^��빠Umz�z�T8FDdMG#�:�k�=�w4
��@�u���RG��ވ���a���=����>�}�npҷhCձ1<�dM���"�h0��+�`C+�(%+V����R����Ji�=���6d$�$0�%�XT�}��˂\/#�tV,!V4a�u��C0�(l��	��P�Qb�BT��ѽ�6����+ D�pN@�2��WP���J$*�����h��f2�O`,�H\BH�Xф"�aXU�!�5r�&�K���H�!q� �LC�a@��BLp��	-��b��
B�ˑ�!�	Qa����v
n���X�Z!	��
�c
b���lh`@ �w,n�IsBݘ]���F���T��$�f���1e#HQ#D��^c� �ԤB,mgb$(Fe�a��K���\�d˘T���1bq�f�T��C,��`��Wi�x�6�� ��@�ER"4A�E>���*A���}}�ٹ'�e��܇�yAX�ĦLF9����k�>]& ˓�T����WY�n֗�̍H��Z��Z�w]��k�����_�Rg#	u����3]N�1��9��0�չws�8��E[<��Go�F��)#�:�k�=�w4
���g�fg�<���@��b�bJCRcq�n*@K�b����rb �+2�2���Jb�$��k�>]k�:�k�=�w4�˕��<��A����& ˓�T���V�Q��O�"�������$=}�%��2�6���Z��:���k�w9��?v�!jH��[�����!9G��,J�팈��-t�h�݇��I�hͨ4����7 %�1�rg諭�'5��d��Ɠ��P@�0"�I�$��Ɉ2��7 #(qR�� �s#R=�ֽ�V��n�U��=����"S�$�@s.L@>�R\�q�@?��VT��,��O~̱d��( ��|$�nk�OV,�d��(�:gJ\�p � H ��%��  N��t��U��[���t��z͂��N��vl�Z����d"sZ9����ы�en��v�x^<��es�#m8Gq��t�7s���f��4q��^��]u��Q$ໆ�f1���y!n�unL*=�ghD5,{PЙh�{pO9�f���Ү���g,�[+SR4�RB��4*�Vl�p� �X�-�������J�S�t�I��o.s���{Mf�ݙ�U�yۦ2H\4���-�؀�bܹ5 �EHL�SF8J���rH�޼�~�$qjݚ~��s@���=���P�LDoqh��h��h[^���Z�:��$�1���=m��*���ڴU[4�+�x�Ɉd���Umz��~������z۹�\�J��j8��d�X��&����r0����ֶ�4�L�ԐMl�:Θ��tL�i̍H��j�9Ul�=m��*��翞\�"D�8%�R-�Y����e_
�g6�b�:��vI�^b�� �H�H9	LB�p��rY'��~��*���ڴU[4��ه���p5#���B�k��d�Ǻ��Ջ2Y?����O�ƍL �E@bi�$vI�^b�O���������N���Ő���^��J,Q5Bpo&.�ݜ����ݭk5�Ձ!�%�"��!�%�$�� p:�\E����Q��'W��,��fX�*����-�-�c����2L�!�.'%�~���͟/{��;��VI�ř4�+�bS&#�M��*���Ͼ��"�B	U��("�DB�`  � ,`�)��s/o|��{��ܓ�a=�a��B�p6�vO� P��o�VI���K$���,�P�����y�'�)�(��2�H"�VI�ř,����un�zs�h���MH�CqHa�M�.��&��6m�;r�gn0T�6G��s��PW��m�f�	��&�r|~��s@�����-D�ջ,�st6�:�eF��Iř��=M���+$�����~��� x�|Ǉ�)PnI�}�O$�b̖u-��Iջ�ZI$>�����c#%HyĖ�ɪ�+I%����$�<�դ�k[��<�IPoI�A!0�ˉȭ$�fg8�Z6m�\I%����I.�S"��_|'q�P��t�aM�;{[�kt�,H4�lф���Ƌ��`���BmJRn�I-{5�I%����I.�S"��i-��q$�sl �2[n��ZI,̼<��mc�6+I%����$�<����Z;Ph��F\)Ӈ�I,z��i$�389��T�O?O5i$��_�8�]��FQLB�q4��ZKj����s�%�f�i$�2��-���o˞��I,���FT`��A�$�<�դ��P� �����$��OEi$�;��Iטq�	 Xa�[@�l�Ĳ� ]6 I�+���[��f�K�'c؜��䵎�@tOE�M�ͺ���S�j�*���9:�ۯv�v�c����4F�q�w0��f���]vkr�6.�㶻M���=;f˝9{t�Q��q�l��u�P,b}�O[�݇�&�p�)��v�CF��ݗҞ�!�����~��C�I9a�
*J V�B�6m;ME�G$\%=�+v��U����mY}��';c��B�����2��� �A�A|q���0Le�$kRIg���8�]x�E�m�}��:��B	�D�,R���/?O5i$���ey	�@�̒�S���s믵w�G�$V�$�{��q$��<դ�����6��z�Q"��@Ѫ�">�6< �HL ��r+I%�o�9ĒǓ����  DUI=�q$��OEi$��8�)���9����[z��H"���s�]�m��oǜI.�S"��� ѡ'����Kȃ�X!2d��)��Y��<�IhC&�ظ�Kw7��I,y1�I%����D���9$�'�����<�[l�nm(�'n�j��i�7呿���={��5H8���$�=Sb��Y��q$��ƶ��*��$��q$�h*&�D9
Q��NEi$�;���0
�%T(0�P�ƅ	ȿ>O�ZI/߽�8�]x�Ez*��m%��ӣ�FT`��A�$���դ������@6��������K�1��f1�䑫Iz�z�U M
���߼yĒ��=������[�@P���{�m$�5h^E�c"�$���-�����]�m��� #�{��Iy��ͤ�����$�pL�R�1#lm7��ν�9氛u�<��L�,�#�:.ŨZ"h6��  ��,X��!0�ˉȸ�Kww��I,y�ͤ���â��(P�bK_��V�Kr�NPDi�M��$�<�f�U  �U
�%�z�yĒ��=������4 kQv�	� ���i8ͤ�����$�^)�ZT �Gj)��/9�~���9m�����vڰ}P`��2�MӇ�Ih�MW�ZI-��q$��[6�ڪowy��I#�DւL�%M$�V�K33��I/�^�^�{�~I%�z�yĒ��2+I%�b�G�`�B]p�ZĻa�[����x]�F뗞G&�2��yvy�{��oW���8�$�Bp5#��I#��)i$�2��%׊a��J�~ϾI*��c�Ɋ`F1�#��Y�xy�M��T�-$���8�Kdw� m��F,Qp��D6�Rq$�j�e�������T�Z�c��[�zyĒX&X��Ba��ZK@<@{��G8�^^��i$����ĕ��BB	IbR"���-B)V��$�0��^�}�߸e���A���@�"���Ib̰�$�� V�毾I,Z��i$���~�?��ξ�-A	>m����v{/�ts�\g��pƙ��hȣ	�؎?xTQ Td_	� ���i8�$��|�Ē��0�I%�fpxxUP�U�ė��a�I/�<<�2FӉ!�s�%Պa���P� ��{=�q$����Iggqs�T(U EP I�D׉&HR.�p�I%���9Ē9�bZI,��/�I.UJMI$���U���'1��KhT<�B�~���I{f�s�%Պa��ڠ*�(UT$�{��Iy	�	��\��-$�vw8�_����A?� ~����k�m������[l��kv�tg$�!$�$�]�>=0���P'�y�x��V��l� !����OI�"@�!�=>X#0$^�<aL4P�A+����3��
c�.�,�r�<Jh	#tj�R)�H�%�O��V�R���0�$3o)*r��I_�}GA����yI]�)��|\S�7t覀׋���p�����K��4I�f9��Y p�kA0�iD�>A��#;�R��h�>��hHF�x{��\Iu6Ra���D6�i�i/�w��~�~��jmT�\���v     $     �    8    m�         l�             �     �     6�     [@    9��%��t�N]�Zg<[5�?���?d����י{&���lu��[hT��Խ�暢£��B�Xv�Z�k�n�	�f���U�יېmm����Y�*�؞��"��Sk"v�ܥӭ��޻��[st�L�%�Kq{,$�@���G>���&��ģa�,F0��`��,�h��q;o���
�';���;\n��M,���y���6Z��3��G=��ۀW��	j�"�LE)��'p���R\�m�n6�D63������ݦ�B�Ù��ON�:x6��ՠq���i��[�csH�&�WQ��(<�z��m��cuh�Y�l(�=W1���a}� �n^���j�d,u�T��������$��d�l^^^�z�k��Ǉv�p�����ݬ��R��ɠ;[��f� �5 {m��i�a�5ź%.�%��@w*]U�e�F�^{i/1ɸ�4rv� �7vЮ�
�+�lR�V�]s�����pm��O�⃮KOu��ۈ�������Uʵ�U�)�
�5�9�)j��v!� yv�,Em�N���wj�\�����猀�<v�g�n�\�lvr�v��t��۱Y���dN�
ڲl�D�u�]Amp�� �6�rjW�I����}���p �۴�͢s6�M�3� ��ɫ$��������q�W�p�<J��89v��62���N�׶tF2��l\��}�T�dT��} ��3cu��]������3�<Y:�d9v��v[0�ٜFN�@R�m�����y7��%UW�Ύ*+�v�k��vF��ZM���Ͱ��튥t��]@K��^�zL���mB�-��ʬR��u���߿#��(q΂�@�
��"�!����Ab����w���~���[� �8h  H �6 ����vå�&�2��I�*eɓQ������/\�p�ͷ\�8�q�=9xg%��|��v�{)�[���3Y峫��q����zwXj�N ��^��\���kk0�ܶgU&@H[���:Tr��\\���1�|�dzq�n�q�[�OgR�[���0̴�ܔ�i��������{ϻ�篣e!�4Eǳn�^� �~�8>\s�{;���ŭ4et���r���w{��.>4��W����_� ??y��I̱6�U6�ܙ��I%��e�8$&\P�]��ϳ89�ުRD}�X��K�7˜I,�fi$�c����A!�M��$����Iggqs�EM��f�i$����Ic �X!2d������Tٙ��I-�f�i$���q%�T��	i$��D�d������I,�fi$��V�w���$wvĴ�X��|�I}׈�Q�Zq5:q�:;XQ�I��]��q�µ�<a��Ө���\�.MTm��j�0�Z.�p�$�����}�I�ɩ$���J�J=I$���)b���p5#��I#��%� hDI�G�y��@N Ec4AK$E��	�] �M�6֌�Y����\�]*q�5�P%%"P��,�+�$�FV*�ѸCDm��⥲�*���9o3�~�r�{�M~��m�y���z��� �//	�3��˒8%������K1���[@Pm�wx9Ē;�bZI$>]Q���r>q%���ݗ�;I%����H�rĴ���ٙ��I.�S,H.(�$���g�$�mܚ�J����$�s� ����?
B��jݫ7<�x�"�vщ�e˔��m���P#�6�3��wx9�N�P�)7�$����Ic�q�%Փ�@xU
H��{��Ik � �2[n[�ZI,}�>s@��H��<]���{��I̱-$�02�(5?�Ț���IUe����p�/��"��(���
?�# �b��X� ��0�
@B  F����5@P�ύ��%������IgB�ߡ55��f�[���o����R������I#���I���z6�P�
 ��O{�0�w<
�}	���jG�{��	8[B�V��}�O$�ٖ4�Z%"q��2Lf)����^���n;|=^sgS�z��Y]�sjm]M�닱�f���[sM�t��}�W��������Y$��/'Q�m��vI�d�z �	��$��زN.��  ��tn�ؒA 1ˎ$�wlY��i�vff%�[������Rw��	D9I�,���P}�|,���'�}���Dv�*�W���rO�f�&Am�KpY'{��>������'��X�Os2Œy�f"ڎ2��Ǘ1�*�]��-�Wv�8.�9w���O�K�N��8�pɐ�jG�u�����[w?ff|�������i��N���9�e�ڪ��n�$���d��L7��	�Бef	N���@O߿*@Knbɰ@N�R�pLp0�0(	�����
��wޞ6I�{�,� PY��I#�S�(���r;$�2a�N�T>��swlY'���d� ��b�&�G �8	  � ln�    ��h��8n�q��w���<p�[{{q�`2�p�ݼ���勫�엜���7]���u�n�ӱ�'�8�4����Ь��G�n�-p�����v�uG��W]"���eCv��&��KA� ±�c=�f��
�i�xb9#iCl�n����9��:n��3�������:H֢�֡jꮱ��cW:�8te�P3Zk�6\�8{������{l=1K�2L�!�p�[�s@�n�����_�
�]������$�����HJ!��pY'��b��@T=[�vI�zx�'��X�Oȃ�`A2d����x��vI�d�g�C«�P"��@�"�Rg��Œ}���I��1��a�5�N�j�ֳrt������獒{��I�fX�v�W���@�@�D��w��'F��>$I�i�y���H�T���1�l�m���~�(c,^��3�f���ڰ�����.���3�YJӝ�3������ow�w�p�@B��E�8�0�E ����X�O{��?fL:��5F��+�Ow}b�9��f1�$pY'���`}B��*�Se�L6I�3,Y'�̱� �?�20$Z��_��\�[�4"�1�쓿�O��<�rş��?j�� �4*O{��I��~vI=���6�hۣ����r*@zۘ�����AH���s�߹�nI��$�p��(�m�d��2Œ|,P� `$D�AH����������빠{=��q�4�jd0]X9��[��D�˨y�V�xy&�I�R��digQ�t�b��L�6�9�˺���h�߶~�$E�H � �>d���,�с�y��8�bBԙ�'�}����O�_� 	 `�D �HE]j}�����?~��ٹ'/�����U4�$I84�4����}�s`���	 �4��C�X @" �������ܓ߿k�ܒ{�ų%>ɣZ�5��˭����� ��B*1T"u����t������I�@y���TY�t��`&2�$�w���*�@��)V*�) �s��Ow}b�=�e�$��i�q4��q	��%���ʇ\�tc�;�6�X�c�˘.˸͛&Y�5���T�$T�b AH 1 �.�e�j�a��̚��`~��� <�T�nEH[s�ņ@��H@���<�r��������� !�$Q֧����7$������y���o���A��P��H)u������33R\ԖV�^fm ?����H[s&���$��?f&HCm�ZpY>� Ш�X�H+�����}���M�9�lܟ��PЏ@�O�"$��~��I��c��8�!�R;$�67 �R���_v�?!��[��s�����R���y��`��m�u��Ie�"�{� h�\��q4��D��������X�O{�b�<]�=P�����I��H������ƤI�s,_ꪪ#���d���6I�{�/@�T<(6s|=n"U8�\��d���b�� <�T�nEH�K�2�v҆[f9��K����?fm�$���,���3]�Nզ@��H@����r*@zۘ��l[���}����w�=��O��t� �� �`��%� m�N!&v9�:�n�8�u���8�ᣴ6,�ڌt%�-���G�7`|[	�4i�s��	v��ѷ\g��\��Ӄ!\�gng�܇6q�v��npW��Z�hŚ����y�k��:���֋{dz�݀��8��6ŮvɈSmfݮna����݅�����4���65��Q��#	tTE�v�6]��D��y����)�z����n�=ދ�~�z��FI��3����s@�wW�[e4������qba$1��9�˻��@W���C�����'=��,���b� �A$841��M�� ą�����r*@I"�[sWU���"I�Kp�;�� ���I���I�w������   g�߾�l�}��E����)�8,���b�?.��l���[��w5�N'2E�����%nӃ`fص�Ƭ�-�)�s�e �4��?ނ���Q�4g �D�pF2��m0?_���M��EH	$T�F.�iȒ�[f9�s2a����� �E�)���`�TC����@�]N~�7$����nI��߳�$�� �w����f���q�l����Y'32ş�B�\���߿OƁ��'q�����OF����� "�C?~���rO�w��9�0�?�}��I�A�hA2d�������y}��ܓ�Q�(�XE{�������Y'�̱d���,ME�4$!:��Y8����s`�9�U�Nݝ-����\�Q�]H�s1���O�o��k�'=�훒{��l�(~V B 2qn��$���4�2D����O;�b�T=UD@-��zŒqn��'��M �\Hb�Gx�q��;���O/����8iH�2WY��"I"!7�3F�Y&�T5 �P�	/�3�H�$X'��!҆��)FHE�@����.����J� ��T%	Y`��mm$Q$�7��f�1��7 �9�q�(��@�h@$�@ 8��#�ўx/�
)�D��~\6�*�X�x
� ����t�'��X�Os[�N(�Sq�d��B����d���6I�s,Y?�~� ��{�d�4{Y�ND�0"�77q�lr*@s�R���������CB6ƌ�Kk،��n,�	w5�<��d�D�	A�<< 5�Bx�dpM��Ҍ��Ӏ��� 9ȩ����}U�a;���N�~I��p�R��@s�R���s`��R��W��D��FHCi�m�d�[�vI��`��R���]YRffV��n\�'���	y�獒{���$��͛�� ��P��hTB*���u�RP�%-&�-�%�`�R��!d&����~����si�Ń�C�7�q���O���\�߿��l����]�%�-�U$��q���z�'�6��p��Μ�K2�	��.C��&�>XH���q6�776�	���R���s`��R$�0e�T�2�e'I�w��� �P��o���{���$���I#�:�4�IC-���?w&$�,�U P����Y'OzA�r8$�#�����EHr*@u�1�U}�j�o��d�[䟙l@�% M9Hr*@u�1�lr*@��z�ޝ;�9�{����[߼�,0�?��}� ��m��l �8Os���sx(칓=��ä�ê8ۗY��]=I��2X�yF$��u�J����F�C�j#@�N(����sc/4�c�M]�΋���	�iv]8��q:��[.�F��Y���)ˍ�d,�4�ѭ����	M�v�Ǝ�f��>�r����؝��d�U�8�:&��������BՍ	=[sѬ/b'e}qe�g9�.9�;��e���P^��^��]�UQ��9��h�m9M�>$���;$�ܘl���X�P���nزOGC��	Q��R�vI��0��I�vŒ{��,���qފ���>���%�p�3D���R����� 9͂ ��
�j8�
B�R'¨W�o���~��9�@y�� �J�6��ͣh�Rq�d�.��|(WsoO	?fm�$�[��}�U�JD�Q��$k9��^ð������|�w4n�$�ܨ
�CM6�:��IB#dr?���~4����s�@W?c�VI9��#�Hb0��n�9�l�4��X@��H� F 2�@��B�� ��*��ꪯ��1ȩ��-�l/�T(U�W�^��'	DHn$����*@y㖏�۟����?*@;(�E��!4�6�x7�{�	9��6I�t�����?��ykm�Q�8��O�Ɇ�>��g��������,�ξ�>�PZ��i���5�X����1{%�;F�@��75�]3�C��Nk�\*1�m�f�����Hr*@y���?Oƀ^���/�G� �Rf��s@��-�ln*_��%~�_�m�a�J1��pY'�y��?w&.�������hu�������IB#b�-�U[����~T��"��9h�\�ds"!�q�hw]���fu����W-�e4ݜҪF�$J	F�u�q�L���V7�z�UÎ�{v�ŵ!s�f�8�D���LN2LM��u���9h�a�諾a�~T��P���CNc��}Ϫ�=l����r�=�e���#����i�T��㈧���o� ۊ�ȩ�Z���
�Qp���������-��f��>��M�H�!��߳�h��,b��F�h�f��n��3�ߧ���;����;��h���8�Mή��kg]�[e�ێ÷.������ݞ�/>��Z�us0vK��p�w�o��Ih�`�m�_��XI��_�~��ND�"1�)"�=l����s@�b�=�&�����}�#�H#��q�P���r*@>�I�@Kp��7	N��4�N����d��f�!�e4w]�����Ƣ��Ә�ͤ�� ??ߗ��9?*@7"��~??��z���p� H � M� m� $,�^:���u���A�	���������&�s���Gm��d]���v;B̦�%������ݍIע��K\fN0��i&*�h6]�<�hL����ጼf�9��'<d$ܥ��muh��[I���N��a��W����vhX[�9���7;k�����8x�Xh�ˮ�-����un}ܮ�)3����gFԅru����B=��Fd�<�[\�س㣛��ێ�b��6����@sqR�zç�� 'β��X���{��h��hu��=l��{��Tq��J@7"��� :M����������M����ͽ6I���d��ܱd���Y��I#Fk:ӑ%�6��4[)����g�[����YMަ�J%QLD�ɈY'�GzAM���a�z�˜�=۝A3�������7����f�h���r*@y͇�Xw���Uq~�H
@FI�73@�f�B�j@�E4�73�k�rzS@�u�����EFU`���ۘ�pY'�٦�?fL6tP��7���d����s@�;uM�	�D܃N��@sqR� �����	�Y�,�3���T�nEH9�@^��|r�R'�S�,�1�&9�vw=�
�Cqu6�uG^xF����+Nwnb-M��_��s�r&L������)�{��hۮbX�?��q��>s`�U]���� �� #�R �NaZr$�1�����=�w4٦��
���lY'7&�$��1��ݭͿ�ͼ��T�rEH9�@u��.�]"����nf���H�]?/ǀ��o���H	]Y%��YK��u��ínx9�<�qc5��G[0� 8��I�5Ө��N�gMs��lM����}�	���H�Y��&��d�N[)�{��hm��>�)���;���B3�!��q`�D���*@y͂ɰ@�
�.9&B�R'�����I�zx�'����DP���*��e�,^��%�S���I��YM���[�s��Nf�Œ{��I���iC!�$\kD�ȹ�SӸ�uh����;��j�v��ۓ9��K�h\er��m����s��ȩ�ТL��݂8��p�'ﻖ/E$s7lY'���`z�M�b�Ĥ	 #$�ۙ�s�R�6�Wo��� �� %���,��&������zl��٦����h��hg�婧��7��DI�@~������W����Htߦ�_C4���lڱOtc¢D*' �q�#T�RIFA��a(V4�4�6�*�J�*!���~`~��@yg0m��Vug@    �    	        h         А         �   H4P     6�     ڶ     �    ���ۢD�m���^זi��Sέ,�ې]�gi���c��5�sv���=r�P*t�Ň��E��SUWUB�ò��#��
��.YK���{q��&�����R�:M�9�`�J-nFͼI�AZ��Qp��6�j��q UUv����5��r���9�����,��k
c��[q]�n�Ûc�L�p���샌���Cu��m�;3R��d��yA
v['l�^��瑲R��=�MlnS���mQ��) ]�����-�R"�ܗcY�U���"7�Lv�]�;Ja|���ݽ���+�؎
�V۳HǬ�n1�ax9Tsh��M���L�cS{Q�1,��yW�����fΗ��&�Y�7�<�Tr����u�G��E�t��7a۶��h��qp�eܩ��Q�]vݸ�v����ڻ�a��΍��g����S]$#u�,������4�a����&��p�b���6�����Eۂu��%�.9m��5]���Eu��m�Up8���h�R�;b���V�vFG'2l���nÚ#m��	S:m��m�ޅ���e8��3)]��]�I �u:[��$�0����1�t�1�b��+��<�,�.�Ú��$��,)���F�WN�[-tJ�v�k���md�v䀛l�g�'<W���Ŭ
��q'q�<���g�n�;���@0`�����\�mƙOj�8���c6A���
V��'��ĢL���\��4�ъm��.�Չmb�Ь�����7�-v��VI@"��Ut�W�"��IN:��E��V�K�T겺�J�� =\�V��<��)TC�*pA�~�=2ڀp � H ��6��  �g$�d�[�K'd�vz�=��j��)�K]��\c�2�/f��PQvsꃵ���-����m�{wWQ�s n�G/�:l�Lu�ݲ��m� n��.{,q)�W'�,�f3�����7c\����Cl0ॱӶ�z7��;K��g�n�ru"��H2ӋX��M���;:t}�Kj�����K��=�!��lg^iG#�WI,�f�WkA�dc�#��$B2b7��}m�@7"��l2K@ҋ�.�D�A�������YM�ڴ�w,^Я6}�z�	SR��ڊ8,�����@t�-��H�T�*S�L��%�˒+'�*�woM�{��,�޷s@���@=L-q�I���8�����ȩ�Z�� 9�?�F���Ku�]�q�i�mq��K�Pe�b�<�z��3��΋�������me�mx	?~T���-�l�T���u�&8H!�0��{��^1��"@ )B$"@`/�r$��P� F0#�OX(�`���,X�!
A D���V! �Xc� $bE���R!! �!G h�BDb0!@_�"a��'�澛����s@�s@�v<�pI��y���6r*G껟�~T�s?~�{B2�7	�@�[��w[��{��@������1eqB4H4Ԃ�=�e�;A�3&�4����}�ND�,K���6��bX��#�F7Q�v�+t l�OZ�-��DwdGv�"sΨ�n%��̺�f��"X�%����nӑ,K����fӑ,K�������K�F�f��᠍h#A�t�"I�,�ɚ֮ӑ,K����fӐ� ș��~��Kı;���ND�,K�뽻ND�,K��N�5�d�3)��7C��4�����%�b}���ӑ,~z����b�D 2Q� ����x��5�k�]�"X�!ܽ7C��4��y�=M8L�h�sFӑ,K? �ȝ����ӑ,K����~�ND�,K��}�ND�,[��ND�,K���&Hđ�ڀ��4��hwf�4X�%��{�ͧ"X�%�����"X�%��{�ND�,K�
��}��$IА�έn�Y8����Ƚr/���U8��m%6�7嚼��#`W�b5x�D�,K��o��r%�bX�}���r%�bX�w��9ı,O{���9ı,O_Mv�å��2��ӑ,K�����Ӑ��r&D�;���ND�,K�����9ı,O���m9�,K�{�\��j��ɬ�\֍�"X�%��{�ND�,K�뽻ND�,K��}�ND�,K��ND�,K��y�-fi�feֳ4m9İK�뽻ND�,K��}�ND�,K��ND�,��3q5���iȖ%�bS����܉'E�\�]�F�43v��r%�bX�}���r%�bX�w���Kı=�۴�Kı?*���?�� ����'^:�{c(n:�	q�(��ϡD��*\t4�s���t���e��W3Si�Kı;�߸m9ı,O����r%�bX��]��r%�bX��zn�h#A�zҐ�!J�.h�r%�bX�w���ı,O{���9ı,O���m9ı,Gsw��p�F�4���Y��\2$Z&\Ѵ�Kı=�]��r%�bX�w���r%�bX�����r%�bYC7w��p�F�4�т�Ӊ&��SW35v��bX��{�ͧ"X�%�����"X�%��{�ND�,Kߵ�ݧ"X�%����Xt�5�]Rfj�9ı,O~�xm9ı,O����r%�bX�����9ı,O����9ı,H-ҁ��_�kz��$�����$m�e  �l ��󫳝�h�n^���v#!��ݦKWi\r�F$:��t���t�	k�P�����N�v���3�mn�Ku�����1�۵\�� n�[���Y[�J�N�q×S��p�fB��εrK��k���s�΢�ͺ;Ie]�g�����˪tT�L�E9b(RE*X ���������G�,�����Z%7��v�zw..��/aʝ9�u����y�Oař�Y�Y2�֍��,K�����ӑ,K���w�iȖ%�b}��a�<��,K����iȖ%�b~���3E��3L̺�f���bX�'�k��ND�,K��}�ND�,K߻�ND�,K����r%�bX���rt���Y�,�ɚ֮ӑ,K����fӑ,K�����ӑ,h�lO���7���=�u@�@��cA6�TS)��W�=����Kı>�{ͧ"X�%����nӑ,K�
L�����t8h#A���|�Ґ�!J�'�iȖ%�b}���ND�,K��ݧ"X�%��u�ݧ"X�%��{�ND�,KΝ��9��kR�\��+[sѡ:����U���;�,.�خP^�;�����ڀ���᠍h#C�7U�Ȗ%�b}�w�iȖ%�b{�{�iȖ%�b}�{ͧ"X�%��񣽭3j@�6�4��hwf�9A�ꇀ�m�ND�7�y�iȖ%�b}�{�iȖ%�b}��۴�Kı>}5�K�f�˪L�]�"X�%��{�ND�,K��ND�,K��ݧ"X�%��{�ͧ%h#A��cPq�1���]D�,K��ND�,K﻾ͧ"X�%��u�ݧ"X�%��{�ND�,K��y�-$�3L�]]f��"X�%����fӑ,K����nӑ,K�����"X�%�����"��hz��xo�E)�����rX�v�)�������x�=����F����{vg9Z녘p��(��r�t�F�4�����iȖ%�b{�{�iȖ%�b}�{�iȖ%�b{�wٴ�Kı)�`;���AN$�4��hw7xm9�9"X����6��bX�'�w��"X�%��u�ݧ"X�%���Ku5!2B�HN��A�F�}���r%�bX���xm9�b>E#��D� �0x�a�BȊWBZV1��V�+	@�@Q� ��Y@�dG
��PD��Obw�o۴�Kı>����A�F��1f��bH�mBL�ND�,�"}�xm9ı,O�k���Kı<����K��"w��xm9ı,O���?L�5f]h����f��"X�%��u�ݧ"X�%����"X�%�����"X�%��w�ӑ,K�����yu�ɕ�����8��ɻt�s9�uǰ�R97=	�BX�k�9���kc3̜,}��oq�X�'���6��bX�'�w�6��bX�'����O"dK����~�NJ�F�4F�����1���]D�,K��NC���,O���ND�,K�����9ı,O=�xm9ı,N���h��4�32��4m9ı,O}��6��bX�'��{v��bX�'���ND�,K��N�F�4њ΂�&8�-�[���Kı=�۴�Kı<����r%�bX�}���r%�`u��L����Kı)�a;ܥ�љ�˚�5v��bX�'���ND�,K��ND�,K�~��"X��F�vn���A�F��F4�H҆A	F�[Mù2^˷Z �G�m�W=�{e2<q�e靀(J�Y=\�w����,K��ND�,K�~��"X�%���f��O"dK�����4��hy�>~
đ�Y����r%�bX�{�xm9���,O����iȖ%�b{�p�r%�bX����t8h#A��`�54�E�	ME�f��"X�%���fӑ,K��߷ٴ�Kı=����Kı<�o�᠍h#C+�j%1�3Z�ND�,K�~�fӑ,K�����ӑ,K��߻�iȖ%�b{�ޛ��A�F��f�Ơ�a��e����r%�bX�����r%�bX~��w���Ȗ%�b}����ND�,K�r���F�4:34�6�rI ���8h  H �6 ���:9#��g�نM�A�2rj6������.:�3�l���vL�)�=[��{C��魻A�<97�����g�tSv�����Zd��wf(�Y-�mHX喖ɲ\kNFuˢ�ێ��n�<��u�e�7'&�\z���s;rP�+��n��6����8[�rCw{�����`���u�7��N�^nM���a۞k�BΚ�g8	���ۘ�Sj��Wi4�˫����%�bX�����r%�bX����m9ı,O=�}�ND�,K�{�ND�,K�>�N�3Rk5e��&f��"X�%���fӐ�	��,O~��M�"X�%��߿p�r%�bX�{�xm9ı,K�Н�i�$�E9��p�F�4��r��D�,K�{�ND�,K�~��"X�%��o�iȖ%�b{��{ۥ!�B�Hq�t8h#A��h}��ND�,Kϻ�ND�,K�~�fӑ,K��߷��ND�,K�=�tKF�fQn��A�F�ٻ���Kı=���m9ı,O=�y۴�Kı<����Kı;���L�C�����l���^��A�7Y5tE���t%�X�+�k�{��q�������35��Ѵ�Kı=���m9ı,O=�y۴�Kı<����Kı<����Kı:�k��vK3Y�Y��Z�ND�,K�~�v�9
Ut m�T۸��bg�w�ӑ,K�����ӑ,K��߷ٴ�Ti��h/�kLkbl�Z����%�by�{�iȖ%�by���ӑ,K��߷ٴ�Kı<���nӑ,K���n�'tI4��5�Ѵ�K��2'��~��r%�bX�}���ND�,KϾ�v�9ı,O=�xm9ı,Jzw�;&a�3V2ə�iȖ%�b{����r%�bX�}��iȖ%�by�{�iȖ%�by���᠍h#C��x�M(dJ&��\][�7:����ܴ[�v�)�g�6uO��ze�VA��aIf���t8h#A�<���nӑ,K�����ӑ,K���fӑ,K��߷ٴ�K��ܘJ�ӆ)	dHq�t8h#E�by�{�iȖ%�by��iȖ%�b{����r%�bX�}��fӑ
h#A�J�đ��[��p�Q,K��}�ND�,K�~�fӑ,h��E�jwܦ5
��e�a��C��xF�$D�p�����b6H�U���
E7E�H!	$I 0�A�U�y�1HDd!P�5MIh� @ �CHU	X�Y.��j˄Q`E�]h�K��j�ZLC@K�M\�L�s%���Ċ$�Tj�ȁb@h!4b,@9C�K)��{̄31"ā�tY5�A�~}A��4�
A�=����CC��0O�_T؁��"��<��L�{�.ӑ,K����t8h#A��`�54�E�I��M�"X�%��o�iȖ%�by���ݧ"X�%����"X���{�7C��4�����t�dl��rM�"X�%���o;v��bX�'���6��bX�'���6��bX�'���7C��4���qiJD�-�*! ��qz�9�ղ�:J����i9�����۵1D�̉���M.�������oq��{���r%�bX�w���r%�bX����6��bX�'�}{�iȖ%�b72�"vL��JG�᠍h#G���6���9"X�}���ND�,K�����Kı<����K�h!ѺΒ��Bm�7C��4X�'���ͧ"X�%���^��r%�bX�{���r%�bX�w���r%���;��P-�ل�#p�
%�by�׼6��bX�'���6��bX�'���6��bX E��������F�4>Ʉ�M8b��f�k2捧"X�%����"X�%��{�ͧ"X�%��o�iȖ%�by�׼6��bX�'N��l��e�0�[����ín{8��k:b3Ԛ�E���mQ�̎�5����B��M�{�[�D�,O;��m9ı,O}�}�ND�,KϾ���Kı<����Dh#A����)6�rCt8hX�%��o�iȖ%�by���ND�,K�{�ND�,K��}�ND#A��蚁GIFF�I!�4,K��ﻜ6��bX�'���6��c�"}���M�"X�%�����᠍h#A|3Zh�q��h��Q�tr%�`'���6��bX�'���6��bX�'���ͧ"X�%���w8]�F�472�"vL��JGӑ,K����fӑ,K��"�����yı,O{���iȖ%�by�{�iȖ%�b`l�BRA�r�TVswI�D�	$�	$8	  � ln�    8��KOu'���Pw:v��N�;���λ�w!��Y�����O[n���=�ø�v�S/m���b0�^ulKȞ�\s�8�q�����pK�9P�dtْ]p��Nݞ\v�	�$ۧ��l�v�8ᱴݶ�7��m�i\��X�{jz�u�p��X�sZ�k���1�u�zt����v���aQ�$Fqѫ��.�p�q�mh�����OlA�9s��w���Y-��D&�.Ct0�F�4������Kı<����"X�%������DȖ%�����6��bX�!����0��n��A�E<����"X�%����"X�%��{�ͧ"X�%��o�iȂؖPF���V��QHFAn��A%����"X�%��{�ͧ"X�%��o�iȖ%�by���ND��F��ҷD@�$M�e�4�ı=�wٴ�Kı<���m9ı,O>�}��r%�bX�}�xm9(#A���0ji��r�nG$7C�,K���ٴ�Kı<���WiȖ%�by����Kı=�wٴ���oq���C�O�1�(,�]A�r�s�Kn�����h��m7G^��y�8� FG"�E!�4��h}�{�Ȗ%�by����Kı=�wٰ��Cșı=�w�m9ı�Ѿ��+�6��ىȮ�h"�'�}�NB�$D'��q5������r%�bX����6��bX�'�}���9ı,O~>��Y;�I�fKu�Ѵ�Kı=�wٴ�Kı<���m9�ı<���WiȖ%�by����Kı)���왚35e��&kSiȖ%�by����r%�bX�}�����Kı<����r%�bX�����r%�bX���N�%&f�ɩ.e�jm9ı,O>���ӑ,K��=�xm<�bX�'��o��r%�bX�}��6��bX�'����R�#	[�W���.�9p���x��N�ґs���]=9�n#9Z����q��ND�,KϾ��"X�%��{�ͧ"X�%���o�a��L�bX��p]�F�41���Ć6�5�6��bX�'���6���"X����6��bX�'�����Kı<����r%�bX����˓Vfi̹�]kSiȖ%�by����r%�bX�}�y���K �MD�M}�xm9ı,O{��m9ı,N���$)�9��p�F�4��f�ND�,KϾ��"X�%��{�ͧ"X�%���o�iȖ%�bx}��@�q��h��RCt8h#A��3xm9ı,O{��m9ı,O>�}�ND�,KϾ�56��bX�'�?���0n��.2���Sq�WY�-�&���ڹld΀�3��_����E�=���ײ��Y���%�bX������r%�bX�}��6��bX�'�}�jm9ı,O>��6��bX�%<;ܝ�3Ff�.e�5���Kı<���m9ı,O>����r%�bX�}�xm9ı,����t8h#A�C�A�e�-�e̺�M�"X�%���uv��bX�'�}�ND�,K﻾ͧ"X�"4>̽7C��4��0��7QAa�j�5��r%�g� @Ȟ���6��bX�'{��ӑ,K���ٴ�K����~����Ny;�j�4��hk=+<"�l#(��Ȗ%�b}�{ͧ"X�%���o�iȖ%�by�w�]�"X�%�����h᠍h#C�5-ME��Q33�k�s`����%��έʧ�M��Kq�q�Y�s�Љ��m��C��4���/M��bX�'��}��r%�bX�g�w6��DȖ%����ͧ"X�%���_�B�!H�QH�7C��4�����n�D�,K����ӑ,K�����ND�,K���ͧ"AmD������ne�ə�M�$���͉ �'����p� B�������Kı=������Kı=��w	I�j�k%��k6��bX�'�w��r%�bX�w��m9ı,O=����r%�bX�g�w6��bX�%<>�Nə�2i��L�m9ı,O;��6��bX�'���jm9ı,O�߻�ND�,K߻�m9ı,HdȡB2�R$B2ڋ	e�
hF� ���wLi'$�HL�H�	 ����$m�em���'�n��u�պ΍6���Ia�ד�	�j1ӹ�m�c<�C�r7��a]Y׳\��y�0�W2įmϳ��nۃ��]�YD�l�;v�����fwH:�,��at�.�:`q���wn�l�/�rJY���F܆��Q���`��^7mf&3�n�L&�2䄸�Ji�cn�~��9��CB7)xtu��2l��7\�2��gؗ�3Zܵڝ��nԘ�%6����F�4>�o!��Kı>�~�m9ı,O~�xm9ı,O;��6��bX�'O��iM�d0"��n�h#A���ND�,K߻�ND�,K���ͧ"X�%��w��ND�9S"X�3�{� \1%	0�wC��4������"X�%��~�fӑ,ș߻�ڻND�,K��fӑ,K&m3�[R8�4��������Kı=������Kı>�~�m9ı,O~�xm9�h#C+�j	i"H �)��pб,K�u�u�ND�,K����ӑ,K�����ӑ,K��o�i������������.a.���mH=�X6؃N�0���^Õ-���%ó�Ψ�D�9-D�l�$wC��4��}�wC�,K�����ӑ,K��o�iȖ%�by��iȖ%�b{���B��	���Q9�᠍h#C���i�h� ]���D�K��~ͧ"X�%����u�ND�,K����Ӓ�4��>��-�ف�-�t8Rı,O;��6��bX�'���m9ı,O�߻�ND�,K��N�F�4t���aGf�Q�t9ı,O=���m9ı,O�߻�ND�,K߻�ND�,K���ͣ��4��Ʉ����2�7$��r%�bX�g�w6��bX�'�w�6��bX�'��}�ND�,K�u�u�C��4���5��F�2%QH��nl����;�J�c�����l>��L���zd�)�.���R;��A�F�s{�iȖ%�by߷ٴ�Kı<�_wY��Kı>�~�m9ı,OM����i�p]�F�4>����r%�bX�{����r%�bX�g�w6��bX�'�w�6���2����<�^DIC"���E,O~�k6��bX�'���ͧ"X��(aQ�H Da � h�M����ӑ,K����fӒ�4���m���i��M���r%�bX�g�w6��bX�'�w�6��bX�'��}�ND�,K�u�u�Gh#A���(k��1���r%�bX�����r%�bX�w��m9ı,O=���m9ı,O�߻�C��4��fi�̥"q�p��Ӭu�^��5�v^�sۗ��:"��sr�nݙ�V��f��I�Kpr�Ƃ4���o�ӑ,K���}�fӑ,K��=����Kı=����Kı)�`wY�(�l�R2Ct8h#A���7Y��?	��,N����ND�,K����iȖ%�by߷ٴ�Kı�	A�q�d& ܒGt8h#A����ͧ"X�%�����"X�%��~�fӑ,K���}�fӑ,K�dj���(I��#�4��߻�ND�,K���ͧ"X�%����ͧ"X�j�'����ӑ��h|4L�f#$-�dq�t8h�,K���ͧ"X�%������Y��%�bX�ϻ�6��bX�'�w�6�4��h}�t��e�PBY���]m<#Y�tm���c�BdЖ,�=r�5�p�TFE"���F�4>�͏iȖ%�b}����r%�bX�����r%�bX�w��m9ı,O���:�5i�\���F�41�;�ND�,K߻�ND�,K���ͧ"X�%����ͧ"X�%���Zd�jb �TNGt8h#A��w�6��bX�'��}�ND�,K�u�u�ND�,K����ӑ,Kģ�Β��I�K���F�4>߷ٴ�Kı<�_wY��Kı>�~�m9ı,O~��6��bX�%��1���JE�n�h#A{��Y��Kı>�~�m9ı,O���6��bX�'��}�ND�,Kf��Et#�qڢT���0	�R	�$%S0���ĕ)�QR��0�+�9��TӚF�*�m�^>��$�,J�@)7*L1M���4m\ٺ��v��Ro.��\�T�bthI�+H[���HČB05!K"@�"@�@�`� X�lH0 �R�-�K/9�@�{W{�0b LBBUP�*+�4X�aaVD&�lH��d���3�A����!R�{f�u�1��Q�4�T��W����x>�?��N�h'[iWn3�    m     �    p    m�         -�              �p     �         @   UR�m���! ΍أ�1��:�	ܝ��	���qZ.g�y8�'E�qקp\�hҥ�[t�3��e�NS���ȗMt��#�B��`+�����ɼ�1�/[���v9K��֌@��S��"��9ⴜl�k���H�X��m�>[�L�#��xj^��Q�mv���ϳ�kn����n8�Qyܛ�rH�9wd6U;;l�[<�v�C�à���70N�]�(�����p��]�Nv��`�����؛<�#&lvU˧��۱Z���m���!ƅ���E�wm��vE�IA�lr�wa�d;;Vʄ�7V��ݲ�F�$��gP��j�S�i�T��-�q8I��pU[\n\�N<�6C��b��N�&�u�܅�NK��a]��p����k��.��B�6ݻc��X�A::q]�K�{<��z<�w0�a�n�ٞ^�$�c�� \�{3��q�sOK�W.���y1����1ɶ�[�7�[�N�3�]6Cμ��Ѥ��m��l�J7�x��cr�N��Ӷ�>�;02Ɏ�"�n4��$Ɍ��;�[%�7��j^��1��p���2��N�8}��l��<���U�s�v9�<�F�%Nʛ�.s��r�t��ۜ]�U���2e����k�Q����j�֑zzx��u90�;u����ϐv��y̺:���k�T�n3՚B���\�p��&�6x�GeY#���֪9��ݔ�ِ��r.ͦ�ݭ; Y�4]���Ն�f@U.,��k�Z:+ӹ5i��t5�]��nt�Y(۫f��e����v��64nJ:���A�)�u������� m��**z��G �N�`B�@`�|OB9$��$��� 0H��� .��$�[��&	���aj�������Ի�n�q��^D��u��y�:Q�K:����Տc@�rk����;�;C6���i�j�aܑ�A=�1=\�k��l�͍�1T����aR�`ĝ�K����ݸ9�/n7F��;vc�ma��H�ԕ���sq�RH�u!��RR�P  �T,�Jԍ(dJ$����v[���h�!հ9\��v�Uh��۲���2��Ѽ����7�����=�siȖ%�b}�wٴ�Kı<����r%�bX�{��Y��K�hu��4�$�Ԏ�p�E,K﻾ͧ"X�%��~�fӑ,K���w�ͧ"X�%��{�siȔ�F�40h����FHYmH��pб,K���ͧ"X�%���u�ND�,K����ӑ,K����iȄh#A]P+Q�ApȤ7C���bX�{��Y��Kı>�~�m9ı,O���6��bX�'��}�ND#A��f�h�F��4�-��"X�%��{�siȖ%�b}�wٴ�Kı<����r%�bX�{��Y�᠍h#C�
O�ux�"q�(�>�G\^.���c�m�5��z�*��ir��b"�]uś���^����oq����iȖ%�by߷ٴ�Kı<�]�a�	�L�bX�ϻ�6��F�4��Fy��%�-�\��p��bX�w��m9�uQ�U�
�w�,O��w3iȖ%�b{����r%�bX�}��m9ı,J;�֣
1"����F�4<�]�iȖ%�b}����r%�bX�}��m9ı,O;��6��bX�#ra(=r8��#M��wC��4��}����r%�bX�}��m9ı,O;��6��bX�A&D������r!�F�2���\1$0�wC�,K����iȖ%�by߷ٴ�Kı=�]�fӑ,K��=���᠍h#C^j�[q�Zq5�E���$=�����k����\u�S}�u#�kv��1#A�"���A�F�ۗ���Kı=�]�fӑ,K��=����Kı>����r%�bX�>��j0�#*9��p�F�4�����9ı,O�ﻛND�,K﻾ͧ"X�%��{�ͧ"X�%���wq�(�QF����᠍h#Cf�ӑ,K����iȖ?�0"��������iȖ%�b}�~��8h#A����Z��Al���ӑ,K? @ȟ~���iȖ%�b{���M�"X�%������ND�, Y��w��qGFy���)6�SD~����9��v��L�����������V��Χ�&��OM��;v��3�:�����j�[�$�=.�������� :d������,u��$	�܎G�r��ٙT 	��VI�vi�O:���$�1w!P$"Kz��h[)�����]��U����q�l��5���n��� <���\sY_eUU}B�UT�/-Y'��x�X���I!�O:���'@U׹�����VI��0��~�7���Cb�uv֧��ڶ9;j�r)I׍���wh����:J�غ�n6�w3.�3s}& :d����u��tLJ�1�6(��@���t� c����z�a7hl���5!�{�S@�;[�<�k�:�M �S�G�<��16�4�1��bɰ@wc���.�f� L�$����^���h�����Z��7��$�$�L�@ $ � �� 6� MVݶ�x�G5�|f�4�	��8Ĝ�qz9���ZWӷmk��H�ڲ�F��=p=g��ivWB:@��aL�#�.s2���C�T�rlF�pf��u��N'�<ndw�q�c]vz��A��X�������ٺ�f�,��v�����8�b]Uc�a&�gJR�bY�$!�@UW�B���v�n5N&��a�c�����C����=[H�C�V�4!���9 �HD���5#���M�}V��v��|�k�=�em2"H�6��wDv9h�&b��bɰ_�@I����Ƞ�(�n+$�^������`���-�s.����k����^���h��:��u�$�FD�K[���a�܎�.M����1��1�H+�B�q	n;=\u��v�{8۵73�������\曎Ml��
rV��r��L�����*@У�j0�� M��{��n�@m m`1`@	���vv@M#qh#F# ��@���!�F,1���M� �H1�F"s B! �b�� �F0�C�&(BjF)!$b��E�__QG_��@~�"�v9hx��&n��!�ӒHݒx��vI�fX�����^j�/?ߛ��[B&�"`ԏ@}"�v9hy&b��b�V86�S�QL�=��h�kz�ֽ�n�W��MH�B�D�X�*���)�I��6���Fv9ck:�y�]S6�,D�d�C#qh�kz޲�z���}V��z6�*8ءk��@{�T�}"�v9hy&b�:'�U�������n��>��S��ba�!A �_}UO������t���Y7j�'�mbnf�����/�Z����n��[���ak#ġ2cQŠ7�n =�*@wH�ݎZ��,��"��m7���]�\�\����D��6\��\��2M�g+Qls4ƭ�M(t���*@wc��������a&O��/�~��a!o0#��{��m�ٙ�������G�}�2��~�Ȣ�D�ɚ����;�X������b�=��$���X��
�F�㛈t���*@���W�Q���g���mZ��mbTq��4��t���*@wc��o�@K �?�rE�]c�����{����B&�˹���\���_Z��-ΎL�;^�ߕ ;��@6�m�=�*@uײ���d�M�M��=��h�,Z�EH� 
�Q%f�e鹅m^f����m�R�EH�r�y�,u��$"?��H��n��[��}��hϬz˰���B&�#h76��*@{��@7�n =�*�I��~�_�ݒ��p�[@ @6�ݶm�  ��I��I8�N�a�Ehs��;cI�Ygyr�2�Ymf��s19�\Z��;����<�aN.]�@�t�r�Os��[��[�;�ӑNK�C]��6�88�Qq�]rp^)5��ZF���'ne��m��9���/m��I�.{sͯ�ɻ=m�K!�l�9XI��;=9{���A	F4$rt1��N9��ckƢz�<�ܪqۭy������L�4u͈z"��43v�3��@7�n =�*@wH����V
�E2`���;�X���b�?}�b�<������	lQ���f� 9�ʐ�*@{��@7�c�;��<�DȘ�qG3@���@{��@7�n =�*@u�T�f��&�&�hy�Zs�=�u��;��h�n�%"q��IF�1�[^���8���8�s�F{\���jw]�s<�HѓrE�w;c�>�]��n���U�}����㌐��nI#�>�߶n��@b�H*�+[IE��
�-Kh�"!B�U؈�W�|����㖀��@z�K���M�D��f���M�>�@���@��w4�s��yP��9 ��c����@{�T��{��*�TH�L �Z��z�����]��OۓM�y��+$�U
�D:J�l�K�fwm�-rq�Y6��V�WF[{
c7l�ԍ��:8�X�횟����������r�c�����qA(�j)!�}zS@�Ϫ�-}c�O>��zIC�Q�\�Fe&�ot@s���c��ߺ��ꢨ����!�P�Lx�ǁ�
h&
qB�X�bh<����5����%3a)�3III� �-
�(4 y�0���L�  lP�x����OC��'���|
p�` yp1Q׺�5�ܓ�{����0�x�HѓrE�Z�Ǡ}��>�)�}��h�Ac��!��wwq�{�� =��$�7������!jƄ���z�ɝ�N2�pU����nq��n� .�Սq��."-�B�Y�� =���-&9���9M �\�(�E"f)�Hhy�Z������� �Y.�%n܀(A��_X���s@���@�Ϫ�.{�k�G�E�@��{���=��ﾕ��}XM�q ��'��r<J$��HhW�h�3�/���;�=�t���qu�H�Cj;nmw��v��������˞�����%��vzc�n��+�2cD�I�d�M���=��Z��z��M��� �R���	9"�NgfE~�G���d���!��U�{���d�G�q������ZݎZG�[�3wwȓ��I����>�@���@��)�˝EȢ�o�LnE�{��@I"��{�Ih��U}�hk$(҄ UV$'��W�,� �� �`��%� �8����v��������!ЖUlj�r���k�:�gSa��,��5��}�ݶ z󣋭�7����v�v#O[R<F�cam���<�T����X��W��"�k���lJ[��ֽ������]�D祧Y[�h�q�' n�3����;��S��e�	��H���+h
�"��?D�F�grg\����C�-n��Ǳ�a����gG3ř�T淮��Mm�Yk�{���@{�T���-��-+�mbV(�ȲH`�f����hWj�>����4�tObrLJ$����@zd���c��rE����{*.�����I����U�u�Y�}��>�ՠ�Q\��d�37v�H�@{���Zݎ_�o����$\:0ݶ�<�۴��;W=�}�H�w\��zfc�fu�9��'�va�O1�+$���^��\A~���<����I0��	��4�Ͼ��$@�$#H�`6U}_|��y���,�/�UWas�_�BG��ԋ@�;�hm�h{���v�����J�#�[��ڡTn��O�ͱd�c�VI�Ϫ�.{�ky#�"�!����봀��-��- ��;����e����u��z�v;H:+����5��s�le��b-U�R�0�� �7}��ZݎZ��ﾯXs�� ��GA�A��I��y��+�G7vٲO�ͱd�c�W����ӥh�$���nH����l�'�w,Y�@@��B�T��d�����?u�)�j8ˑN$�6N��(�sx,����d�|����*����6I��I��(6�7D�Ihv9h$X =�a�N�ͽE���P@J�	�]�!4�ݣ���͘�8붩@�c��A�V!�5�>���u�Y�}�����$�t=@�
G !CqY'��lފ�?w6Œ~ݚl�ϟqY'�6�7H�Ƞ��f����h[)�}��hm�h��	�㘒�����@zM�ݎZɳ-z�����!!"�H�I ,$�X����י���{OQp�&FO��M�hy�Z[+Z�빠}l����jq4�"Q5ĕ�6�W:���ݱ<��Q^܉�|s��%���z���H��@��ܑhl�h{������}V��t+JF(L����Z���� =���`��geVH���	����e4�������u���է���k74@{��@9"��qR�UUK���d����%��$�n+$�fb���� =��=nJ32�p	 p� 0H��� 6�UU��rG'+�����D�VX�Ku�{v��<�k��XyÉ�Kk�.�7nƹ0g��[�u�=7kP�gU�;K�5M�M�q�Su�Uխ����[�D�B�j���g0nVs�AE�[\�;�.�Ck���`{ju7R��@"%�A�;p!�Z���f:�6�K���i�c���}���%��2��j�k�r9'(k���:�[��rnuɢ#��,P1̩��sE�vY��~T������&b�8�'S�bJ&����>�S@�Ϫ�:�[�>�]��=��dd�6�f��c��rE����� �(� ,�F6�@�ҵ�}�`��c���Y�n�{�}y���hs���`��c��q���m�����VK#	v��p��4�<9P㋝՚�]�2[H�%�M�WB4����j*F�����HG�@{��@8�e�}_W�A4�e�ӊd�Aǁ1��3߮�m�Vk�os��˹�]��Қ{X+�)#G�{2�n*Gﾯ������Oր�J�<PƟ�k@���hW�hs��+Z{:6	��%]�nm =1�@y㖀s�@y��@�֚�MF̑5�&@�L& �.��!��Nk�]����)#��G&˜�qɮ��I1��@��U�u�Z�>���ÿ?� ˔��
!�21�$Z�ހ����?ր��-β�L#���N)#z��s@���N���̀ �"� �Ȭ��*=����9V�|�o@�gT�Q�XF^m =1�@y㖀q��A�����Y$�FkN($j�Y'�>�:���w]������MH�1Tsz��p����źC��Ҧ��˞��u�6��h�=��k��Sr\�I?_����s����=��%s�˫���pq9�I�>�]�����>�@�ҵ�w��`�R9�Q���f��ZݎZ?}Uw?M����?*@;����y22bi���>�@�ҵ���߶nC�K,�Ł�<���@2�??آI#rE�u{2�n*@zc����-%c�]�1#lm7��λbPz೷]uZ9��-5'mr�	�\�r�qls:lZ�i>����9h<r�z�~��-�S���(��bi��>���>��hzV����z�V�S#j?�csm�Zǳ-���9h��V
��J'�N-�Jց�u��O1���@�L�d���	kQ�����ܴ�����<��@8�eܓ��d�I�@���vF.�l16B��d�HI#HɄ��ჴ>W�D E��9���V"�ekF�]��T=#T�#	D�� I	T��G�B$��5C	Y�V%"BWI�#$&�0��� ����4FA��w�e�j�UֵR(9�6�l�@     �           �    p     [Am          �   �     �     ,0    �    	'[,��F�jݸ9!Ӭ*�n��ܙyfy�:н(�������ŝ������<�vG�݌�Z⪪���PnM�z	�-��«Q͉v�/n�����ul�rW��)�ǉ���V�Vkcla�S��^7YZf���K�䗬L��م�/%8x��֪Ԡ�Om�Y����W2I�{m�\���ݶ�3t� �� ��y��<�e:�ٙ�%��X�
�̳��1k�d\Z�l�G�"ꌝV'K�6��sgr��u�vm9X�m�w"c@[fX��؉[�;Y����n��I<�pn��N�R�ˉӌe�<����Z@촦�%u�n�%�Z���'���[FʁQ\˱i�w�jᬇ5ml�H.�ɳ��p�L���|=���r���󬃉��9vu��y;DBU���Lԫ�a�mϓq�V�.�n66��`�O3͹6؋I��.tbd�%�8�@�Z�H�@Y,����,kN��n(�j�/6��팒֙|�W+dN��C��k�XQ��1sqc`CV�i��Ё�MImlAnJ;YX����D!�tm۵FV筹9�����Tp���z6�93�z�c+ڷ��H�U�rz��t�%݅i�L�f,1�`��pc��E*�R;��8���REn�yA�u[c-Ԭlbď =R+����v���(f݂�漳jh�n�/T�s#���%Ζ�y��ū�`7m���!�K��\Pmss�n��%��@��F���������-�cm�Π�V���Zj;$ti�[��d��"q�,U�m[m=)am[pm�u����\��Ō�j���+�]�&FmH�jB��P�
���_A��6�	��D��R!�ꮹ��h��kZִkZ֎�� 	 ��� � q�k�/]�n7c�΃�u��Lh�m@��]և��4a��^����sS�C�c�`CK�-0�[\���z�j��Nz�Hw1��p웯����v�;lrK��ub/v����I��Ù,`G��݆�읚�ڋc$�ڞ.ZwS=�Μ�F��m�cRY�ʎ�v�V���O�Ĉ�5!-�L�4�͸�t�uF�Oc��$3�9w��lX.z�}�\/8��9�Q���g�:��hs��+Z�빠r�eE�<�jbi�-��- �ٖ��8��Z ��+��I��1�$Z^���u��>���>��v:	��AI����ܴ��HLr��r�=�h�uJ�DFD0&s4������Jց���hqԪj(�B"Hq�gu����ۇ�ה�O�S�N8-v�2u�B7	��h����,��r��������kzX���s@���@��:�VI"�<��h��j��ď��s@���By��+�UPH��F�KZ��.d����HLr��r�=�h��ǉ��%JH�h׬�>��'�ٍY;T(�sx,��tf���@���3swu��- �ٖ��8� zu�v[�IH�Cj'0J&���^�VC����Od(Mx�n%뇭�	���k���Fz�~�33wm �ٖ��8� z9�s�v:	��AI���r5�}��4����J����ď~y�%�(�FFc&s4߯�}��i��d�H�=т�ACEa�H�H���|�7��˹'�{��@=s�R)����C�hy�Z�fZ���9�]Y.��e�����i{��q��@{�T���1�}V���PUGML�4�
�8x�x�I�8�p�<x�l�ԍ����
�(���$�h{���^���U�u�Z��sx���%JH�h�� =��{2�� �S�,#ɊDcmI#�>���+Z�빠|�W��⻊!�?�rE�9�f =�*@z㘁S��������� | B�y������S8̐�1�RF���s@������-����'kte�����(��%2����d;)�m0�<0�nq��ۂ�ںH�'�P�
(�FFc&s>���������ށ���h�r�D�6��0�����- �9���8��b�VU�\��Ey"�:���{�柳��=���\�F�%A�H�S��w1�qR������b �g7��9�Q���f��^���U�u}[�>�]� �;�X��I0@$� �`��%��� �I]����M�NjI�od���@�ۣr�`F+ظ,l��/�Y%����3�>v%;����`x۷Ͷa%�fL��g�nhpҹ�Gmݮ���{F�t����r��i&��80��ۯ%�t�u�AN�Ol��Q�M j�2�%��a�nWT�� �eЗhpW�ۯw�jpP�Ro6���:ݯ�z�c�A�.��z�EѶkWr:T�ӦeC9Α��b��RH�W�����zϻ�?UP�"~[��GFzE���fn��3� =nL@{���>��ed����I�>�]��ֽ�>�@�v��}^T��<Q��ɀ���ֽ�>�@�v��� ���sx,�{���P�N;!��-�$�@{�T���1���F�;	=�M���>'{\��{և'��t�5�\��n�N�*H9�Q�2L��EH[���%G��KP��jREd�}�bؠ+�uB�����@s�-ҲK@��VT�䄣JH�OWs�~�����IwC�VI���,���P1���ڋw��:VIht��ܘ�+�ӏ�� �i��~���tUW�����_ߞ��>�@��*�M(H�.�����H�;@̻��cg������;v^���gOC�u]Q������T�v��v9h��Z�*]���ĦFc&s4]k�=��h��Z޷s@>�UR'�����;��@t���]_U*����� >]k�;=����D��E"�=q�ht���L@wc����]]�d�G���@���h��ߟ�w;�h��� ������7���2�����;6���dn.snt׫��srd��٘�Q��I�JH�h�k�=��h���@���'��زO�`�e�H������v9h��Z�"���4=�WqD<�'�cNH�\}V��R�I��r�����&����$b8�� UP���Y'w]�~���� ��X��y�1%�6
�2�36��L@wc���X�=�*@v���z�n5N&���\m�S0��!"�fl���sf�qΜ]���Nw��!����-�U�}�w4^����V%rb�Hُ�)�돥�=�*@;�1ݎZT{�uwS�w7/~���@{�T�w�b���>�@/��ǎ�$����f���b��J�-�R�N����&)��)��>�@���hz����zٿٝ�.��9$�$�Xa�[A��� lK( �`p��>���(�>�>v��Qɕ�8m�z�]ע\=Ԙݺ�[��'��n{4�-Ց��ql�nͧm��'c=�s��I�#T.�6�'c��)n�C�n��+�V�1��+��n��V�7sv�t;��Sc]{r�`Iw\�s'����,�>���V#���,����t��/3��%**� hH
�fY��iC"Q5i	ю�6�p^؎Zځ�k���ʯ&4��=I�
�� �i�I;�{��<�EH}& ;��@z:���nV�Q�[�[�h�*@;�1�Z�c�~@$~CI݉�T2�	'�qw��@zc���X�8� t�r�r��A��8���\}V��빠r��@�\ubV�8?���@��r��T�w�b������1�/kV����9'9�fZxY.m�ة�F�E�:�ډ�4�����K�-~���:�� =|�@��h�<a��G
)���$�}���g�9����/�]�u*~��ܭ�&!6E#�<�_�@���h/Z�>�aO$���I#�=s�� �����1u��'�XH�8��]���z��z�>�@�T6�Pi���"(�����T:L״�Ձ���3`�g���7r�I�Ɍdē��r��@�^�@���h�WHE��N=��J�- ��H}& :�d�ɎD�f/�H�\}V��빥�̛����.�b1b�XX1���RJ��q�&�`X�Xq@�X�>�	��H�	1!"B� E��r��)+b�@��!�#�D���^1(D�eZ	u���6H$H�Hf���y0�p0�,d7*C��A2��jh����y�g���! �P40�$Y		14\"X�%!1V�F�)�,LA6B!��b	! ��s7�1b�X)D� 1b "a�	��0b��H��X�a@#��u11]`�Ņ���#�$�h8D!��&��|	@����C��~_ i����S�Si�  �����*�^�r�Mˊ"E$k'� �����-ұ�@�6�0b�Y$��r�^��}V��U�w��h֚�MF̑cQLOQ�]u��]˵��CA+�]��/;����	��.sL�Ǆy1I�M�8�����Z�㘀+�Ún]�n�Vᗛ�h+�� �1�Zݎ��qǑ@�,R{���������Z��7��ɉ'3@�mz��Z\v��2��]<@�S��}��nH}�9~qd�PJ?�#�>���:�h+k�?fe��~ME�H�co��u�y�YT�;y�PY�'���T�s�Gb�az�����������]����ϐ{󿖁�:��,��"E?�n-��s@�mz��Z\v� ���;$��1d�f��I�Lr�VIh�*@z�`��&)1	�I��}V���@�u��9[^�g��#I�1�$���Z�䘀��-��{�ߟ���}y��m @	  �l m��I����n�v��I�$�÷4�9�>6�<f��7k�=v�q��:m#�a���ֺ���{n����Ta�[L9�d����d��͵�Z���vp1B[��":�n4\�Y���f�����jvt͵��#����� �`6�t�d��J�:0�W�z3�fҍ["�%6�+A�Gow{��Q��"�m���Z{k�%�%ݺ뚓�ᖚ��lY�g�Y��uI{;7*D�"��'36Œz�1�'����@Uqc��h�?�x)���s4VL@zc��r�K@>qR �D��YD�0���hW�h�hm�@�\yV
�q70�R-J�- ��HI5�Z�=̻\�)�1���]� �٠}_U�[�ՠ_5F�N$d����.Yƞ�wΛw7N#���%P�$����s�k���%�I2< �I&|����@���Bs�^��Nw6Œ~C0�,D�.@��ֳZ���=��<Т�������Y=h�T�$�Pz�sM˼�ݠ�i��n;V��빧���H����{󿖁�r5�܉�P!��#�@�u��m���Z��Z��7��ɉ'3@-�hW�h�h�%SQF�J&��?�!�z7/Wdϵ䞇�B�)Ō���;rצ�nf+����A�a1E$�>���-�j�;�w4�f�����r ���hVIh�*@I�Lr�����q�E����@�u��m�{��ϽU_}�R]3��V9hs��3&�x��I&h������v��
;��d���:�H
�"ےI��$����T�$�P���
�Cp�۳kv|q�`w �Og��;�h��e��9��י�U�NF�@IY%�8� I&�=1�@t���b(L ȄqY'�w,^�D�������qڴ��bo 1�Ww�HI5�bJ�- ��H��<s	�����z�Ͼ��{�lܟH8
�Qy�{��<�l%��$*2Gd���� 	$��9�:��ܗ0�\��;��<v.��1�#-�x�Vس��tmp���
�;�,������ 	��9�	+�9�`�Ŋ
1d�f�[�h+�����]��;�ǑI��ےI�\sV9h��	�^��4���I����: �D�VIλ�h�f��^�뎬n���(�E�E�w�U�����z��ߤ����������p8�-� � ln�    <I�n��ޚ�qm �<r�l{n�c����.���拡e26�5;�']����-�\ח=���Ж§��&�lv�)y빶r87Hq�>�`*�q� D�	�H��AE�{3!�[4����G����I��C��[�7��cv\"����n�NyL[�gN�ۂ�	�=ft�����}�5>)PBD��9�Dv/#���ή9A�p=�s��\,��v^�C��b�s�6����P�� $�r���@�uq�H5&(����z������ ���=�%rc���7wV9h��	��9�G݉�S8p�ܤ���UR���d߯�|�W�[����m�1��((őH�޳@�^�@�U�w�U�}�e�8��s��f)���W�Ge����{n�Χ��=���Ϸ1��Nz��LCnI$�/���-Δ�;Ϫ�z� Ͽ�\�'�2&5$�@�:S{1@�x< ������O<��n��z�:�����X�4�r��j����<�5&
��Y�(�}@U�se�~[��s���}V�}p���A��LQI,�ŝ�d�n��s�5Y$�v��%Cj8ƜML��,l����xv؝�0�ؗ���˻�H!�wn���Nj;p��Nb�$z�n��Қm�@�[^��,�b����L�;�Q I&�=rL@IR*@�faE\ւ�FPq�d���,�ř��
ʡU ��(�"�P7�h��7$��)�}^Z6�G�8��$�@�[]�se�$���l���[���$}][���FɈi�$z�e4��m����z%[��	���%8n�9���!9G�q��k�"cg���3�n�;v�25�̘�`��!�wt��[l�>Vנ[�S@��PV$�R1
C@-�h+k�-�)�wt��z��ǎa ��&(�����r�h�)��4ˎ��1���_���J�o`�$�P%�}O�`�!%\��`�!H��TC�a (L�X�A�,b5�B)��� 
�Q 
��9g]�x3���!j������Қm�@�[^�nYM ������7��̐q�1/����^��ᑻ\���M�F��x{v�mTj�wn)1AF,q�@-�h+k�-�)�wt���yr�#y�ےI4��ޤwF�6I�ɦ�'32^�H��uh֓�15$�@��?OƁ�Қm�@�[^�뎬n�C��X�4��f^�$���d�,�vNСUT�N��@�y���Hd�) �٤��(}7u�IѯL$��Ӧ�> *��Ѐ"���@U���"�D_�PU�@U�Ȁ"��� �����"� �"� *�"����"*�"����@@�"����"�@�"��",R(��"",��$`��V(�",�,Q",P ��B(�"(����"����_�Uh�"�D^
 ����*�� ����"��� ����*��"��"����
�2�ɣ�P �������9�>�r|�@$� � (� 
���E $P�@ W  z�B�      ����I�
%DH%(�!B�QAJ@P����$�)B��� K�  5EJ ( B�� ��&[�n����q7Mŕ>� �[�{�O&�n39��9��F�{\�r��� ����qn�w� w�i�{�*Sܰ�9��Z.Z���
{�=N��q l�;k����� Ǆ �� �T
&6@ޥX�|A�n4����W�}� �-��,\�\��[�85�� �I��ۮ��Ӏ �r�� >����Vv��'��e��F�ʻ�@�zk��y���3s�����ԾϨ�    )�`��kk��e9={7�gJ��ڛ�@G��cs��I�k�zyx^�6���x {�>������}�e�r����@;ϥ����t�n�����m��H y�����:ynz�x���R� ��P(  ( ��4�Ծ�3���x�)@� h��
3�����@�� b�q�` "t4c  Ҙ�h�� 0��LM
bh�)gs� .3J
[� ��14PM(��hS@( 㨀* N���1@҂�3J
1��6PQ���E�p��T���8���>�>�n@�K�S�/� q�{���+� ����Ů��ݵ���yn��Q�znm����ׯv�n����ï zBM���=LA�?�SoUR� `@ ���R��=OSL�4=��I�IP  "��J�ڥ)P   ���l�*�� ��P���/��W��������3+1FJ�JB��C2��"��� ����*����*��DU`� �����o�>k��!�	K�s�q	M!8�'@�d�R��"h0ap �͕�`D�@�8l��VBHH4�a7�Fn�H�54`����M@������b?��BR�Q4L��]jm�%s)!�v��}��믩�ލ��aA�h���bD�6SZ�@�#tS%	���
1�q�C���7���\�9�;�eu���!���(c)�4�+ �,JJ�1 �^|N&�{���4�?��h&Î!����f��vF��7�'j~����d�K�pe�I�9��?���u��|:�?��tŢqQ|_e|��W�ƑmM�`�D%0����C��q"�`�w��W�~Ja�t�9�$� ��P�#	�!���h���I�A���c��?0�?0&~4)��\6�H�@����R�JNL�Z��!�j�G���BD��>�3��t��~q�щcH��U�4E�1�)�ȅVfs�O�k߷�F���䡿���-��>�p(@�ˀC�!�JS�d@�MK�8�_p:�����$[����������$�P �M0���+� ���WF��0��
�u��?��+�6�1�a$n�fp�i�%4�L�p`t8�����tQ`i`��WR)�44F��DSoJ�l \����� F-d`�:���}��`QdȐ��@,��܌&��|�Ȍb'��t��rNd �#��GM�F�͟���L���$��	�qzO���"��U��ీ����Jes��a
��#u
BC~��5�t>�2�B�$bh �4���0k
�$(ĠhX�d	�'�����[���d�D������d!L�p���
��B������Nk���a$�H��HI%4
h>��~?�i� �8����o	�w�hH4g�,
�2o����Z	�f���D����)Y��ʹ��2�?k98|��������O���§L�cP��{.���5��_��G�?�]k>�2�o��5M[���F HH0@�)�Z�$tƐ��_��F���PLD��,]�H"P_M$�W�T+���qp;#HT"@$M��6BXX��"T�FD�$J0�	X���~2Q�"�_���M�?k���.�]fӅ�Ji!X_�$`@��,1�WN@$�K�4�h4h%�|�(J~?4�w����l�l��6��5i�5��V�5�a#��
�i��D�u(�a�##�����%ѕ��8M
����*.u?G~ہn��)����ڔ��tC�t\]�9�er��	 ��9!�~H�%�H\��
Ť�i�g?r��6Fs�n��Ԗd�,�)��
�����+�#Z�o��<?')��g8�����D�#D�tj�����C|8~X�!u�?|`߱	�����H�6?M�����"SA�ÌB�/TQ��@�BH�tj,@��сOݍB]�¤��JB�D`M:�	4RLE�PC*T����R�8���d� @��H�`�HT�j��H]],(B,+� �*�(@%5#�Ѣ�HY�"Ȅ�V�[44���A�R�
�i�ZV��R�WEV��ԅ�$�9�4�n��A�)�VXI��� q�6jӣ��X�]c��%�_�p�wL�@�d^����ۺ�ԍ4º���HQ�����k`�m��
��g?O�8�C��� �����5�S�!���o'�FL.��Ny5Ąԉ�Dv�>�R%���&��}?$*J�ѤO߂A�")+EҎ�ʡu���]��S���Y�:%>~+��X�"�"�ĉ ��/�D�����Á�>~H�O��i	�__��'��P|�Ŋ?:j�����T$! �&L�q(C+
F�&k|�4f�ji���f��].`U�@�x�X��4џ?~��d�0��s񳟏��`&��NR���]�ӟ����JC�ݯ)����Wf]j�j$MA1  HHW0'ND'2��J�	˔J�ܜ�J�ڕ�/���g����c9	+�m*H_�XĆ�	aWI.�o��2	 M!4���,�ς���vU�ME�T����ҔHZr�	���!SB�H��A�H^��NsN��F� �"�1²A�In�CP$!���b� D�W�ʫM)��'NR�IU�!�~z�/܅H�a�=4I�b�XĲJ���k�|`m�H:`X���Y��8�D�$�1�B@� !�����F"ؐFB$�`; v�6H�`�:�0cCN;�l�F5�6�(iKa��A@�f�]l������gN?$
k��?%ѣ��i?#��[�Iu����B0�V �t�d�SXm�u��.Ï� ��`W@~a�	���'ٚ�9Ns��.r�_�&��!�L��+>�e�]�o�U��J�� �N��	1HN����4��1�����a����-s�)�M"R!�2rc�GWs���|�,�qd	��^}��~�K;+�Ѯ~�k���X��3��Ǫu�A�_��$X0s��s����fn��ܖ���W���A���v���1}�|��SJ���M,���C�Hk�V�D�HEÁ�ц��S�i�?SI�g��N�����8��>�,�d�Yp��R[����Cw���5��d`��s��SM�s�A$��v���K��NU����R����~0��ᧈ�:I$"I#`�[�|	�e-���d4|�@�H���	a�Hm7&�!�6p8|���|?��]8l�������4c��~�|}#�4m���~�5���>X��~�]?�!MT�I	aߎFMr�;�v2�즜HXSL���,$$��
Ma�p���C���>Jh ��I#]#���ğrGo	SQH,.�p�oS���lm޳z�ϕ%_U��\GGw�J��9��"�X$#@�ffr�޹�9�k���5���|�"C�@#�c
���>�>�C�Lv���q��|�(h�|�|�,)��g����b];x~?}��5�a��� |*��o?Ѩ�t���2H�$! F��"�����1���4oSZ4�@r��I#BWl]6X�X�?	��"���,b�B��4$� BȬ�+HSF�4���5��@�k
i�d�t��6� P�����$��M8ƴ�L Q�\����ј����M�`AH���N�����ӄ�~�l6�����ՄX�F�a�n��?HȄh�ɳ�Ӥ� � ��X;KRW�|CG�:y���㱌#�|��i��}{x�%4F�a�yL�$i�7�t�ǿ�5�?lp#�����Dr�_1}��b��]|��J��L����-Jj�\_H��K�(�J:��ur{��   ��                          6��#}��                                 mp�` �llإ����ඍ��	k� �E	���@,1l�R�{$���Mi��`��`m���CSamI��J�Zj��;tUS�յ[Uʲ������2�o[�`�n� ����m�       h m  :�i -��;�����kw/l��5�R�a1�vX�F�Tt�5*�]6��mNU����U��l kX �nm[l � n������ �-���   ��0�n�j��oP�I�  �� -�h�mT�j��B�@      M��m�m�5� m   �vm�ݶ H   
U���-UR��Ғ�;`�]. ͮ K(���v 4P                             �Jٲ�           ��  �rD�                                                         �|                                         �                                                           |8 �m�-��  ��                                                     ��    l�j�M� �+m�n�� R����-ҵM��i�l�ۀ$ lv�V�m�I,��h�o�I��(�R�lL�� ��Ԥ�ҨUT�� �Ͷ#m�@X��6�t-� �ն�����k�À h��sn�h,��E趀 ��l��$�d�m�h��l �`�(k4�M�Um�M���UR�*���:�� ��� ���l�K��ʷT�Y{a�Pk�e��  �6�eR�&�ԄEvq�t�}��}�d�m�Zl�gm� � �l��Y3���k�W-��@$JKP
��m ����մHM�I��I�z�F�L��e�� M�      � $�H�:�v��׋s��r�ʫ�ͬ
WjjB@���*�UUUJ�P   #�
�v�_9E	
@P�36�M��� �:��N�l   *^y�E������UF��lӮ�e���E�-붳H�%�h�w� ـ[�2�Uj�K\�(VU88�;	��N.�kN�Scvu�k/)��ګ{ $6��-bBm&I�mn�ݷn�tV���m�6ٶ�  6��$@n�p���`l�XĖH�-�uu�J�l�@Pn��5Ӱ�`z�8�b����n���h-���M�m�sAA���Ŵ 6��Cj�m6�� 8�r��ֻi0[\m[p �t� v�l �	���Z,�h  l���p�u� M�E�� �m �MCl�FZ��6�g[�� Q�@���l� Sʁ�eͶƊ ���!t�mji3]06�Q#m������6C�pp�I���l�;}�
�� 0u-+p�m�U��ZSk�^�l -��5���iT��l�uU��\���� p�oQ��zۀ���\6d���Y�{6��H5� ��nٶ�L����9kelL�*��T ��G��a�䁙��+ec^�j�ŶӸ��ktS���v��5+�0Yۊ�̭b)5a�,�UUAƃj���3��Y$�ڨ	P㝥�4�m�m����gM���6��Gf0��PYzM�k,���[A�R^�2�		;e�H lv۵% X�նRIkbt�: �*�&(�R�V�U@A��j�]���B*��6�c��q/@��(ҭR��������V˽���FP�g��@T�쫧�j�	��V{ܶ�T��F��p��+���G�u���% �i'{�a	X�4+�K�3�����V���
C������=��[4��[@��.�m� rlXkh�`�Y��)B��V����*�Ͼ��&`:A� �cl�tȷ+L�X��ҭPmR���f�3m�t�K���'Y�Hm�p��e������u8�� ��Z��I��Z�-mT��mK�UR�ڭX@AB�s�T����F�VU�+[�� �����8܁FEz��uV�l]*����;�������uWk��죜����7S&�s�vl�@�v9r�5u��湨���9pb�l���1e�"Dk�v�#���1��歬�  m�Z�ndm����"�m�Hpp�� �`'H3k*�
�u)-]UU*�  vԢ�6�I�h�'S�jA��{nsm��l�� ��Þm� K(	�[uVʻT��.p5�X�۲CF�m�!^P+Wb�٧�5Tݲ�*�UU*ʀ�J�*�*�T�P[U��J��x �m:l89�m�%�M�6�A���6� ��β����i0[*tXiH ��8���e�m�jvͶ06�kI6հy��m���*���`(0S�� &;l���
�U*�UUmUU�� Isм��/.m�l�Wi�κ�Z�T���:�:�h2�UEq�g��gN���V\������`���&�!0I��M�lU�aVU/���kn�[�C[??}���6�b8�),gw@ş]v��P�1�v�"x��";=�I�����=W �5u�=+ř��K�c����|����]d�l��ʑs�ӕY㪣���p�ny`�㱺�a�U�k��;M�������ݶ���k�.�v�N6�vVH��gl�Gc�VW�[l��Av�	/ZM.�CKy$Zk� jض�pp��6�䁴�F�[�H�t� �8  6�m��r���m=bK��@d���ϛ}�� Ą�mq�˪�z{e�v�n��[T %i��mvƵ� H �� :@Y-9Ͷ�Ҷic�6��ڶqm m� 	�vum��0�>�E��m�m���l�@��p u�u� �`@���w.��/��m�}d�	8 �l�    
��WfV�6GmR�l�u���`h��9�   l �7gi���n��7�]��e^ Ku���%-���)�ll �غU��]��Ƥvһm�n�7$�����Hm%��n��E� lI,��+�v"�v@6k��jLbjԳl�� ��"�����-H�<�.�u̪�0����M�ӵ���y�m����y��ݩU��avt����-� V����$�cf��`��ztm��d��Y��m�����7�:�HZ�F|=Ut9���Uʜ� ��/[�-�o����>8����ն�m&g�}������mJ��\��(�R�h *��T�U �4���6Z�j�I�t�I�zIIgW  ��m�ehjI��p5W[e�<�m���rN�[�!!y;m�|�zIwH	��MN�m�F��-�6��t&��m��I� #�]n ZѢ[d6� �kj�TjCb�
X�mR�!r�����H ��Ddm�6�{Mw8��`T����f�8]����n� 7mi6��Ygv��    6͵�$kX jB�m�n�d��MT�Um�iV���UU$ p=&��	ХHs��Ӧװ�l H�   �km� �D�l�����8I&�@h����)U��U�b��@7mj�Cn� �6��fIbR۫�] ��5�<v�j��퓳����O2��36��:��Q�YV�I�b���� �v�]�Mmxmk]�q���`�rD�ݰ 86��d��4�ۖ��;V�H�dm̕���m��    � :��j� �UUPW)�9P:1�(|�� �t�ũ�m������Ơ6j�m�e,�ڦ�	-Um+Q�}�eM]^ٻl �TcUW)*���&*�+�yZ���cQ�t���p�m�K�R`-�M�yg[rNk		��ll8   ��   �| �"Gkn���	  �ݰ4V�m&�:*�%�6��*�v�]���T�V�r� $�',0����ww{������� N(?�- ��G�
�A���UO�
�J�4����¨�������@pS�B(�C�Z"� ���a F!�"FbIIE ?+�W�|"@��>:��PN
@ �~!j�P�EA8.��""���Q5�@��'Db`�X*j�qZ��? ����(�����D_�:T�
LA䢈< 4 l� �ӊ���i?��Uϐ��1�@$$	$��,H@���� 28'N�"�+lEJE(�P��	��8��W_1H�B(B0$�D�`$1!?(3�H��� X��IC�Dd�H�$XH�UJ*-J���
�B�EGhAHB�$�+̀���'Ep�B*;�`=V+�Av�*�P�DC������ 4@�"�=Pb�|��S�k���v"�*@U�P"U� �]� ���*�Q�"�B(� `*��
7���0    �`      ���۱Od��s�V͎�]�{=:���&� S�<b��u�mZ��v��5KsW2�\��Ί�UV����(�6�V��u.�     �  m��I0        6�  l             �     k�Y�      �   6�9�ml.��^�^6��K�V�i�S�H7/:�Jq�u�I�!�Gl�g9jC��r��[���K������7;T�tӤ뭶n٬��a�-� �Ղ�͞��n���9��:6���-��\���dE�^E��tY K����Yv5.6ɞ��A@3;*���.��4*d�::^�1'��5Hs�,�9#�]�49���cjm��»1E]ڑ�=�Ш�C�조Pe�kI��v�p`�Svh�Sm��[b�[Ҩv��+<t��[Jt�5eu��/3�-�2���]v��(!�6�ڭAl]�:��F͸mq�(y⇜J�j�[�!�	`�q[mvG���p
�w%ڷL<y�M�l��o�9��\�'5�*KgHv1�"c�բ�U]�	v�ΰ��F�5�z��S<�/m��\�@��t�'c`z<�H���p�u��1�݈8���< ��"����e@����:7R���8�'��6�GS-�K-۲m�i�h��-���6��뇂�1��gj{EUt�:Þ�"ZB�0o�1�II��2��9��'�&8Ή�=i�r��5(��A�ct�8���ۡj��ƢnS��++ƚ�V��]��Ɗݻ>�L�V��Xh�:��FX�	�89�v괥ʬ-���Kz[��-�z/9��ザgF�]t���^�J�����P��d���<�)Te��g#�<��[:�7U��f���N�Z��!�����.��0���f��k5�_���]
�mv�QW�A~C�D���G��pW��Wh�E��33-����V)5���v��S���� � 6ٶ�	 8m�6�ފ��^iZ�A�=�g.�!�[�7�1͋4;�\f�܌�pEV볒�.��z����k���vM��ϧJ�ʝn0�(ヘ�6Ixu�D�{j^9-�SR:�v�m��v/㫷<Y��a&Ӗ5��zB�i'��P�e� n��?��w����w���_~������ >a;;r��L���<v9{��<���cƚC0Ə�	z��C��s@�zd��Ɓץ4��kHF9'�^�@,����Ԁ/2��/�J`�D�s4zS@��@�PYP���C��f���W�y�]H�* �* �� ���W�0�c��C@���m���)�[e4}�6ҹ@f&���1%�[6v��vB�Vz:ݶ�uGM��4,IF�<�#M9�Ĥ��w4
��]H�* W�c�`n��U�Z�5�7$�~����0P<��v��7wmX����4�$���^e^Y��@<���T�e@:� �L3�H� Ȇ�i�@�����Z�3'��6"woK ű�-6��	8�jL�;���-}V���w4�����7q)m�y1yj��(x1e�&��Wl*&v�훌5�6}p�E�Y�^��P�H���T�w4W/�����&ӆ�m� ^e@e@� �.����07v��wt�/2�
��?~��Uub��<�͔�?[)�~�[�yF�r
���+�{��V�V�fVg]� �ם�dQ����s4zR ��y� U� �g5y��V�Z z셺"�Z� Z@��n?����>�8���x���#�ÕZ��[���o� ^e@e@� �Es�e^�ٙvfi ^e@e@�4l��v_-kX�8�jL�33-X��,��gu����d�����5�h���k�h����f+]��9[���0j%X�OH��{R �* �� �:*�lveZ�W��C�d�����N�ZY9�Ew/��qfL�f���Zy�ݪ�n�v�ڐYP�H��ǑA�9�Ĝ4m��-�M�j�-�M �ם�dQ�o��j �� \[�/j@e@�b�Lm�"oCR�ՠ[� 
��ڐ��+��*��/j�2�͸��VT{R ��	?��W���E�&�cYcs��]pȮ��#UU�@T ���	     [}�oH7m�Wn���i�[qW�5�f���A�=��m.�h�Pf��瞽����Ҫn�ݮ�u+7h�=6��{��:��1�I�u�ㆷ6�qv�\�I!�ۋ�v�g�ya]�Q��n��lNsd#��!�6	���s�]�p]N��\��4�����.���{�ܱ&�^���r�ӎ�ZL����sǧU��=��:��n8�8�uF�2�i�>���� ^Ԁ.-�� ,�\M(�6A�G3@��4]�@��4m��9[���0j$)�m= �p�H����ݜ�V9��I��9�oJh۹�[Қ�ՠ~�[�yӐɌI� U� ^Ԁ.-�� |���N�e�@��+�='Tt���E�®�Z����w��SR<z�蘁xxsJ���a`fNc�3;XyBQa�����/�i��M�hjC@�ڶ��*B�R*�B��GR��8s>�,grՁ�������:��S#Sm	Š[Қ�w4zS@��Z�|���@�s/4�<��ڐ�n �� �Y|��SM�jD�h���z�h���z���U�4�r"F�I��z쳂��ɥX�0��tn��s��9�4A��Ɯ��"�5Jx6�4�S@��4��h������2�s������@� ,����RR�P��n�ڕN�%�P�H��`nnڰ3;XYP��(ԡ*��ZX�V���; Ȥ�4��	��/�S@��h�S@�n�w��m6���Ya���R �j@YPΤ6���~�?�� �R�W��w1:6���ɴ>Ӯ�	����؀�4�ۙ��\�hn��-�s@��O��<��ﾟ���|ň� �N��@:�u v���W��efe闦��� WR �j@2Ձי�*��M�PL���a({�zX�ZX��V��
'2�윕�U�c0�x��C@��4z�h���oJh�q<�1$�Mbē�mY�s^�v��9�xӃ�{m���7.�G6y�sE4�2cp�-빠[Қ�)�[Қ��;#Y�F��3j �� \��ڐ�T �R-i4�6��5!�Z��ޔ�-�s@��4ʬ3�H�28�ܱ�;Q�r��7wmX��,6""ݭ�`�7di�f�L��˚,ŕ ^Ԁ.-�� U~���]s�U*�U�O���h����zB�.v�]�һj l H  \�@lRi��[i/gF0e�!�w0<q�p��F4nyӳ�;m" [ĝ�����=a�q���ڮ$��y��;�ARã�q��̙u�ك�ee����&�m^rv.��r#�\�9f.;[�=��v�vݐ��U��<�=P�\�a�؊:�j�%{��#Z=��@eZ�W�e6�a=ZM�=K�s��x�݁n�d�qO:��]�K%�����w��.-�� 
��k�Q�Rr��	�4X����!$ٻ�����j���a`}��,jiH������p�H����qn��LڕU*IuT�)�,6!$�wx����@�ڴzS@3��dk	$yYxfQy� ^Ԁ.-�� n��j��V��&�R6��#�n���\�:z"�3�����vl/k���lp��*pM�h��k�h�S@��ϼ���kK�6[�5S.fX杁����D$�J�&d��Z�9�XX]�@=��֐�Rn8�p�-�r��@�ݩ ���^^љ�ze鹵 �u �p�Ԁ-��+|xRLMA"xcn�ՠwv��e@>]Hr��\�����S�]��t��g�/
m=�wI���vU�ɷ2��Z���߃�a�c��$�?#�h�)�|��˩ ��n��̕����^��maw�@>VT�Ԁwg7 ��M���������$��&&��hn֖{=�gVE� MG�v�M���k
����4X��bi �nSI�h�rVa`j���H�.�D�ʰ D�@�c�����G�,���A��I�4��	��c?��h�#s`��(�H; �B(K eHUV)#cD P��T�P��F���B\�54��HM�7��kY0��n4������r I�H9�̒�6�X�J!CQ�+����tB��o[��Y��%e7��ѣAHJi!tA����0$?Z���T��&�i�2WX�@�30$
��
0#�0R}F��X�$�A�A�+���	t�D#�C������:bA4i�E�9 � j"%A�^��?�W��*
�W�7���g��w�nhz�h�Hn	�m`�4���ݩ �YP�R �tW9vU�H�m�8���?w]�����}V��^�'�D�`�m�"Q��x��aV��j�<'D�r��y�c=����\�l���8�bs�q��~�e4���%
8�3+K�Rljr�3.�a5J��@>���ݩ ��� ��9��$Om�@�Ϫ�;�S@��w4��h�a�c��$�?#�h�k��Z�9�XXR""�4��$G�P�%s��vnlͩR�)�ST�nh�9�rՁ�b;�� ������������?�]��k��U:�x֖vt��o�N�q�h嚬�6;����~��T�%�i|}��`s��v{���%a�_�4�G�������C@����ݩ ��ʀ|����WNeيdj&��@��M��w4��h�}V�{���#� �#����XX̬,}=�a�'�������j�t��.��f������J#�wo|�ﾟƁ��S@���<�vInI$�J/�VA�j�
ҹ��QV ���  ��p � �`�{k��hZZ�{����mt�<\�T�tg�Y�.b�I�m��C/Y�ݵ�/g\"m��sUь��^�J70l�xeY\��*1�"�������we�R����=���l]tma�WC	O��T�Нl����|<��4���An�N'UCqډ�_��=����伢�)Uk��{b�	w"Vu\<���w�y�[;�q�Z%x����4�ԦʁL���;�Ԁ}ݩ �u �r��6��wbb���;���"G�N�׋��x�?wJo��G�����8�r,�Ĝ4W�˩��W~]� 
�� +�,DJH�ƘФ4>���oƁ��@��M�^ۿy#��CpM�k	�,w����J����=��X���zԦ� ��ȓI��&�9U;^������+h������Ў��.+_���ݻ�;��k�-�ҩt�e�4|�׋��a`s2��^(QHwg|�ǽ%����fk.��nIϾ���A�J��?��0"�E�	@�B��9��`wg|����������Q� ��s'ο��֮R���L�`g����9��;5$��"!��J&wv�Xݯrr$1�'5*ٌ5�dܟ�P�G����s��w$��_���aa�	'���`w'e�kSJDTЦ*j������?D%п
#=�À���?�@�Ϫ�/�&�V��D�u������x��r\�q�۵�4��Bϼ�<kT�y#�nE����=�|X̬,v{�R\a�������l��M�T���luG ��i~���Nk�72��9����S!���2�3C�S,&��;��vw����P�(P��R�:�4Ƅ�!R]FAX:
�pW���\�=���{�g�����L�*��ә�9�a�(��/�IW�{�Ł��~,�+�
�/�QY�{�_���!����.h�9���^""=�珀�������#����+*��ǵ=s���v0��ˁ+�&gl֩&����2Sʇ�@��o�q	�Đ7@�����?s��)��%�BI@�	(_Hwv�X��Hy�Y�ٌ�ֲnIϵ�n�ª�� � JJ���W���z�}���Q�@�S2{�_�R�kBf�sY����W���{XY�$��D(��}��|��Z�U�y#��H�x7�"�"IOwy���z�X����P�P��n�ŀ.�l��M�T̩rKQ`g�XX��$DB����{v�X�Қ���Hc�O#r$�I<���d�f0 \ͷ����S�Gn���^.��b���{��ԉ�m!�&�C�:���^�K�Xl(�(��=����Mze�T���hN-�Jo�y�$wY�}�O��Nc�ℼ�Jd1z=�!�.�˗4X�^,�+=�z%3ܟy�ݯ1I���t�2M6幢�a(O{����gu���	(�DD�o<X��Hy�5*YPI3E�ϧ1��ЈI$(!(��<|f׋>����ߟ�����u�B-%�����.ێۯ*���  �     6�#]�G��T�"�� E���3��pe���
�2�B܈&�)c�<�Sn���5_$�L�HƉ#���F�/:�u�8z���r�<�v�3���ۓvy�m��e׉����@�#sz�5�������G<��s�{v;7�GV�Վ�����fQ�l��]�s-�{�ߝ���p� �J�lFY-��<n�Ӯ4Ko3;I�kF�����L52SY����"�	E�9-�M)SB���z�~�$����ܓ����G�b+ �D ! ��@�!$$���������jUT�����A3E��ݬ/|BI" I!"!L��W��>�3��/c���A		
d|�����fT�$n��=��>��g��_�P�W�z��O���"Ѷ��x�!���DD)�_��n׋�XXl%��g���׍ޖ�RMT˙�9�`g{XX�%����7�ZX�s�s��i��w�QW�q���X���6Iv��.���<���:��o������Ⲕ"M����ϲ��9��=�
<�H{v�X����c�&�r��`g�X_C��� �"������ͯ�v������"!%
d�O�CΨ�i�P9nh�;��;;��͈��BH��!
g3kŁ��x�3���;Ma�L�MHf�.����"�$�
I	D�w�,ͯ}�����"�*B$R������;��n<�7#����4}�M��!@" �"^�s��w'�vw������p��+��@�]�R�i�Z�Ա]��3�lv'&�֭�5�?��w��v����	5�N�Jh��s*\�7T|�����Ә��k����+K ΍n�2�3C�S,&��9��;���%	~""*���~,�W��ϲ��ICf>�-�[U$�L��c�v�V��v���B\���BJ5DG9W����Nk��Fd��ꉗT�˚,5x��s7�,g�Łϧ1�j�	D)��<X���&����3Rܷ4X�V䗡D.����=�^,}�M�U�<K7&GNH�m��m�Y�L�X�0��@st��g��+�c��w��������(Oғ?�?�Z��=��4��Z�*�<adr����a~��%&f׋��Z�9��;ԗ�"��y�Ԫ�SS5ST*�f�3kŁ�fZ�aG�!D�r}�`{v�X�'ܥ5Nj�J�$���D)�{�+�>�3��,DBW	$�4�"�hX�T�Ī���@����h�Y��M�7�6����]�@�J=
��������ϳ-X��c�������7�&1�d���vq�fM��N�oj�e���.R�k5l���,�C���[U$�L��c����a?~�;7$���g���1�D�Ȅ�B_Hw'�v���H4�Q2ꜹsF䟿}���"D���HI	DA
d�{֬��������P�?ʰX�Eb� H�Eu'}'�ɩl��I�ܷ4X�zՁϦՠ^�M�zS@��*�x�<.��7'��E ,��D�(I"$B��_��n׋�XnO*��!�Ea �@׳��X���/554J
��`g{XX�(�$�~" ��-�}�����V>��`\e�*HQ�8^Z�J�P*�?���SL�e�.�L�К���0 Y.��h�J��a���BI$BO��6f�����#�G�!X�_�7N+L�0W?�0�
�#6��_�ģ
�#)
b!j������D�ec�Б���@�1f�I��Cb:`�̈́�@���#[w�|��j�������H.~��P��o�����P��L���HkSD��#|�$<�(A�ĂF���@&����lq��a
$�B��<[��U�?D�4I��"BHiC�ŀA�Yy����p   ��| [@      ऑl��t^I}��Vm��jam�j�<Yh؀j��59��pE�*�>�J������p���U���3��@������`��t��    v�  m&��       m�     �     �     m     $X6�      >8�    /{C��1�8�R�F%��vǮۮ�6��˳]]��f)��BOD�a�tv������^�(����*:Ӳ�� �m��v͖�uf�XGҪΊ���n�ؓ��ՌQ�&�=la�B�uRe�	�&�d��6�c���ֲ�Z�).k���'�ڮ�ڲ�;���r[mn.D3c9w�\=�q�{*vܳ[�.һ���f�P�v��5��f��Ƴ�cf�47j]ٴJ���Z�`�T��m�0]X-�ۧ��t�NMκ|9콫���S�y��uEsm�m�g���x��bn�մ�γ�&*�I���ĝw��ŗ���ܽ;���q�C��
,Һs6;��\�������mO7�?<��i�y�U��&]�m`���� �izyj4�O-V��+%��62to=ـ.��Z1��U�;;#�Y"+�5���vc��a�*8|��I�^:��`c�]��u/4�R��@ϰ���Zx4�̏mkd�؝X%�	�����6���
:�������tP7-Y�s�S<�i�v�g�ܸ��������+���>�����Qsڨx8uMP��XN+���f�ݢm�ԫ�7nx'��ja�ݗkkq�n��f�(�GFb�gzɁѶꃷ2U骚��U8:]��g��j��t�n	 $5�W5톓AmU�ԅ���ٹ,.u7lj`�6�=�[SJ��'i�r5R�6X6�e�`�}�>��4�Ս)��"f�2d���a����D��Dڿ�tAv(��W�� �W(5 ��*�õDT:o��fZUU$ƍ�+� ��ۦ&�^r������ 6� �  �( ��g� �Լ��c��y���R��%�g5��ñ8�7�q���zay�-A-����3�s��r]gوv�B݈�c��U;@���\p�]�JJ�:�m�ϛ=V����܆Ŏ}[Llõ�����˂�UA����H9�]��)ג9�O"�^�l�nW��ۘ��mY�r۲���#��mu�gۈ��8�]sԴ9���w��ow���~�]��Y���{L��?{�~,�2Ձϧ1�B��̭4=�+�b��LBR����G�y(Q2w'�v�kŁ�ݬ,�fK�ФCx��h�v��Ji��fb]�|hw�nhza��,�qF6Ц���	=̽,�+K>̵a�BO�|���>���Rr6�p�=��4P�{���>��;����wP��@eR�U��M�5����n��5�-%�y�)����kn/���V��q�k��-����Ҡ�n �� s*��ꉖ���庥`gӘ��!B!
�UliB(@��ڻX&h~]��i?���1��!�M��U��R���@�`Vb���yDF����,�}j�ϻ��b�%&��/55*������mx�3��VjK�P�}��V�kŁ�;K"�S5ST*�sE�!%���V�kŁ��aa��%��x��O}Jj��8�bi�3@�۹�~��/t��}��h:��Q�Cq)mb�Hc��]l���ԍ��K3u[&Gċ��������d�E]�s��e�U)je�����`g{XX�d��	B^Q�D	BK���~,�!~�Kj��u$̺sE���a{���!!(P���o�Ձ��x�9��h�|���Rr6�p�-��4'w;78�T� C���D��/��� "AUX"0Q�0A@�)A���������}����^dbr4R�6���+�!B��$�EX*������ܓ����Mn�o}��r����  �A(I]o�SM��ކ[�ҩ�MUCr���[l�����oT  D��RK{�i޶ߞ�mU��ϻxs���g���V
y�
�r۫y���.^��9:M˻ip��<y����e}�;tsy�=F�6~o>���6�Orꝶ�ϻxjJ#�P�	!DB]�6�v�.�m����SU4�Y��WY9�m���.���,#(�J*��fߎq��v�.�m�ݼ9�QВD(@�UT�羥5NJ�je��fj��m�fߎq����K��$���r����߶E�$���-m�ŒcX�$�-�W�S��Aa7���jn�o����Nr�{��y�vߞ��D>��Q��_�q�ǂ�Kj��u$̺��M�m����[o�W�@�
 �s���1������9���s.Km���q�R�U#T��z�m5��9�V{Mvg�N-��a{rX�m�b�^��g4�[~�@��]S��y�oq���I%�"!}T��m��m�NF)��n�MU;m��v��5D/"UT���e���m��k��"߼���_�F����A'�4�?~I/��Q�$�����$�۲-I%}�Üm�ɩhX��J*US$uL���(S;��9���ݺ�m���9�ޤ�N��m���-lSU4�j*�fh�o��uN�m�BQ��i�ͷ�ݹ-��}�Ün��{�����`M]ZuQ�ۗ�h&�V6�qe��)u_��|� @ ]�`�:�rnmh	t fm�����qu�s{mб�1,LA���c�l��l�0�Q�(v@����q�\K��5��z�B��9����n��;v����;0�Q����b(�B�&�֐m�=n��Vv��s��V��,s��Hu��e�,�g��?��>�TC'�M|}�t&�*�.��ฮ��X�N+�:���M�lq]4j]Y�q33UO���Ϳ�m�9�%��ϫ1���=�����RI/xY�Ͷء1�m�9����[/b��o{[��m��Z��I+ݴ��$��Z4�1Ħ6Ԏ3[m�՘���}�b�m�Q���
!]��z��m���r[m���̖7Q$�L��>q��^P��w�T�߷o�8�Ne�m�P�L�ou��L�NF�JT����$Z�J�m?~I+��5$��Z�~I.?>�����g�u����V�s�����LB�E�����:'=�9ذ[��p�;���b؍Z�H1&������}�ԒW٘�����]S؈��os/Nq��f��k5���3,&�57-������ �?�D%wn�2ꝶ�����m�k-��DyB_�v�~=k�SU4�j*�]S�o����;m��v����"!]��W�e������~�@��~~WR�̣�Z�����8�y��e���՘��ި�A[~��-I$��?��m�Bcx���~��W�-��oT(�$B����������m��m?~I"�R�6d�N7"M&�y1��nM٢����Za��������2�����:ݺ��4ێ#RI~�j��$�۲-M��{xj�QQ@��m�k��m��l{Ħખ��e7T�����]S�Дz""?B�D(Eݷ���9�����l��|�j��$�3�������s"Ԓ_��}������ݱQ�T��Ub0� !�?�`�~����y����N�m�fs�U.FBl����ʈ�*��3����f�����8�o;X��m���Üm��t��M'4L�2�K�f����o9m����	$(�*��ʟͶ�v�s�����[`��������*��ɬ�,Q<�t:Kn��ۮ��y�����VB35L�f�k%f�%?����D,R��8�.f�e�0Թ�������S��w��8�y��g���o���6����I�6H8�bII�jI/{���j��_�P+��_���o=_�>q��v�S��B^I/���m�{�����2�Z&��o�����m����y��N�I{ݴ��$��Z�23&&ێ#[z�^Uwy�>q�߶���m���Üv�����~ Z��������ݶ��ߞ�����旂��� ��ߝ /{���$��u�K�KW��$���N2�������Q�;��Gnͦ7.m�9p�:�npp�;��{_k�p�k��C#t��o���8�Or��|�f=���[o�Z��m���!��L��hM��q������D%
f[�wvy��}��N�m���9�Q	(^�UO�}2�檓%JA5%����ޞq��ݬT��{�Üm����RI~�/�b��I�q����3&{�������Ӝm���:�ߒ�U]�{���@��?�Ժ�Npv� ?��~��K��=I%��_��${��5$��;���￟��u�`���i��/Y��]�Y4�:  m� 	 8  lR����\E�+��sb.�R>3v8;.Í�v4E.�n������{p�ػ$��jy!�m��8��ۚ,��38M��f��t�8ֻdX,��z�u��g.�܌!���g�-�6��l�E��*�����u�����V��\M�{�k�+s`zZ z�M�m�p�.f���zA� k�.�c�Y���?c��W:��S���7m��m��'���6��K�Ԓ^�m?~I$����$����M����d󟒄�����^E[m�ݿ��>���$���B��ޯG�����$���:��m��m���oq��_U5$��ֿߒIV_.& ��'d��N��G�~HJ�}��9��6}�ն���2y���I~�+��ߕ;m��~�C��c8bCN�$��ꦤ������I/z\�RI{ݴ��$��6��NN �J�v'[����޼N�ٖ��kg;r�b�9�\��JyC�`����af��jL�2�Ͷ�;�O8�o��*v�o�������;9�jI/iw>�,R5	<�"R?ߒI{��]�X�?%CdS���I~H�K��|�oq�̝�m�����7�����n�wTc�����2��c R�m��v�s��}=�V��	L�ӻ��4��>ȵ$��賫m�)�6��~�o�"���T��[m�Ͻ��m���������$/C*�FLc�0lQӫm�����oRP��B��|S��������I��jI%���5V,qFܑ)r�N{�x��9ll��]�;V����p�����x�d�ݫ:��S�� ���� >���8�g��u�yG�L}�{�`��bch��'��&��қ��y������̀s��V�Cʪ��Bn[�,���8�2l�ġE9��B����%"�cX��k$Ed�դ �X#`Db����\4%a$i+Y�TC��Hp��BX���c"A"q]*eR$�� A�X�.�dM�hW �,a	t~Ӏa]�DМ��~���0���!� 0�!ed��;Xq� ��>��}�� 0"Md4���R"���U�$� ��_����$,�V�+�v8:"��*|�@ >��!��È��C�(�D�
�C�N���lo��@��xeY&!�&<"R-�ġ?�wf�>�iV{���В}�f�ߋ3�"�#P��2%#���&��Қ���@���@����\F7�&�l��6w�s,�q�=�c���;p��F�
<_y�Z�8� �KI�~�>4���8�2|�=���*�;�[�m�)�6��h���� ��Rh�)�y��3��ԘF(��=_}����&��Қ���@=��0�d��#�C���4�}7$��_v�C-�]jV$@!Kh@���	��!7v��"a�R\�!R�7d��Ŋ,�' �#��{��$��y�u.���9��3TU��{XXQ��k�=�z�ޤ�?wU�<�L���rE^��̖^Q�q�z�9��7g��z.9kQnM]��z��<{b8bM'�w;��?.���z�@��S@��xeY&!�&<"R-��^��y�A�_��u��@���h��/�b��I�q��z�@��SO���K�ߖ��|�
����#� �KI�h�Jh�����^��g�%�_���e����o@�4{9��ː�rl�ڐ�~�H;h|�b�41J��������Qlk(���Uז��v�X� ��� H    ���u�D�t7^�.x��D�%��V����vc��+�/d\�SHi�W2�oeg�c۬Vq���Z�X����zOI��mvx�cr��n8�n��OV�O�PQ):m��V�N���q����Ʋ��=JM��Ў
V�`G�us�<ݸy���W�/�D=�{�����Ђ�J9]��;w1u�lu�ǎHdч�u�\ys��䗶���.����*EK�����9�aV��a�"z�����>���A�F��= ��¯�&��V�Ϲ�`q�2oT(l7��>��Ҙ��'��M����W�~]k���M�+ǎ�BJ[�,6!'��6l�ǹs�¬�ڦ�y��ʲLC�Lx���Z���sUp�V��ɰ3��r��	��8��v՛�-��xz:����\!��8�a��t�b��5C�+7�I��������8��N��7f�͑<�J�F���im��nI�ﳳxQ����+ ��(�"�B$*�PF�
�EAJ��A�<
��.�e��u�r�@?{�&��$�"�M���o��=]~z�ֽ?�H���4�i`|���LSSIԺ����ԡD/*�� �o�X�zP��f�>]�cň�F�H�5"���ɠ{�~?����?z�� ��I�"ƒq�Ԉ�z���f�qƭO>�����(nc��됷cM�)<���S1��2h��M����9����������ԍ��$%P�]�����g7 >�5��ړ��7'fP����ER�EUM��gu�>�*��P��Ir"�~�a`|��60�e�$H�$�LQ��>�/z��@��|h��^��ՠuf.�d���KN�U���XX��Q����d���9�s������TC�4g*�[Hc΢��8�褭,����d8�;H���_a����(��1�x����{����Z�޹?���	}!���`c�^~1T�S����1�>�*�>�+���ߒ򈉐�����U.���sN�37ʬ��@>�.@=�[�
?��/.��ښr��*��(�Ng�����zl���¦"���_w-U��KČ��la*�幢����6��"3w�> �o�X��h��B�DiĤx�%2a��V�"��Q{0/%��}�8�xv|���u2�e{tup<$�I��t��~��M�YO�? �u���Y�y$Jd&Hh>�*�9ܬ,?��`}��7�'�t��L�t�M�T���z�Xw&����h�z���GX�m�F<o���)̽�3'|��f*�9�V��ʨ��I1H(��=��Z�����H����Vn��fn��)qi�5u��L��v�5�n�@&�Wm@m��	  ��6Z�N\2��*Ⱥ�^���n{en�y�!*5�!���;o.�p/.x�k�2}��v�nD�v�6�q���&��!��l5:u�n�c�&K�M70gC�&4u��S�NB�����;�¦#.L\��x3��o8�k0g�]Mt�Oe�lo{����Ӂ�J	W�8v��x�Ʃ6���� ���7!m����Kz��K�$�����s�}�������0�g5�i���t���yW�����@=�[�{���{nM�;���� y�N��T��n {�[ �s*ݎe�nՙF�i{� ��n {�[ �s*�(�����7L��M�M�T��T�8�-l�̨��p�����8�뛲�|}�t&�&�S4b���齶;Z�X�j;b��n(��[�{�� ��*�b��9��-l �$u��ڄc��9���V����ȡU������;�n�I>�ޙ�;�r������X�S)��SC��`}����Y�7�͵`w����w�Z�,$R$�"�}�&�����=�ڴ��Z�����S1ŕy�[ �s*�b��9��-l�~���~jݰ��J�k�9�R)�x���6�����';�y�#��p�<��&���iw��� {� 9���[ �s3@�u�2���8�4��Z �k`�e@�H^���ٻ{�T��T�; ϳX��jƒI		%Ĕ+�U�����'����}�J�R�"K�4��?Wj��4�$u��ڄc��9��Ԁ|�� |���e@=��^�1��*�s�vn�&�GW=X�����`�Ϣ��5��R4Iʒ�VÙғ�>qn >Z�w2�v� ���V�K		�A8��nM���{�4�ڴ�:�&&��Lq<M��w2�v�������Jrj�������a�'��������YV
(��E�%٬�>���5T�(��Nh�9���B�D/�~��~���{��3+��s2�Q,�N(�N�h!��sv�]�'V�e玷f��۞���˴rr'�ȑ"�$�L#qh�,�;�� WR�p�����n�^���l�UV{ܵ�~P�O{������@-�f�_D����P���Nf�����̜�f�ٻ�j��͵`u�3��Q"L�`�4�ڴۖh�w4l��~��X%���D�杀fbʰ<�%����7v��9����8���UaX�#�� �P-�V�%���M�	�l`T]H̒P"%�b�tI�"�H�I �J�F���0 ��Aݰ��(ēB;��333333    �      	$ڈH�4f��H�N����ghn��5�� �e�`�r�.�I�¤����<�:إ/r[J���Uj�U�)	Pnĵa�v�e�kX     ���  nۦ�        l     �          	     rA��      8    ]7I�m�v6�U��ƞ�j�X{9���^�R�:�,����3�g U�uT��^
8��٧b��嶭ú��S��]d2c5U[Td7$b����qO����F�Tܛy]۰��]Z�\��X�kA�$���Ӌ��re<���;��I[0�r;�gdoc��e�&�+0��8��nls@66s���O>{mSj��Shɵu����g���5���ם�ד�4V�^��6���VƩWt"bpc`����Ƈny�a`��ln�Z���8ܪ�Nd�n�i�ݺW� M��qq�rP�1:.�����VDا�嶶�Wn����G6��#���H�l�uJ�3�]�=��܂J�$.���5���j�(7�J�Wl�����ɳC�G��K;S��s���T콶s��ʰ�^K&�-���Άs����no[��<��z1�[6�ɒ���V�"t0��v�������KK`��88�ghm��$��P����]�rθi�rM5�$ p�,�0��C�I����M!U95:���w\\�v9��-$Pr�EV�Kj^}l#u���۳cIuL[$<���s��"���^����(���qڞkn�u�s��!챌��\���A90J���mSm�ڶj�k�m�W�61T��qD�ƓrkBK��[��ct�GD�jɲ�P-Grm���T�ʆ^M�1Yu���W+.�l%MՀѻ��
қM)-UI���BS�&���N�{��w�;��_���ꀑ@�x��Z��D��N��M�ٙ�����n�x����t-�nRJ��n ���  � ��zC��E�.�e�z�%���;��pNzl���Pd� x�Yۓ^'�-	<��le�v������\vۦ��%)S���F��F�M������c�!�{��/F���e�z뚏,K�ϵ�䱧:E�b�k<e��؜T��j'=}�W�@��0R�������u���Py�<�m�F�+ʏ$Succͫ�����m��T]H�-�i�]�V.F�������S@�_U�Օ`w���I�읙B֪�%R"i�c�pZv��T]H_J�cd�)QT�MS�؈P��յ`^�nh�M�v��w��2G�d�wWf�n�;�� WR�p\�@���Hc�O#r$�m�0���\%\��m��_���b��k�a��k4�$P��l����|h��h�,�;��h�9P^E$����?w]��M++�>P��R D���,A���	_��S��2�
�@��s�E�j��D��Zm�4�S@�]�@;���I�1d&%2M��Pu 8� �`_5X��H@�	H���)�~�ՠܳ@�빠~�Sm-c��ē�(�y;����m	�x��e���\���ȝuּ��v9�{tu1	���@�]�@-�f���s@��h=y�T�0��1F������!&���V�֖2s�����L��"K$�4�SN��)SB��d� UBQD\BQW�M�ά� �|w*f���2��LҰ؈{�zXl� ��w]��*Ȉ��BSH�-�i�w2�
�@?����?����q醠��Ӟ�-\��;�6@�]�:"�ۅNM��Co#!����tQ�D��_�>���h�w4l����V�wu�&�Jb�LJd�w]W�Bl�����gu�f,�g�r1b�JF�h�M�v� ��w]��:��Y&!�Df'�9��31eX�rՄDDD�EBP�������R�1I䘣qh�-X�rՁ����̜�`l%w59\n2�@� ��f�fÛmnI��8@��;`��Y�®x�]OP�w��� WR�pZv 8^U�Ԓ'C`���)��${��v��j��{����^�U*f�f�w�@>qn +N�;�� WR���5���:��T�i�jI7���`
�J�+� �Ÿ��뼻˽���j�kv�̨���[�ܳ@^yg�d���bJI$��$�`�Y���l�����@� m� H   ���h�N��mj�.t�cp��
�r�9,܉����
i4n���ú۔�uӰ����3d��{coS�'�WS���ˣ��A]���y� �/fۅŲ�t�[]�:�9�[��j.8�	��ō��]mp��=6�#\=�K���5,�*Fk.��?�C� s[�-�,�3&kPD�ײɦy]��m���v3��:��Z
9ɫ���T��5�
[�6������|�� V��ws*�cu��n՘���Ӛ,d�;�J!��յ`ff��/;V�sם�HsD�G�7�^i�w2����obh8� ��߯��h� ʚ�����+;9���Nc��	(I��[V��u2�j���4���;Д}�����j��{w4�sc(�&�q)m��^�v㇄7	�0�N�.ݰ�X%��V<E�맖���ۀ|�� y�`�ʀ=�p^�Φ<K	$y"PN- �r�^`�S�� yrw9훒{���@�]�@=�$���L�ĦI`w��Vvs����w]�njڰ3���#c��1�H���h�j��,�/u��?s�U�b�c�v}9����5mp��Vvs��,���>R	�曖�mʤ �պ��og��;m[d�hŎ��sԴ9�r����)<�#n/�_��^빠^v���Z�;�t�#�2D�$I�h��W���=��;�>��,� �=����X�'3@��Z�ڶs�B����-�V�F(P��B 4�!V0CxEP�8�@�čFEGA��
`�H�,	B1��L6��	@�~|2}�s٠w_�4ɑ�EG. ���; {�P�n��Y�ǉa$�$K"qh�hy�[�������/�ՠ�I<2ō$�m(%^���fm=v)*��=�1\���u��됷cM�F�<I�5<jd&%2M�]���;>���P�����ؓj�IU,�#uS4���;Ԓ�%2{'�v���X����jV5T�(��	S�3��v��U�	���V��3ם�Hs�'�dmŠ���]��;��۹>�@�
bw��.䟯s�����	4�w4�����������fa�`|�&e�yL�8X)T��C/u\�����[�	s�v�;P��4��<Q(��b��9��k�3��v��W�J#�73mX�L���"� �-��Zm,�/u��/;V���Y�ǉa$�$K"r����� {��n w�s)�u�Q@�T�y���X����ՠz����|e���h�ĲTҰ;��v�D,��|�ul���蘭���඀j-Y7S�/^�i4k�Ֆk�p-���p� 	�� ƒ�'��ҙ���<��]J��5�ẋ�q�u����ϯ;�����D�Nם\�<aSy.��rt۱�^3���8d  �@���N��
N�����;t�.�kə����[���5�0�G7�۠�u����,��7;�8��k3ʯ+ә7{��ww{ݦ�|�h�0S��]v��j�dSs >���x�.9��>ո�z9Y_2s��n{\]��ݿ��9��i�+*݋p��db��26��=V�z[w4�j�:�V����v"G�d�]^��n@9YP�[�s�pZ�����#��Cm'3C�[>�h���@�[��m��/tE0~LP�D���:�V��+�:۹�w;V�~�Z��"Ȓq�F�m��4���8��Qms\��lue1��N�I��+4qչ��IH�D��=V�z[w4�j�:�V�w|M�Ƨ��	�z^�f�x�� 6�+�M�]��_U�z����|e���LbY76�ط ���� ��ϸ�*�)E'H%��a����:����m��;��@�;ʐ�F)<�[��pZӐVT�����~�����4�ƾ>�N�Q�J.��\N���v"���gD6����Ľ��}���戒���}�����w;V��ڴy�^�v�����i6�s4�j�:�V��:��:۹�bG��|`���R4Š_��h�;��.g�sA�D	uJ4b`b@��P�%֋	
���j`CH�!��$��$��4�@$t�� ;Y!��P�54�ѭe5@��,xQ�+�H���X�C���b��S.�!.�[$$@�i&X@�Z�.�:p�'mV0�K
@���@4�@������&�JE?O� ��D�C����V�B�E����'�'��G8(�IF$�C���Z�;��v�]�<I$K"�h�r��]���;I��k��6�j]A4��r� �*݋pqn�Zr����5���J�\��OFv$M�֭[Oo
����;6Ɛ��Ǚ�\���j݋pqn�Zr�ʀ}}�Q���B�H%��`w'1��Q�{�f��ݵ`w�������ɥR:����͸�i�+*݋pqn���t�#��X�S#�:۹�w������TA1	B�0�Wo)d�a�ʹ��Ɠi'3@�v���U�^�׮�}}q@n,i'@���8�f�8��c�����#`GdmŞ�k��B��F�`���$h#�@��Z�i��*݋p[W\��XI$J
E�z���z�h�ՠZ�� �:��ōO	@O#�-�j��g1٩7�9����[6|�"L��%�t�mUM+Q2�]��9���+�-빠~��Ʉ2Dx����`fOq��D};�g�n�ڰ;��;Qbĉ��:g{�kY�k3335�qq;�Eoc�0C4;t�8��m@m� ��t��c���Wn��ͳ��fA.������q�uhq�0��;[p�����k3�6�݋Xu���ݣ�����Sr�	�ldwR����q��pb;f9$\h3��؝��7,<��$�G<K;���Ӕy�A]��:�۬" n��tƄ�{Hf��]\�̳J�X���5��j�N�݆(�V�`�9�h�'n�<N�f���k][w$��T�q�נ�ӊ�q4�o٘�l������
#�7g5�<��FH����o]���Z���?+r� �qʹ��Ɠi^m@;���.sp�i��* �DS��� �A$Z���?+r�޻�s�UŝLx �,�;��n��9 ^e@;���.sp�~����Ü\L���{kQ���ș�nyێ�#m�졇�փ���x佨By�o]���Z���<���纶lꝉ6�d�Mґ�U4��{��!%��]K��/f��=ճ`fu��?z���	����ŠZ���Zr �ʀwg7 �r��vf���LQȴ�ܯ@��������h�|�&E�$�F�G�[�jݜ�qn��9 �9���Ӈ�� �ݲQ���nx�]�F�E�zA�tb62���Z㵒��� ��~�3'5���vb��.0�͵`ne3DLR��TK�T���;Ԓ�M�=ճ`n�ڰ;��;�]�JUSRF��Z�nW�[�sOs3��c}U�Z�Zޝ|M�Ƨ�� '��
������ZӐՏ�,��D�1,�L�;�U�Z�Z�nW�[n�����i~c��ē�(����M��޼N׷6E�F��y�[j�s�v9�t���*	njx���1d���h���;+��Hs#�I�9���9 U� ��r �� ���I�dX���S#�-�s@��^�k�h��^�P��6�s���MҰ�J!��l����<œa�P� '�z����	��s}7$���O��� �DR=�j�?+r��w4]���U ���JF�Ę��E�NG;d�K��e�`]��x9���6�;�,�0�$j
E�~V�z��h}�N����v�3a̦��E+r �*���qn��9߭⹕�����@9wW�r�P�<�	C|y�&��ݵ`s��*E
�Ji�˼܀.-�>�� 
��}�h�;�Ht�Ry&(�Z�nW�[ܵ`u��6d��6(|�J L"KA �HĤ	a0P�J��)���������_��:� �IwF��w���#"�7jڪ�ڶ 6� �  ��rQ����!��[��.z�u��,��ض������N�kbq�uk:�G�N�&ޝ�h��G��ܼ'�Cv�q���=��m�[�gZ�=4N4��2g�5��K��l�G��ͻZ�gJfؙ�sv%�V��j�e�c��%b���5��{�7�=�q�Z8�lш�5�C��Ss�)�{qpv.x9ܖK��)bW<q;p���Bjd|�n�˺���h��^�P�u����Fbm&�h��@9�ִ�y�?��������0^FI�h�G�}�-�+�-빠r�@�pκ�`�L���92�a$��wV́��j���rl��V��r&e5.��(�r�l6���_�*ʀ}kN@suw�Y�V��z�Y4�+���Cpb�8xκ�vx�'T疎(���7�Sˠ���]���~��VT�Zr �*����4�45��j�f�$�{ݛ�2>T�����,�3�j���robQ��i�D�b��1H�h��Ϟ�m��.��m��?{�N�"Ƈ��� U� ��r �ʀ}kN@=]cj9���I9�.��m��?+r��w4Z���<���JJ��l��+g�:ۀ�#'<���R�;�t�K�4C�MIi�)�m�� ��`
���9 ��u�YE�miUR蚥`�,��ٻ�j�י�`ffZ���	��ت�MS�*�)�UV���nI�����#A
4H>
 �B]��T�$���� ��ʰ3�rdx��ĲG3@����w4�r��w4޻ra��s	��q��P�N��P���{�����)瀺��պ���Eny{um�)���D���{t��\S� 4�y� o���*��1c�dX���&I�[�s~�>V����nh��C�XڎB���w�P���/2�杀/34x��yR6�h�G�[�s@4�y�����mUUUe�s��3���0�!$jL���4�Ͼ�~��|�������xe�I��PJ�we6�UVӛ�=m�%���{o1��u�:f)s�$ŐS�8�$�M޻����̨ ��`��;�Y���w[�� {� ̨�Ӱ�s@���d&c�O7޻� ��`̨ݩ �{h���6��f���� |Ӱ�T�Ԁ/]�����2,hqH�$�-� {� ̨ ��`��������ЅV������@���HBI��dHD 	 ��!R�0c!������ڍ��!IB�"D$$!��5��"��F0jc6�	"�FE�HT�)�$@�#1��
� b��"�[IL+���0�$$��R0�C���2Ĥ�ņʑ�M-4�R�$Db�*��0B ��L	� ��Ñ��H) ��)� ���!	�
��-�II��$Ml�a�)�i ��E�t�P��s�ᴊ�A��$�B~�ao���^�{�W�]�������     6�      �d�-��m���II�c��5-来s+vH m��r�����s��C�Z�[i�I���vIAmI�m��BXp�J�lԬ��� ��]���     ,�M� �4�        l     �           �     7e6       �    okl�Id�٫q��������g�m.d�6��^B�^[R�B���+Q�uV���-v�i�:Y�$���pػ�8������V�.�m�UeiG��g�`U7a���nU��gvv3�۳cA/�����Qk�(�QK���+������ 6 |��GX��y��Mm�f�,��%�!�h�Tq�狇`\��2g�$�-�t6���'�@�V�h��ax{�[��k
�ݪV��2�)��dx7��6�k�'c���S�����1��g��nU�;r�ͫ��[�d�4)�YHM5GW[c���u���)�94Θ��n���\V���sr��7Y�]y���U �N�UU�zJ�(���;e(�VE��yҫn���ɛnò�b�&ZU	֝�î]� #!�89���SpWPa�=3�Qq�a9�l��D�n�v3g�2q'NI)C]��=/)Q��{q��z6�=Y��u�����gl��\��a��{ml���Z�om�LH�d��;�Y�U��x۶+��n2
�-��%�8{\=�)��v·���-���t��4�<�3ѝU�-���U7$r��SS��f	6�nNu. �d�l��ǈ�ҫ&�gt<OkEf⸒�*���F��(��I���j�X�(���ft��AS��ru\��2���% e�I`!�WeU�<ۇ���pF�����훳��2�����UVQ�C7��:��6W����{���{�w�?!�C������C]S������{�$�ߠ�h3hKPɃ\�RB�L[kUQ�  [@p�   �`ֹt�]tK^�ڱK��i�P�ݎڷX��W3�D�*���X�En�n�;���[�sֶQ�Zش�[1흍�s�]ln�F�٭��b���z8�^�[it�����y�d�z�S���cO=��4��	�V���� �����<܎��W�-%��T*/�ff��][̳,Ժ�[��qm!�wU-t���)sY[��;V�`9����lp��#j9Fcm��pޔ�;����e�����:e0^Fԍ���n�� 4��ʀ>�H��-Փ�LD��I3@/��h�* �� �* {���ݫ�/�u�y[�+* �� �* >�f�}�|e��dIO	&h�S@��Z��U��fZ�5(�Qݬfʡ��4�]�w������>�v��\��;�t�h�++�n�Z�w7k��o����vՀgز��2��DDq��V�V�&����.�IH��V�bʱ(™>�P�BiDDM�v�������Z�?{Ѭu�,x�b$�4m����;�����4�.��������ͨݩ �YP�N���������X�)h�2�\�a5E��YP�N�<��ݩ \��5��2� ��8�&�ӹ����!^;��9؝�S^e0Vh�;f�T֫�杀yYP�Rܲ�{�$�AO�ȓ�4m����;�����4�;�,�"�A$V}����s-Y�S����ڰ;���}=ȤQE%4e��$�����Ձ�fZ���z_�L��L��}h^l�)K�RR*����	���%��ͧ"X�%����ND�,K�w~�ND�,K���m9Ļ�ow����U?�]���t%>�x�'k��:����y�9�ۮ-K���m�c����rkY�e�p��r%�bX�{���Kı;�w��Kı;�{�ӑ,KĿ��ٴ�Kı/���Z�����S333J�p��L��Yܽ.�X�&�X�����"X�%�~����ND�,K�{�6��bX�'�2ֈqS55-˖K�.L��L���p�r%�bX��t�m9���������"X�%���o�m9ı,W����b&�*�j��W�&Bg��D���?�iȖ%�bw���6��bX�'~��6��bX DW������ND�,K���L��2\fk)����r%�bX�w���Kİ�AH�����~�bX�'}���iȖ%�b_����r%�bX��{ut{7�X)U]�<朻Ӝ@�Vjٶ�+L�bs�6NǞ�:��F���]���,K���ߦӑ,K�����"X�%�{��iȖ%�b}�{�ӑ,K���w�2��1���M�"X�%��}�ND�,K��Ofӑ,K�����"X�%�߻�M�"X�%�Ӿ�R�f�5&f��r%�bX���{6��bX�'���m9ı,N���m9ı,O��p�r%�bX�������h��K-ˆfӑ,K?��������iȖ%�b{����r%�bX�w���Kı>���\.�	��	�cͩ�STU9jgZ��ND�,K�w~�ND�,K���6��bX�'����m9ı,O��p�r%�bX� �v�*�x���lFX�,8�u�7�6se��\�n�[P �`8@ ��UR�T�6�#�î
�e�"z�-��'b�ns[mpX���ǟs�%�q�&'F���q��y6��	�Mq�F�)K�y��u�oZF'1��ӛOn���O�z����i��#y�㘧$/[#��Z��᫜�Ƌ/���2&y�����i�q�WF�)��]ri����=�����PTr-
���voN:kc�g7&�u묎�.lt�)��b�ZzݏK2�W2~O�X�%��{�ӑ,K��_{^ͧ"X�%��}�ND�,K����p��L��_OS[����L��fL�6��bX�'����m9ı,O��p�r%�bX�����r%�bX�w���O�ꦢX���?�\�.33)2�Y�ND�,K�����Kı;�w��Kı>��iȖ%�b}�w^ͧ"X�%��y��Z�fj��6��bX�'���m9ı,O��p�r%�bX���׳iȖ%���MD����ND�,K�翜&e05�cu���ND�,K��m9ı,O�����r%�bX��}�iȖ%�bw���iȖ%�b~�wt��kc �D���j�<��k�׬��Hf���|�5�7\Kיח��ey��iȖ%�b}���fӑ,K���ND�,K�w~�ND�,K�︮L��L��VH�f�jT�H�3S�ͧ"X�%��w�6�����1j�ߐ~4��ċ�8��"8&2��6lc���#�?�!�� �}�'9��M�"X�%�����iȦBd&B��gj�p��p���O�n��]UUM�̍�+��!2!nm��\�bX�'}�p�r%��	D�N���ͧ"X�%���p�r%�bX�i��C�����d���p��L��Y���ӑ,K��_{^ͧ"X�%��w�6��bX�'~��6��bX�'gY��0�L���*�\.�	������m9ı,N����Kı;�w��Kı;���ӑ,K�q�~~M�|��`�U�s�sO�6�a����J��=��4�j���r�h�ދ�52L��fӑ,K���ND�,K�w~�ND�,K��m9Ĳ!v{��p�Bd&Bd-�j�D��ə�ӑ,K���ND�,K��m9ı,O����r%�bX��}�iȖ%�b~�;�	�Ld��fk�"X�%��w�6��bX�'�w��m9� $>X���Ћ��D�N�p�r%�bX�����Kı<}��.�k.8L�a��K��`j'���߶��bX�'����iȖ%�bw�ߦӑ,K���ND�,K�����%5urMK��Y��Kı;���ӑ,K�﻿M�"X�%��w�6��bX�'����ND�,K��x�MfSd̴*�l���A�qYBӵ����'�ү��f���6�RUM�����O�,K�����6��bX�'}�p�r%�bX����l?����5Ĳ�}�p�Bd&Bd,�!�L�T�^��̛ND�,K��m9� ~H��$�����&��	����m	�.�ܨVB�	������`�M&UV�&fND�,K�}ͧ"X�%��w�6��c��D�Ow=�v��bX�'����iȖ%�b_���kDup��n�fӑ,K���{�ӑ,K����]�"X�%��{�ND�,� 	r%Ͻ�fӑ,K���<�x�ɭd�,.��ND�,K�g}v��bX�'��m9ı,O�����r%�bX���p�r%�b]��???���u$0D��Ģۛ<u���f��s�	�&��cb��v�����kYv��bX�'��m9ı,O�����r%�bX���p�r%�bX��;��Kı:}ݔ�.d�.\p���iȖ%�b}���fӑ,K���{�ӑ,K����]�"X�%��{�ND�,K�{�S^�d�Ѭ�R�Y�fm9ı,O���m9ı,N����r%�bX�w���K���ݝ���!2!=3j��UV�j�։u�ӑ,K��ﵴ�Kı>�}�iȖ%�b}���fӑ,K���{�ӑ,K��ӻ=	\ֳ.WVfk5��Kı>�}�iȖ%�b}���fӑ,K���{�ӑ,K����]�"X�%�<}��3l ��ӯ�v�ΚHMIt$`p]W l �>���@��Z�u�!�\̶.�6^����U�i��s�8��Ń��:ڍ�Ƅӹ�nɈ�h���8����y���֍ۅ0Z��Xs�{q7c�ه`�З�cc!us]8;tOBdK��k���j.Z���U������L�øD�z���+\�Ю۝�w^�����.�8X)G+ �o1g������,O<t�g;[�b�y��6{q�q�kU�'�,K�����fӑ,K���{�ӑ,K����]�"X�%��{�ND�,K����+���d�.����Kı?w���Kı;���m9ı,O��p�r%�bX�k�kٴ�O򂚩��'�r:�ƮMk%�au�0�r%�bX��}���"X�%��{�ND�,K�{��m9ı,O���m9ı,O�g��3)�����f���bX�'��m9ı,O���ٴ�Kı?w���Kı=���m9ı,N���z�2a�.8L�a��Kı>׻�fӑ,K���{�ӑ,K���ﵴ�Kı>�}�iȖ%�b{�x�9�,ֳZ��m�mZ�z����9pQ��8'd��ε�%s&E9��e��������x�,O���m9ı,Ok��[ND�,K���6��bX�'��u��r%��	�����R�f��Z��9�p�Bq,K����ӐҊq�"j�@(VHA"�,�@�%!�	[�O"�y"X����iȖ%�b~��׳iȖ%�b~��iȟ��Os���~?����c��p����߬�%�bw����Kı>׻�fӑ,K���{�ӑ,K���ﵴ�Kı=��麗Y5����ə�ӑ,K��^ND�,K�}�ND�,K�g}v��bX�'���6��bX�%��=5tWWpɖkZ��r%�bX���p�r%�bX����v��X�%��g��ӑ,K��w'j�p��L��^J^��M�C>�X�*�J�{)�WIɫ`ݰ���]�ۏ'T疎(��쫮냕�n��{���7��bw=�v��bX�'����9ı,O���ٴ�Kı?w���Kı?}��̦�Ln��e�r%�bX�w;��Kı>׻�fӑ,K���{�ӑ,K����]�"(:���'�{d?�s&s5&k2�9ı,N����ͧ"X�%�����"X�7�6JOթ#p��h�u��ȁ��>x@ ����6 ����?�"�*H%�^~#6���։YF��Y�#A0���vq��~W�UP?(��v*@�ʻU�(=:� / �C� TO��'�f�v��bX�'����r%�bX������t�9T9�SUp�Bd&Bd/����Kı=�w�iȖ%�b}��ӑ,K��^ND�,K��N�MI$�3(sJ�p��L��[�w�iȖ%�b}��ӑ,K��^ND�,K�}�ND�,K������Fp�R��l��+�n=v���٣u˸�u.�𐝣4�qX����h�n��k.ӑ,K����]�"X�%����{6��bX�'���6��bX�'����9ı,Ok�;�Xj�&fk2\˴�Kı>׻�fӑ,K���{�ӑ,K����]�"X�%��s��ND�,K����+���d�3Z��r%�bX���p�r%�bX��;��Kı>�w�iȖ%����;W�&Bd&B�ѩj34j��.a��Kı=�w�iȖ%�b}��ӑ,K��_{^ͧ"X��y, Sc���r%�9��r%�bX�����fSY&7Zֲ�9ı,O����r%�bX�k�kٴ�Kı?w���Kı;�w�iȖ%�b{��p���l��S͔n�Z:���a�e6]ŶyH84l����1y��+�/R��f�.ӑ,K��_{^ͧ"X�%�����"X�%�߳��ND�,K!w+5�.�	��쬖��t�L��Z�k3iȖ%�b~��i�*�Q5��s��iȖ%�bw����Kı>��׳iȖ%�b_I;�e˚�MMSZ�.��r%�bX��;��Kı>�w�iȖ%�b}���fӑ,K���{�ӑ,K��^���+��e����f��9ı,O����r%�bX�k�kٴ�Kı?w���Kı;�w�iȖ%�b{])�M�W	33Y��]�"X�%������ND�,K�}�ND�,K�g}v��bX�'����9ı,LS���%#bVF�$+H�#'�:wO�?�u�,%-��m��zn���ut���� C��� ?���  ��v��׶i�:S�]�mn�cn�3��S� �������#ڧ\��bj�F+X{9�:�iܜۭ'`x6�4ԫ�s�^3�ƛ�k��굫9v]��jͱʒ>��+JݮM��K��%�m�Fu����b����k���Ꚗ�+3��~{���۾��2�A*�ݔ�ڦ��[&7=GrڹN���piz���鸤�����ˆMYsY�O�X�%�����6��bX�'~���9ı,O����r%�bX�k�kٴ�Kı;��h<K�\��X]e�6��bX�'~���9ı,O����r%�bX�k�kٴ�Kı?w���Kı?}��̦:�f7Zֲ�9ı,O����r%�bX�k�kٴ�Kı?w���Kı;�w�iȖ%�bt�vCԹ�2\�&5�v��bX�'����m9ı,O���m9ı,N���m9ı,O����r%�bX���wS�e r9����\!2!2ٻ�pr%�bX�����r%�bX�w;��Kı>��׳iȖ%�b~�}�hC����K<t�9�T��9[��np�<V���R���Q9��챴�Kı;�w��Kı>�w�iȖ%�b}���f��)?D�K�]�{��p��L��Y>{+��h�D�Y��6��bX�'����9�<V"�Bl��"r%��w���ND�,K����"X�%!gr��\!y%�I	��:���)t
���uN�p��L��Y9��\.��%�����"X�%�߻�M�"X�%��s��ND�,K���֥up���sY�ND�,��}����ӑ,K��}���Kı>�w�iȖ%�b}���fӑ,K���jZ�r�$�'4���	��	���{6��bX�'����9ı,O�����r%�bX���p�r%�bX�w:o�v��AK�Wn�v��{9t'2�3��q���N�m`ܬ���v��:#p��m9ı,O����r%�bX�k�kٴ�Kı?w���T'蚉b�so���	��	��n��t���̆5�v��bX�'����m9���j%�����m9ı,Ow���ND�,K��}v����:���'��=�Ī@�((s53Up�Bd&Bd.��iȖ%�bw���iȖ8*	�)�2'}���r%�bX������rBd&Bd'�fm:u5$��̡�+��,K?��{����r%�bX��{��9ı,O�����r%�`
�!w}���	��	��}�xL�*�Iuf�d�r%�bX�w;��Kı>��׳iȖ%�b~��iȖ%�d,�^��&Bd&B��w��K*���Z[nOS�C�4�[]22��h�v�a؝�S^KIi2t��NT�1)=ߩ�,K�����iȖ%�b~��iȖ%�bw���iȖ%�b}��ӑ)	��	�5h9@��n�����\.X�%�����!� uQ,Ow���ND�,K��]�"X�%����ڸ\!2!2�V���.�IbsO0�r%�bX�����r%�bX�w;��Kı>��׳iȖ%�b~��iȖ%�b~�;�	�Lu2�֮�m9ı,O����r%�bX�k�kٴ�Kı?w���K��y	 HBA �HE#�BI $$d D����N��6��bX�'ǽ���3&�2L�e�r%�bX�k�kٴ�Kı?w���Kı;�w��KĲr�]��	��	��ݷ3#�L)�M|}�tg��ɮ��؜ݷ;���NvݴjK5)l�8#N�n�;[XYk���7��������6��bX�'~��6��bX�'����9ı,O�����r%�d&BzfӧSRI-L�Ҹ\!2���ߦӑ,K����]�"X�%������ND�,K�}�ND�!2gL4L�H��ꋅ�ı>�w�iȖ%�b}���fӑ,K���{�ӑ,K���ߦӑ,K��HwܸMC.Hk3Y�s.ӑ,K��_{^ͧ"X�%�����"X�%�߻�M�"X��f�w�����	��	��o����MԔ6:�fӑ,K���{�ӑ,K���ߦӑ,K����]�"X�%����ڸ\!2!2}�\~��m�UUUK��]�)�ƞN�7�$(�5��m h � 6�  �Y�xmv���]�1��m;V�<�u��u��[r�C��=cP]v�^9���O/�ϭ���
踁����x�F�Բ�d5ʜ�^x�ku�N���v�{��@`�<f��CP��v���^���Ys����g�]��.w)�Gj�ڂ�H�<�Nd}��Ȣ=f��+*���rԙ�r���gb�p�@&]�	��5�'c�Ou"\�	%��:��.��	�����\�bX�'����9ı,O�����r%�bX���p�r%�bX�����fSe��]j�&ӑ,K����]�"X�%������ND�,K�}�ND�,K�w~�ND�,K�{.�kR�d��"���.�	���ݝͧ"X�%�����"X�%�߻�M�"X�%��s��ND�,K�f&�B������U��	��	�����"X�%�߻�M�"X�%��s��ND�,K�}�{6��bX�%4��N�MI$�3(sJ�p��L��Y���iȖ%�b}��ӑ,K��^ND�,K�}�ND�,K�����n��*��-ٺ�t���\ܚ�כ�:��a��甄���՝��]]���W2m9ı,O����r%�bX�k�׳iȖ%�b~��a�A'�!2!{6�\.�	��څ��He�fk5.e�r%�bX�k�׳i�D8+s`~U�ț�bk��6��bX�'{��m9ı,O����r#!2!>�ՠ�iRP�S5W�%�b~�ͧ"X�%�﻿M�"X�
�Q5��]�"X�%��{_ٴ�Kı=�WW$Ԛ.��m9ı,O}��m9ı,O����r%�bX�k�׳iȖ%�b~�ͧ"X�%�����&e1�[��֮�m9ı,O����r%�bX�k�׳iȖ%�b~�ͧ"X�%�﻿M�7���{���??�
���fU��W���[V4����u�4�.��y9��Y�4��c��ۣ�f�5���f�.ӑ,K��^ND�,K�}�m9ı,O}��l8��� ����V(@�wM�I�h!td�.�sY�A$N}��n'�K���ߦӑ,K����]�"X�)��;��p�Bd&Bd&���N�f�&��h�Y��Kı=�w��Kı>�w�iȖ>0� D����C@�CD�Mk}׳iȖ%�����\!2!2g�n�*fh�&��&�&ӑ,K����]�"X�%��{��m9ı,O���m9�b^�I�{�p�Bd&Bd/j����.Hk3Y�s.ӑ,K���{6��bX�'���6��bX�'����r%�bX�w;��Kı/�u5m��.&
UWN;ni�k����5g�u��	�
�.�m�0���lݫ0�~ND�,K�}�ND�,K����9ı,O����r%�bX�5��[ND�,K�d�x��䆵!u�0�r%�bX��w�iȖ%�b}��ӑ,K��w��r%�bX���p�r%�bX����̦:�sP��Yv��bX�'����9ı,N��}��"X�5Q>����"X�%����;��!2!}�;B֥T�5T*Fk2�9ı,N��}��"X�%�����"X�%��g}v��bXB#!����bP�EJ�P� �"k���.ӑ,K��g��>uP'*��*]T�.�	������Kı;���iȖ%�b}��ӑ,K��w��r%�bX��9w��3-
��%v^m��È+�l�yzW#bɸ�nk���Zk�]r�#���"X�%��w~�ND�,K��}v��bX�'M{����	�&�X�B���W�&Bd&B���r�f��h��W2m9ı,O����r%�bX��}��"X�%�����"X�%�߳޻ND�,K�!�r���fk5.e�r%�bX��}��"X�%�����"X�%�߳޻ND�,K��}v��bX�%���Itɬ&d�[I��m9ı,O���m9ı,N����r%�bX�w;��KĽ
$,U���.�	���G���䆵!u�0�r%�bX��=��Kı>�w�iȖ%�b|k�����bX�'���6��bX�'�:�`?��wt1�6 P�© �J��)(�,0�1B#"iX�Q0k1ћ�L1rb4H��'D`�q"��ā��4o9�h*����&����.�c������"`�Җ����>"	� ��!C��Xw�N��~~�{���    m�      �L�G5m�[rM6`b6��Z�dN��5�tH� �kik�Q�n�Ret9��@)oe���F�B��Z����t�J�@*�����H�����      �&�   䲀       ��     �                �x�      �   S�+n�P�D��k�v��$��}���ko;nӥ%�/	^���6�;kc:$9�ME�l:1z�j�J��[V�;FyM��`������]	h�tT�RJ<쳝-U���Ik�PJn'�Z�n�@ӑ-�f����0���4���p$��F�/l�v0,�܈óUP�S26y6ta#��'l��j�t��7F���E��[R�z=��gai3�X�m��m�V��0�s�<�5p���c��.����d4z��]I��$�X9|���]��`HN(����(q�������L���s�`�`���q+�F����(W<��՗��x7mۓ��ݶH�vxݥ�T�Bn�.�㎸�@�D�BPM�5�n�L��2ؓ�.N��"�4�D�m�ˡ�j�9*���B����9uT�X��.�v=��2Q*h@8�@���:$dwT�Cl�n8���d���ׇ,�����]�f۰m����lr7e��,37��Z��Y{��PnN�mhv-��6Ne��a��u��%UI��q���[�<���F�AlG<�\�q�tr�ʭP1p�k-6��m]t�#�
\+v�n���&.W��|��jM���a�$�|�.o;�8׶4R��ܲ��g�K�L�\ ��V���P:B�lo�#��u���s��p�-y����_t�v��n�3Yz������*���砉U�誙� ��em�ڮV�]D6�$��NS ڦ��0��3a���]�������
qWi�'�!�@ؠ08��C���fkZ�h�Z���^��k$�2�`E����� H ��l��F6��bI]�K�n M2'&�1�M�Î.��L��<����[ny�h�\��$��YZ_$��Y��q� r���ɗ1��J�]kj��e���bGϙ�çv�&�l��,�#jj��`U��['n8.܇a0v�Ͼ��à���:�nW��l��a'Q�w~�����tD�D��b;t�s���v�vwn�w<q��]I[�q]�p޻Qט'p��w�Kı=����r%�bX��}��"X�%�����"X�%�߳޻N�	������*�I��R*j��Ȗ%�b|k�����bX�'���6��bX�'~�z�9ı,O����.�	���2Ч]T
d��ʗU;ND�,K�}�ND�,K�g�v��bX�'����9ı,O�{��ӑ,Kħ�{�2�\3V��%�ND�,K�g�v��bX�'����9ı,O�{��ӑ,K���o��	��	��z�&f���哚˴�Kı>�w�iȖ%�b|k�����bX�'���6��bX�'{[��p��L��O1��;29�n����ś:�q��"�c!�=�0��������NOE�4�(�����{��2|k�����bX�'���6��bX�'~�z�?���5ı;����r%��L��W���4��i������ı?w���8D�K�g�v��bX�'}���r%�bX��}���/DD�RBd/eK�n]��Q��Kı=����ND�,K��}v��bX�'ƾ����Kı?w���Kı?{;�	�Ls,�B�Z�]�"X�+Q;����9ı,N�������bX�'���6��bX/BPI2��p�Bd&Bd.�мԬ֦�2L�e�r%�bX����ӑ,K���{�ӑ,K�����ӑ,K����]�"X�%�����3�nٶn�[l���X�g�L�{98m��X�<���6�˭�<��9ı,O���m9ı,O��z�9ı,O����r%�bX����ӑ,Kħ�{�.f���M]��"X�%����]�"X�%��{�M�"X�%���m9ı,O���\.��D�RBd/N�s$��:NU՚�e�r%�bX����6��bX�'ƾ����Km@�RN�+�ҕb�t$Z�҅��q9[��m9ı,O����r%�bX����������d�d�r%�bX����ӑ,K���{�ӑ,K�����ӑ,K���ߦӑ	��	��(�U7ChuSp�%�bX���p�r%�bX�}���r%�bX�����r%�bX����ӛ�oq���?��9�o�X���z�Sf-U����7l2a�:�˹�����n��&�ʺ�7.�L�rMR�\!2!2{[���Kı;�w��Kı>5������Q,K��p�r%�bX�z��H�j���"s34�L��L����6��bX�'����m9ı,O��m9ı,N����r%�bX�}�vC�њ��k&fd�r%�bX��w��ӑ,K�����ӑ,K����]�"X�%�߻�M�"X�%��hS��2PP�f���p��L������ӑ,K����]�"X�%�~��9%������,H�h�i@�aH��S+��z���524����������^�2sflgrՁ��DF~G�S����
U^m���:� ۯ�V�m�.�5��c=���U�6��B��p�f���<�� ��s <ʀy�HWZЗ�L	#��s�ށ��T�j@;ݩ =���Vhn��q��빠{zS@�zS@�}[�/�������&93@������������~�w4����E���U�^i �v��9̀|�*����w����h��ۭ�d�K�zy���jo���|� m[ l ��  �`�j��V�-gJ��4�HM+fN�gU�#� �EvCD��6��b���"�]+r�����/k��<�nt�
8�b4�݊Y6��g��`�I�4��F�����l�-��h��\E鷬4qHCt�rS�'�������gF�ba���`]^�w��n�%`��뷖��݇v�)��-��AŞ�l�*�i�S+ٕ㣞�*�Ē��ߛ�?^����?��3����mS?��� ��o@�z�hޔ�;ޔ�;�V�/.�$���ƞ&�hޔ�;ޔ�;����]����nE1<MHh�V{9�63�j�b(I���`n�>�c�F��G��o@�z�hޔ�;��h�RO�d�8�jA*��wm��ۄ���ȧW���s��,�����qF�dlp$R7�~�w4�)�w���=]l���2��P1�NI�Vs���(U
(��;���������s@��|�H�y"#16�,�=�`|��Uf�ۛj�������ɼ2�y)'��Z���@�z�hzS@�_U�~�S:��8�Nff��grՁ��,ܽ8vs]���d�?.��Ҥɉ�MĤm� �-�ݝ�Л��Xڭ�1���J��9�F�C�X�����Jh��W[&�����?*ajm6�S��Ԇ���n��݀|�*�j@�]�k�1�$r
E�z��4׮���ĒN"*��XXvs�}Ջe�c� �I4׮�ץ4��Z��&�}e̸$�l11ɚ�)�w���=V�4׮������}-�E�0R�]��u[�5�����y0�q� ������޻Qט�@gg5�<̪�9��[	Dq��V�s+xg�&G�I��9��ɠ~�w4zS@�_U�~�S:� x�!y��� ��T{R��n�Wv��RuRɥM�.S���b!BI���`gg5�<̪��B�B�� ������L��77$�{	�&�n8�x���;ޔ�=V�4ץ4_U�}癞.��S���n-�����R��U�he1�m&ہ���u�I���܌k�2$n�����4ץ4_U�w�)��\��H�0�3@����j@9�{� �vh�\˂M@����k���4U�M��M�v�0�@��*�36��Ԁz�݀|��s��=��o�((�	$4U�M� ���ڐ���n��UN�5lRɏ�W�n�e�1� 	 � @   m�[�����{F�R�=�uF���Rƺ��ڦ�)�x���ꛓ�*]�xx�����]�C0=u9�q�>,��V�(90�r���=w�m�.l��+�Y0gӓ6� �tX�&����	�r��s���ٽ�vB�c$����.m��X�ݤ��l�%��{���w}���?M|}�t+�ݭ����tiF�O'��nѩ,�sg�d$�Ŏ7<N2	�䞁������h�Jh�l���Y�Ƈ2$��������;ޔ�=V�4׮��bG��}�m4�'�qh��Z���e@9��K7Y&A�#q�3@�[d�:���-}V�׮�{�|���s	���$�@�P�n�2��w`Ny����V
UWk�-\��p��3;ۅ�v�0��bwl�`�y��v��ۇ5_ ��}����fh��T��L$�����qhޔۛ�g/3�|���\�n�*���j�̞㽈P����)�ɑ�8c�I��}&�}빠Z���Қ��,�Ȑӌ�m9Ua��7��ݜ�`gݬ,�fUX~�[�D�IcOs4_U�_zS@�[d�/�w4y�� �2A'@�[8�f���v;R����:���[�</Jmv2��f&�MIx�qhޔ�=j���P�n =Es�]�n��F�Y��֮�y� \���M ���[I���$�@����w���s�w*�@Y��WK$ @"�hed�х#$ ���&�TVt1(}u�;�aiMDI_:5]��A.��h�O��z�?H� �`�1 �4|B����`@yKьxU�~��$m�3X�q0� ��U��X����H��� �� ��]l!4�	t��sdH�E�0(h�Dx$3+�f����"F$#���#
K�Yt���j% ����VGaib$!%��Ў�;�! �Ӵ�+z_��O� �ߎ"q@:�� W�7�W�?�j�A��,7��yٹ'/~�f��̸$�l11�h��@�����ɠ_zS@�o��%�����R�Wv �� ���aP�kc�*�J�lK��f7gӀ�zz^Ę��o'8�k2�K��r�;Zz�4۟T���ɠ_zS@��_y��gƁ��縲G"CN2	����4_U�_zS@�[d��{lD�%YyW��{R �� �w`�S@�����i�#OCR��4�fUX�kIEB�$З	D��tD��E�Ex�����7$��C��!�aCp�=V�4�Jh���}�M�<��{Uhh��QĩG+�8�i���A�e�q뙰�p����u�oa��?#i#ȅ"iI$��gƁoj@v�֮�����.��`Uᙤ{R �� �w`�� �o��$����_zS@�U݀>�T{R�awGV�囚V~�� �w`�� ^Ԁ>�M�Z�H�Hi�&Ӓh޻����j@=j��.�~�T�twv�k��ɬ8�Y,�Rt���u�Mz� �� m�  wM��j�j���R�v#�]�Ei�/a+ju1C;���l\sr��;���u�x^��Z��7b�H��.�##`+^Ic�4Ii'#����_(Uk��Ict�땣p�k�ݭ�7�Ym�pn�%6s�\���b�S�Bu�	�7]��tz�λ �֧�S-l����+˦6L�@��v�]������f�0lk������B�2�o^���}i�)5hG�����mx�3���3*�DD%���Vyb���i�#OCR��4U���ϻ������n�n�S5H���h���4�]���hޔ���I�D)JI&�}빠.spݩ ��� ���h�˭��xf�@9��Ԁz�݀>�w�o�����C��`�W��8(�ܚU�v���rn�9Ɂ��qf������N���n-�Қ��&�}��y��;��;������1�$����ʫ����!bI$�]�rՁ�Oq�ޔ�?u�qd�D��di�4��j�̞�aD&��ZX{�U`��f'��bX������hޔ�=V�4�]� �V+Si���<M�� }ڐZ���ʀ.sp6�~����{Y��r��9ۺ���ѓ�;6dؓ���	�=�1�7;x��̘9o7m̳3H�]��e@9������I�D)JI&�}빠.spݩ ��� ����w�[Xc����Vd���v��RJ�!BJg�m�@��w4V��A��
x�n+>�a`|�2��ϻ��5BP�k5��K
|�dh���C@�[d�/�w4��hޔ�;޸�k��q&�nٶo\�Ƚ�����#<��6rq]s�2�����G�N2		�h޻�˩ }ڐ�M���v�+r�e��r��+����Cf�+K ��*������b�Lm�#OX9�� r� }̨�� Z)rı9�6��4�I�_z�h��ܐ8��A0z�f��f��Π�c��L�Bh޻��Ԁ>�H � ����*�ޖ[*�J�{)���s�p��iq�R�χo#����R섘6�3&&�58I3@��M�j@��� ��P�闷{yuxfi {� �l�ʀ>e4ޱ,8�&F���$��֒�ϳ-Y��v��72��9�d�j�j�&f����a����V�kK;ڦ�^����;2<P��,i�Nf��Ԁ=ڐ�6 �e@
��]������U����{EHc����*�ڋ,��E.ـ�  �.� m�[x�J�3i��b�f�^{b�'E��\�]zɂ�l�QPUF�m�Ѿ������-S�;�+��<T��q��7/2ue�����@a����q����r�h ��L�K��\n�m�:�&���5yz��ݞ@��9�8c��$n���R^�`3�B��]��U;�� �R�mmd1���b7ţU��6rܼ\;=	���)�*T�a����{� � |���Hnա,Nx��7 �i4� |�@�H�)�vVmm��xnn� |���Hݩ R�d��'-�2YD�5J��=�ސ��� <��s*����3K�˫�3H�Ԁ)��ʀ_l��}�ų�j6�R<x��0�h�m��nÍ;e�@�� ��>���6�e{8;Zkkr��2�wt�)��ʀ>u4�Jh�-oq�I�m�A!HM$�ﻳu@�@�C{�߳�rO�v|h�h~���EBƞ&�@u �Rָ��2�u�f7.f]K�NXMQa�
"�/K ���@����/YM ���,Nx�2ɚ,;�V��[��.���������wT��ɂq�ԉF���Bm����j�<'h�9���87=��b�\�l���d�A$�drM��s@�e4�Jh�f����q4�!�D���� {� ˰�*��(wr�X�N��m�vg�瘼Ĉ��P�8�������=��rOޱ,8�&F���$��m����3+%��zXa�3jU4��f��{� }̨��ݩ l�*��M'E0kq)m@Ȓ��iK��Ͳj�M��m]`�9gd�sMY�J6��<M��-����4�f�}빠��cmF���Ԇ�}�H ���ʀ+�?��ꪪ���챴�)9�c�v��V}�j���h�U���F�1�$�L�w`w�{Pu g7O�?U~�4P���HP�T �� �L��L&�r�T,$B��ID%��;�`o�ljr�!�f�{w�Pu g7 v �eh�QdM6F�JF�Ra��C�l��>�Du<��
��vy����9k��=��lm���^i {9� ���* ��@��Ê����ȴ޳@�۹�Z�������=��7��,M6�2 NM������h�U�����; �Fб��9�y�$�k5��������J�w��/$|&6�j<M8�Ϫ��3-ޕ=����I���}��}w$��*���*�� ������1EWB(���Q_���*����*��ADU�DU�DU�"����EU��"�DQ^((���Q_��*��DU�"����EU��EW��"����
�2����2Pb�����?���������\}$����� �    #Ŧ���Z�X�\6�n�>�{]� v<uU�UUb�����iJ�6�(w qi�B�g�)J��W����W���JR��-�CӜ�WM8ڕ�[g3^�qj���Gi^ ����k�J��U_x!EHl $F��&�"�OSjM26I�4x��i�BR�@2 4h4h�� �~=UJi� � @# �2���T&�R�� � #  �#L����R�0 # � &  D�@�SJ?T�P���M�z�hѠ��4�^ͦ� �@��᳚@�!h>LP���` ��*�#�>���?��9PB�d�}x��_����?rF��dW�o���?L�;�g�k���N��_̖דJƒ� BkwY��:�s���D�P���
�!G��,Wį�N���&`���A
�m��h�O�n���/lk�I�;�c�d����V�]ӑ�𑄺vL'�C=��%[VS�"3=8Ċ^���uE��-MDل�V�q����F�� B�$�HD��iD�
��B�D�(Y ;݉�j�
S�
I0�6����=�b�j�)^V��=KS �$���@��������k�T�T!z|�b�r�TZ�(��
�e1��B�F#D$ɓM�C����je����4M�^N_��^aP��b]ZV�G+u������JxB� B�1���(�0@�F��G2�P�bI1( �J�k���r�!أksڮT �P�M�^T�	 ڀH���B�b���L��x�v»�\��:ͼ��c���D�5#b�$�!X�#@F1"F�Q� F��
�IH�B�0$	$aRPD�
�H�@�5
(T)7�р��e
�*�8#���1�B�(�(m%8n�4�`0)0ʮ��/�u���C��'�}�:4@�KF�y�6�� �c5�&X�F�Zs��9�s                                                             ?�=                                           �Z�m�It�Z�Ͷ mQ$W.��w�j�
�5jH���jH- -�mv�x�m�m��m��G[;Ci�9E��s�                                 ��                                                                             =�       |﫷���m�[@$ �^�kCm��[�� նݶ�e�ȓm�;e�v�E�G��՚IW�m-��-�j��N����@�[rN�M/Yv�YH� Uk���l�`H�v�@%�n��>�z8 �L�k�� �������ŶM���m�@�Aj�[��u��$]6�q$��l�Gh�$^����I�m�-��l��x	�񞧯^�-��mRlsm�Hk͛l�c ȶ��[\ ���Y0 m�E�mmƺ�� �P�We�:^�kyo��qj�M^]*M�e��p�$�(8RV b���VŖa�	DB���26ն��#XA2�PlA��P���B�d@���6�m�f���bI�-K��!����� )���n��)��WXۖqp�v흮l>�c��Dn�0<RH��!cs�h B���! 7w]����O?�\3	$ 1����Ow���Ȱ.� A��B! ���rD>�m��~�6��b�D*uL)�/QNpRĂ�EP�gt�� ���ʚS�H��Z!�z�� GBЧP؋�i� �������AF0�d��x&��v
�� WP
1��@           6�        td���z�Z:(�yδ�      6�              m�.��]in�)5��3�d3µ
з(bF�jY�����P��A�(�՚�[`�І��&+�\�Y�ڲ�':A�KN��Rd������@B�(���e�#�?�|}�>� 6� �v�:l�  �N�7+j�!a�)�Ac��*(���Gގ����~�p]���ʬ��7��.���ws�:�ϖ�I��Z(1e�r~�"&��S��w}�*�χ1���Ӹw|_�ueZ*��2�︆����챘\�_q�K�>s�o�j��p,p�����ws�;߻���iWsꬼ�7��V�ޮJ�"*L
B#;ӯ�s�p����N��k��7�3�����_yUUUUUP:6��M�   ٤�׎�[|H^i-sm8\�
��YqiH�p����窲��v[]��3.����WbJ���uH�t�k5������f�͍c�9�=��vҮ��Yy���ҪH��!D�� �������"b=�N�����޶�z�{����*�U��P(�<@��J��Ue�!��:�>����N�_s�j��r�!�Y8q-��a�UKz��C,wǈ��i.�����   �H�&�   �u�3$��;T�[��� HP4R)R*���P�;�����x�$���瞝;���eZ* �)�J���17ZǼw\F {��vҮ��Yy�}�nr�o�Օh����Yޝ]Űizf&;�<4�ؘc�'�{�E�J���e�D�F���*��X�KfZ $X3&��F���膅P�hX.�Q����u[�us��{��s|�s��r�V����o���owޣy�umv�X�9��311/���KI|���h�\#alt�[_�y����ǈ��iWsꬼľ@^�I$�H  ?�ٽz�z�    X��U��޹5�N+d�Q[��eZ*�)*H��v�����3{�>�X@=���V�f2��Y�f��3M��2f"�Q[�䪒%$�Q������.��݉����8 �P7�j�PǞs�\΄���Ù����L����n���舋�ߗĪ�%$DJ*LA6��d�߽y�n�-ۧ3}�m�|4�(\ҍ>�y8��$>�u���o���؈���/�������5X�t�5�j���xA ������Ǡ�S<��ʃ�ߏ7;�m�0{���s5ZvÙ�`-��y�����=Ϋ��*��I%PM"6D��;u�{�0�>��̨�0o���s;w_>|�3�TD�w��ɉ/,w{RI$�  9��t    	�:��j��ګm�-`*ڠ�0XR{Z�Uj�q혉�>f:�q3.���u熗;�U}�q�☺�=㻱�k�ؐ������DU�/2&������mEw���s����q��E�َ�2V]�^߉U$JI*�*�tD7w\���M��V]�:�χ1�x8.�U��C/1u��UI�B(�R�Aյ��a�ؘ����<�L���?N��+�^;����*�U��A@�����U��C/1V����sS��/���ΐ�y	�D&B!�".$sn�
	�:����                    ͛��d�Ɖl�kJ]WM֝@                       ���k%��e��R�����6��i��Ɨ3��Zѷu���v�k����)4�l��`L�Յ��\�Ih�b�&L$�-(�Td�J�]]SM��Ǜց���"������  � t��[&�   ��݈�io%�a��b=z-6I%TDI!X{.��[σ~�+v�_ϔյ��c��[��/x2����I$�B(��$RT2�o;��0!�?w��a�����xq~��N�|>YV���U5m��s ��!ڈ��w]ݴ6������=��V�V�**����b�in��b���nb".���ο;��T\�A-JĜ�����y����e����u��Ky>I$�  -��&� >`�  :ݥ�gm��Z�ős���`�{YV��4�Q�!ǹ
[�j�c��<AwG7ž�=ow޿S�YV��!�,E��]��3L�^��,S--��a�B�u�3�s�j���#�{α��!�J��Ue�DH���1�t{,e��{.w�_�c�o�ڠ�0\-F^�_r~s��M[C,wǝ3Vx2��Ϻ��YqB���o���65��c0��b�in��b�6�$�H  ��wK�   ۥB]��l��]&֒��w[��`^��%M[C,wǋ�W����W��ow�{����|��mPWJ�HDg+=��30.&&S���2��ަ��q{�t��*�U����s|;��9e:�c�\k��fM�Rr���+Ŭ�DВ�S
/ �!3x�`� B
F H	#H�`���
'��ӫ�L�@�#pߑ�!�x*�ۅ��GC�_UDUL�UT8��EQ/C�P�o�-h�Z:zΩ
ǂ��y{�֏��CBD��V�~y˪���u����qb���"����rgf����!�x*wn�r-���T<f��֎ţ�@�n�;������  �me�l    Fĕ8km�e�l9��n���󻼇�D�����T�5#�X�T8�^鵣�h�Qݕc�P�8���h�]іC�H�c5��umPUm�Hb��vh�٤^&�����O�m(�Ȭ~�襣�h�Q�:�Y�i'�����֏�L�o�EUV\����uɛ���wg�x-�2�x)6��{�Z9���o�x*
�]��*�TU��7y٭���2������pT8�/t���t(�ʈ����4�����vk�;4���ŵAU�J�*��x)
��ۅ��GB�7ļCپ��k��^�:ϪG��������^�   K�e�`   ͎�`��u]��E�[ّq�uT\�A%C�vk�;4̾�n�V<;��Z<���d<�S^��ɼ��3�L���ʴT�q�JMQ/C�P�o�-iM
ţ���=��#�X�T8�.�mh�Z:weDC�75Ɍ׾}Օh�ܸ��o;5ȴt.��!�x*wn�r	��F���s�z*
��tZ�شt(�_-�
�����)5ɛ���j�g�-h�Z:weDC�X�T8��-h�Z-e��7z)
����*�j�E3RB���-h�Z:��%��,z+�>�-h�Z:u�T�c�P⼽�kG����(�$�@�*��C�|����                   ں���:�]�m��$�Y�                       �<��k��[XT���6[�K!ZjVĲTT��UYDL��崄 �aG%��L��b�A��.*L2�7-Ύ�l��n99.H�Ukz�r��<8�Qйox���݀  �%:޷    Im�2KfE���k�r�p>֥����YXɉ*��!�z*og�x-�2�x)
��ۅ��GB�7ļf�}�-�
����n�[�٦(��R<<�0z+]�t���t(
ǂ��vqkG������QS5T�&(���x)
��ۅ��GB�7ļ�F����赣�h�Q�I�L��&3O_���YqiH�kG��У�rx|�FEc�}��Cq�y�k2�C�)|Vמs�'&���f���mPUnR�1�rc
��}�kGb�У�uH�V<+��Z<���Q�V<W��j�   u���   F�����.ٛK��Y�uľw�5M�q0RIPpı%��X�%�B{�p���P�����P�o�-h���3>V�UYpiL$�&nk�P����b�h�Qݵc�P�{8���h�]іC�H�T?Ov�j��r�!��y٢gf��C~��*
��}�kGe�ci�cbi��أ�uH�V<+}�6�x-��l����U��75��\�����Z��Z:�FY#�P��p���h���b�YĽ�$���~�����*5n@�#w�����3/�?$�&n<+��Z<���Q�V<;�zo;5�3]����{?wj������M�Y6    hv$�v�d�m��M��K�.�·�D���um`K�R=~�p���h�^&�����{7��v-
=gT�c�P�ݝU���!\�-7�����3/��ۮIi�IFE����֏��wFYMrc5�{����;4�}_,�EHR� ��^
�����tZ���أژ�)�3��!�TV��x�D� ID�"�h�x��������=�1����M�P�Y���m����rc5�>�ʴUmȶASTZ��t.��!�x*wn�r-���T<&���e�Z�ػ4��x��AU�\E&�3s]+��&֏��GvTD<�C��qkG��л�,����r��uUP  ���`    �]w4�[ea��"�h��I��
b*hŃ�h�^&�����{7��v-
=d���X�T8�wD��᝚fz�ʴUeť"��\���
���֖ذZ;tm��R<{�Z9���o�x*
���ꨊ�Un�V�;5���f_�\��4у�X���mh𦙣�G�mDC�X�!	�����%	Z�*��I!�SD�4C�H�T>��-h�Z:��%�x*�YŭEK�,ML��I�n����Lf��ߖU��.2��7����GvTD<�E!N��h�Z=te��R<��Z9���s�T   :YD�(    ���V�J�ꥲ5K�!&Q���n���AU�$���^�����VqkGB���D����X�T8�w�6�M��z/����75Ɍ׷��dUUf
-f�Z<���d<�6������i
���Z��^���x*
��Vq���3�L�ϕ�h��ZR낱�q[��h�Qݕbԙ����8���h�]іC�H�T?O�յAU�J��Y���3�Lϡ��T<ެ�֎���G���x+
�M/y���j�&ׇ�[ñv}7DUVRQ�m�&nk�����o;GB
G���v�kG"�мM�/C�Pͤ�M50�6!E$�� A�b0�I#������                    %�"���d��͝6�3k&$                       �� k�&���,[��gf��.�Nؐq�4Z�$�Xai��P�%��u*�Di[1�HHXDɔ�7d�uӴ�-��	t��.\�w���Jemz�r8��]���݀ Z�9�    "��2Km�v^�:i�v�K������3MQ�B�У�O�c�P��kG��У�rx+
���֏٦g��?���EVꭖ*ˮ�&��
���{K^1�بZ;��T<���Z:������{!�p����V܄r�4�vk�;4̾�TD<�C��qkG�&ѣ�wF�E#�P��p���h�U�]TETT�0�B���%�x*�Yŭ>I���أ���
ǂ��{������(Mc��b����X�!	���HRTRI
QR�*j�Z<���d<�C���֎E��x��^
����՜Z�н���<�}��   �s,�    lZd�H�&VP�AF�sZ�7��AU�\A.�3s]��W��Z<���d���D=�EC�v|Z��_6��F�E#�P�}UDUH�2�-Fo;4L��3�o��#2hi B��\�����[��6����0�V<+��M�GB�{�*�U�����rf�1������x-�2�x)�5+�n�I�P���!	b�:�*��I%QJUEQkGB�У�OL</�-�/��M�4��}�Ec�y\9=��yٮL��4��mPU�V�
G���v�kG"�мM�/C�P���-h�Z:z�釂��r�����{   $��&�   ���]]6�B兙��b�a)EV\ZR*әɮL��2��m���ǂ���b�v�Z��^�,����׽��o;4L��5~ߖ�V�*ATU�T<ެ�֖���X�x(���c�P��kG��У�*"L������{���EUVe ��f��t/���
G���v�kG'�cA8 �"8�)�KZ���i{b���_�C�P���-l�3�L�ϕ�h��0��&lx*V��mh�Z:weDC�X�T:�5ٓq�7
mRK@ �l�3޻���k��{�j��r� ���Z9���o�x*
��VqkGB�У�OL<�C��tM�GSϏ��   [��    i�%�\�,V��LH�H`,��l�EU�
*Pm����vc5{�=7�����2�x)
��ۅ��GB�7�k��Lf�}�,�EF���f�,�1u�?�x�]�.���N��=y���U��upd������nr��o�=����#�.���U$JI*��J�4Ul���l��N���s����<ss���-�
��p�P�;��2��7��A��.���O'�����|�@   �j��6    f����-��H��6��^�	IQI$)R0
�PU������v3��p����8p��~[T[����]�DJ���8�M���S�Fu��l��ss�~��-�
���Tg/?kK�?,��e��ol���]��y�*�U�����|'~����{�ss���v9�;��2�V�%T�)$�(�(0� ��­��9l���.���N��:2�z�� I	!�!�㪦ꪪ��                   -��l�w��k��ņ��$�                       �����2�pqe�Ԑ�	���Z�6I@�,H�� �XY+,(UU �VU%F1i�ژ�`L!a��e(��̾Y{&��s�i������k7��g���|'~UUUU �݉f�   idݝ�1��J�M�۱���`��R�2|.w��L���;��2��7��O�Z*���EZs|'�߭���>w=]����Ȉ��Æ&W��c)���%T�)$�(� ¤�,���#�.�"g~�����~������Ȫ�̤Z�T��&a{��e3�y�t���#�E�H�ŁPȃ��~L��
z�syslEϹ�۹Wu����wX�\�Ɛyuy�"&b3���� � � �A�|׵YA�A�A�A��\��D��>w��eqq��������  <�N���   ��-Iz��潦���M'3��%.�M��Pwqwn ���&Pwn � �A�o^L�� �A�A��\��������w��Pwuwn �>y��Wx����b�wx�]�������u<��� � � �A�oS(;�8�;�7|���eqq�{z�eq���������b�p��������;�7k��D��5������ �#�B����^w�T�"����u<��� � � �A�<�wuWx����E�%����"�|"DL�}���A�A�A�A��痯fPwn � �A�o^L�� �A�P��$b���~{YA�A�A�A��^{�n�񋻻��*�(�jm��i<Kh���6�O�ϣ/�����?~���^��UUUUUUP�V�:    	1D"[rA�m1�0�2���&r�h���7�ÀŽN���v���A�=ǚB���HR�`�
�����SZ�1�{X�üw�p����8p��~[T[�����l�Cx�dv���m)fDD	�;UD�A
ی\��m:�1X"R�,k2�XГ��^��R{�v�{�æqj䪒%$D��H�����ܟ�{��2�ŽN����2��;���U��.-)l��O}����v3��æwM�e��M$�H  F��ɰ    ����[�n�d�Xܙ�(Zl��ה�/�3
��Ֆ��;��#��l��\���-�
�("�#9x{���Akt���o�,�[���y!IQI$(�	 ��v���A�#��S��{y�r�����^�o�j��r�S����|dbާl�Cx�u�z�;g{l����AE��������/}�l:gt�Y�7��w��I$�I$�I ٸ��    �Iz��'���]�J�K��J�ʴTj�o7�u���ԯw��^�_�����ær��UI�J�!P0�A�;��2���1o�7�3������߶�
���%@�i}�����C��:��oe����3�ߞ�N�W�o�ʴT.��:w��oS�k�3ZǼw^�{��v��6�k-�jfk3�}��߷޿���[�B�	$[]��3.����S�1TN��
��7o�a�<w��t��m���T" �%�" �~����>��f_�ce5�Wю1���v�PP� 
	����,_g��2�oAGt�q�������n�u��O�~P1D�H��vh������<�*�߼Y�I�5�7�niV�5}�.�qy��K.�.��
�Y�d|Ӿ��ӹ�Z6ަH�cab})�DPf|
i�aK�B+�D�X\m��u����_A�^L>���*��}Q�PPG��I%�L�/��Ex�#T��;mK��S�Фq�oߕq�J�#?�bZ��� ��B!=:����1���_�9,lzwt��.��,�P�_xLȝI��b��\�k��Eq~-�ΪS�h�mw����lk�񕘵hz��`���B������i �|b���	�(D�q�~��ۦ�.0V�*�):���RE�2��a�H��n<�� B��+؈�Qdf�lW�-����% ��=s�tA��sT֑�����;�gv���{���~�����_�Ss�M6�IW�I�T��/Dq�7�2��X�{e��>�RN�t�����E>}���K��cc�2��7'��¾����F�I�vV�OZ;I�f���*p@�\rJ��ΰ��&��\xu��E��a~'$3\��,1�UPF��DA�G�� ����� �3�I��}o&U
&��a�@�M����Hi�!"	����H��@Bd�£9Ш�ַC�)%��B<�*u (j�*�a��4���������!e���Ѡƶ �$��G�4� B�6��8�[� 	!g����!��Y���V_���:5!���R��<��}n�_�����X�:�ɕ��r���"p�cQϣ�Y���w�x#Y�2bw��Q[�l�?{@�Q��9iy���>ud�?���>ψ�(!�(���-��G��]�r4v���9x?E�v�0Q��4���U�|B������T��"�A�RVg��V�W ���0��n$�S�Eb�Ĥ�8g�b\���L0���Ј�� ���l�C�s�`�p���̓L��lf5����U�b5I�Pg{2�h�!zKy3�&LTA��;1�ܜ}�.h��Z���֛k1�!)]�V�t%Z�������'~��sؗ�3��
�Q�ԃ9��ܑN$!�� 