BZh91AY&SY�ʣ���_�pp���f� ����ar��*��D���"�B	R�)J ��� ��PP	 )"�B�+Τ     
*R� 
 
D���P�E�J���J
R�U*��
���@�    �T�   PP �h�	�>��E�C��{�� �=@H��  6�T�W-�5�} �R��S��=�=2���Tӈk�=� ��zj�Mv�8����C/{�����4U �H"  �� �b��ǧZ�x0g��,^mP� � :�6s�v�rj���W����,�� }�Nv�B����n��m�mU^}� xyVv�0׌hdc���n :���l�͎!˪�9�T�;��
    ��x��m���^Yq��\�&��z��$�}s5|��t��[�@�'�)��  �,��c�}�J�xoX\YE�7[�w$�
P8=2}'>X�ʌ��A��J�@�   �� ��,��n]���n}��o4�OyN����1�n�Œ�s��(0	>}��g 8��M����%�YNX˳�:ހ�K����W��gu�π@D(   )@f` ���X��8�p�tF7ݩq��.,*��pP}<�s}#|  ��ۣ���8 9��{h{�x�8�t�7� `��g��r=���:x{��vG�@     =@��J���      ��ЙJ��yOD��i����50O��*�  `   �=��CjRJ0     �S)�j�*�F& F� ��	RLI�Ѩڧ���F�M�=5<�ȟ���g�_��z���a�ﾎ���{��
*����@TU]  *���U_��R��������~������(��_��$EW���UU���_���f����1�����)7E�%&2�)Dc�i3y8_��b���'U�wg�kysq��f��J��0NBP�5'�q�J0�F�v���O��y����[���]J��.�0��"�Rs�ƃ���%%*8���Ŵ���H&T�T��U�Z"�B��mb�S�r��Ӥ��*<���2�o�.�9	Bn����( �ŗ5֫g�[�XQ�M�zw.9�$��]�e�N��Y�[��xR�$)R�5+!�EFEC.ꕪ�r��l�"wMb��Ԕ���饋=^���jq_L:0W�[��F'��R���V#�JST�o�J��*��:�T����V.�A�jVx~2=9X�6o�hn��9�D�)J�6����Z�yy�<~���!(![P�e��f�(a$�:2PhsA���%�g�X�hgx�K�ː��Ra�1t��ѸӪXi"i���(��F&�{�i�K���;23Zc;�a��6k��SDf�7��Y�BS0B�Z��g�*�U��B�A)U�b2�/*S	�&��*��H/$H��LM�&�*%:R������G~.�)J��(J��(J��(g��s�|�J�g���V`DI0⢮�J�iW����U�/{5Ld�	ҫ�R�*�!tB@���c�P;����O�(9Mt��;b�V���N�0�:���$Ut�^O/#Suo+�fT�B���Y�lBP�'P�-7z����&�D�����- ��If{C�B$#nC��枝�Ou�:�4fɣ7m{%uJ�--ĥ�y)Hن)��z*L��Q���p-A�kR%RqՉJ����X�lE���VY/�UVyZY��P��iK�^V�7�#޳�#;5�D4%$�����,#�3���Xc����{�AcS��zBP�%	K ��6����5\��sν;OөY��f�"R���Z+ʡl�$BK���6���P��u�c�uF�*��ǅ���e��q�մ3F���:vl1�3FW떭y8�%*Z�18�*= )NU\Ύ����F�n0��BXh��aR/(I�M����2"H�"PTN<L�6�X���^�j�v���X�ë��۫dW��Cafj�s�W!�lG>���R�t���"a
E��U�����	�n��=[�9bBv���Y^���ݴvZ�!K�\��Ѭ��F��H�%�O�ʮ߮ ��t"ڥf��۩\O��h1Pף�*�ؘ�HP���1$Ԑ�-d+�L��G
�\V/N����D���y�J��N�fѰ(�)Q&�1
�T���..�r -��%5>S^�S���Æo�Ǽ6��ttnt��E:�ѳeF��%'I��[����_�'�=�T��Sˬ���X�|���]-T]�����3�����{,7mya>ڕ/��"b� ��&T��Vƽ�"BY7���m�q�g�g������۬N��5�4���	8RI5NB�g����M6;�����ã��BX�7�e�o�� ԗb)b�Y&��J��dx���T+�zms1��z�P��.�7r��˝wjy�̈́%�}�P�5Wq����ۧ��Lm�&��b�$�M���-�w��TDa�ﳇI��R��f��놜<�;2��P��#4��1͚3���;8\7�]�;*��5�r,� �J���2C��'3<#A���m0�̳�F�w�jR%����FH�C!5%+E�Typ���%�D����at8NBR�'p��P�BP�$(@�B�DƲ��W�y��ݹ`�fw��l9^nd�KHfA��V18o��0됕��4Fr����l�V��
&!Z"\��W�X���Ĕ�5l59���(J��a����Xd��&�,��ɣa��N��ӿ6\��w<ؔa�����C�y�.�ͼ:;7�U��ձ���2��j�-��7���7tf9ْRF���D�Z�؞��<乪���ĺ��L�׀S�a�������@M\��W���f�T)"IJ]e�ًi>��.VW�1)i������5d�)\��@��;KQv3A��[�ӫhe�u�$���:�;i�]	��NΝ)O��K�!SMTct�嶈��Il�g�eTX�:�e�/-tL%-R��5�B���IY�W5fR�Oڭ+�qO7!-	]2kPlr�@�rMT^��J��4Jkڕ�)�"��r����H�,��i-2UBʆH00�9ǭu�<���.�{A�$�q^�,��WYx�������X�r�Js�2O%�����.��b������0��\-�;�83���vR*�VR��0���{01]�SY�>��+ SZ���W�;b�^&�ܤז�6�*�^/=�p��b�"����5��F	�D�����������LJ6𻝟T����}�οR���!
]ZǙlS��w���!�5x����I�O�ޢ�w������`X7\�ӭb��l^J���ϳw��}7�(� �u��C�|�,�R����\�X�S���:���(Jѣ��GXԩ��^V���O�U����Ͷ������uW�&(@�Z�)"p�)$P�l�v�N�Ӿ�p�ڍ�:�KN�뮷ܩd�����a6d&�M%�Mڷ��-M^{o�O\����JD�\��VL�P������%��̈́�R���0���N�� t�2�T��U�Rv���:�X��hK�.u�Z�r�F����)�[��Չ��^́�X�'�J3�p���g+[3T�&��+�)y6��WR�ۚ�jP�<��r�[jP��j���)�%e)�j����ǖ�D��J�yic�Q"�)D\ژ�8�iu�֚�\���U�2���1M��4�/u�!8Z(^�d�:ק��u8md(�5`I��`�]$'!7DFBPboVnp'�Z6r:w	�i���P��ٽ;5�6n6aG�o*���R��^ē�HfJ��r�g�u��7����z��x<�磌í�A�]�z�����ĉ/+��Ef��>����b��W)5*&�Ȫ�F�<�n)
E+):�tgg3�ɑ��f����jH����!�L�+�W2���Z��RCDXȨ�r��ݥhT�&7��e�
h�aW&�'u���ZB�K��*��]?\!SII����8f��n�n3{��Ɲ���$5��h4K��%�$��C2Ō� ĳLkX�E�8.9!�jMF�J1�Z�IY�4.�%�a��9��=nw���<ݸ���!�ݹ���v�����N�d%��9HfXA�ե���3 �l!�$�ye�c��˝�N9TG��"cY��� ��
�	�m�ӭ��AP���Er��&��ʬ��U�8e.�9h��n�|���CBԃ!J"e)�M��6UD�UR�;�kNC��%	BQ�BP�$I�d%&Z�,��F�k�㖝��D�]�z��`���sC��E>A���l�a<�:�:��(
�.F���)Y�I��P�*X�IBZ��kZ|�h�Y�}2k5���n`hi(<�$ܔ�<������Eq���&�L��F��"�}g|'"�tof��O7	JS�����T��dI��$I�d	Eúp�:�&��r�) �Jd�I�t�M�u)��b5뎍l�Ɨ�E4��P����Y�c��E����H�I��%���W
x�D)��,#{���1j1l���Z�PX
el(�����an���BD8�|z4nr��"�zs$f���Ն�+D��A��V��%!�bA�����H��<�R�"'�r�� ��4Jn��2��(J����.�\�!�Z�d�)*�"*������a��᎘֜��ބ��1$ᒈ�;u��*�����	BRdm���t�"`	BP��	BP�%	%�k��:ֵ�q�y9�TA4�Y�o۪,���q�ܹo����x���4l͜[��d&�=����n���4BV�dv�'A��s����:;�'!(L������ﺝ���W$)�+��%g������lx�nӱ�%8�ٷ�C�ၭ;㾻��l���Nm	�5���7	c�f�#���15���ܥ
QQ��,Ǟ��g�/���;�=�T�Rbf&&BE�\���r�	�Jq�ko�Pf��:-���4F����=�4N���]=$d� �F[�=�g���4l�ͽ�'[��ޞ�=BP�%	JP�%	�J8�3\|<�`Q4�V)^UcO|����Y�3t��z�<�k�5�u��۩�yc��S��
T�MZ��v��2��T%)�Tj�N�',T��uO�5JU�J�T	��	���E��MtK�ƒ$�U>�n{�W8@�j���R�Pi��~�4l�79I����b�P������ί_�������]bѷ�鹝��Ȁ�,�%Uژq��8�-���v��$���#V�vo�5P��#T�L1TF�0�\����<)IO�� �T�B�k76!�e��B�%l&�-*���F^�LW��ǈ�T�v�z���g����x��NZ���:=8Wcwv�M�+�$��y]�s>���[�'�4D5���W��'��F��'I1����Yz�R��Ҵ2����{qWb�CȆ)!�Ǧ�)Ɔ�ˁ���Orc�]oν�����:J왲z`�0�ttY���܎����!;�4� Nc��Kb{	BP��	BP�%	By	R�Z���'�Ψ�7�95��71�o�j��(J��)w��}�'#u���Z�9a�%� ��p����kԤ�Uq^M%"��31T�jc)J��6
�v�{D����
aDc��/���xj���$3!�J��2�*ڏ0��g��ߖ��b{Ŀ7�74� �l��t��m�i��$�M,�!�,Y�AmPU�KV܆h� �e�X�b��]~X�|��R�e`Wd୥ej�`
B��j�&�hm�ְ � $#��5|     m�    l                 6�    ��|   $    �                �   �`�                               �     6H�  �  ����[d  �    l             -�   	                  ��     p     p    -�           $ $              ��       ��m���;mʷi�c�$�k�ց   p���dit`    l�����   9:Hm�5P� �ڐ  H -� 9#[v�Z�@ k��l�I�K���ҡ5ʠ�5*�` �HH$�  �p�(n�H���qmpq ��6
Z���m��Qi��H�� 6�Lՙ]� �]�3�,�j��L�K<�u���j�e�f�7gl�yl -����:ؽ.ҭ(<!TTph�j�l�r�2Ψ�-l�ۛIde��M�[���Ҥ���qJm�L��k�� -��H^� Z�"@,�g8m�]�#� ��ZL��[����$[vi�K���ݖ��ЪUUR�K�Um�5ɱu�-� ֶ�]&A�m��u�%�v�l�hH ְ xI��m �ٲ�6٭`�[C�l�z�l��@ 	 �    ���մ�  -� ���� M� 6���l�`H �vl -���-�����p6݁��-��H-[$�}��}h��E$ m�g@ �l  �>ڶ�-�l�A �`�`        >� 8�J �P0 s� )j4<�� ���:*��@R���� )I�� (0 8��5�m� � 
P` 0 8 ��:��DSZ�7l�(�m��Xghm� m 2  �'m�m��   -6 -�-�b2L  �ky�۲ȩ�I�
�[m�iT�U��L N��Im�r@�����s�-�6�+U+̫UU*���=;v�Z��Uj-`� �  �U!s�^�C�٫�wN� -��(�m@$MSK�z��`m*����\mW�i�l��R�egk����H[mF+�į*��&����[Y6���j'H;H,.�l I#%��հ�"۷l-��@m�6��oRFٶ��u� $d�bKkm�J͍�l�R��    l۳m�"MU�m�m�Z[D��p�UUAK*ʻ���*�T vS�vӥf�u�r%�m6�m䜶� �  6�k��lܝm�g kOſ}�A�P�]�6�-��� z���O�ﶩ��<��e�@PՌV�UP��	)��$k���v9qp�������u,$7;%�&���	���>nQT|\��ܪ�uU�v�A[(�56؛`�f���C[��j)K��U4V�*\u����l��c�*�,��t�ZD��J��N9�L��� �����c�:>5�;*�f��*��r��Ig����Vv.mν6���f��n�n�9R��Urdk��uM*�m�UN�)��h
�o=j�V�E=P	�o[��9|�UR���XT�5 T��݀  Il�[zW�x����U�(�ҭA66� ڶ�Jhݬ�{jmaA�׶�j�NQ��
��%[^��t��I��`   5���O��$�n� lrޮ$m�Am��2tݍOT�&�����\p)l��!�f�m�pp��Y1��5 t�㵸���y�T� d6��3v����@�m&&�bN*E6��&��M�7���@)˪Ij���V�eW<�\�%-�V�ݖڍF�D��#.Iv�k٤�95ث$*��[ kX�izX�g�(P�3i^kU���qNҦ�R�WU.��q�et �-���n�@Uیjhx�T�֑I@�����@�kj��}�G,����6����ZuX�n�ݛ;K�O/ca�-@ ��MͲA������;J��PP
nҬq��ڎKi�(��J�M�^��+�@pᮇZ���*�gXqؼj{oL�T��ob:M��L�+qہ�X�5)��/[�]]�5��u<�����'H��,#a�R��4���\�����`7�=l6җ��`,<;\k$J�UUlp�V�b�j٬�2��-����
�UU[R�\ʮ�ٝ�� �Y7M��h � l���8 6ؐ�Ül�`nG�l���m 3J����&m��� %�	�M��v��@  8	 �BF 6ۆ�Mkʵ*�*�W[uǴ�v� �ۭ�m&  -� �mk�[׍�ɶ�k�UmJ�*��UZl &��z�n�ڀ���I�6�m����k  Y���78Y� m�V�oUA�t�UVQ��*�ꭠ m�H��`[B��6�m��%�ҳ�T��o:�v�v4m��\�4Q��m���[z@A��\ ml���_LÒ��,�Zl	��D��j�(7` �)+���f��%c��FtT�k�2�[KU*��u@  z�[$�@[Q�����P �T9���mӀ���)�u� 4Iפ)v�d��oIpm�j�63P  n��z�[\Aj��k�Ӳtf�f��oT��Tjh*E�O�[�);A@�J�@e����We媶���W�U��]�mUJ���RQT��
��[jeブ����u żX�n��� J�un�*�)��҂� ��J�mҭ�	�%ݍ�A �J]��A�vN�E�*�UI�d��������&�r, ��ܑ��m��讠��d�N�V�UQQ�`���vnK$�9�S	/9f�!��v�����:��^j���v��vU���:mӧ\-�ssV���M�5u҈��Gdy����ݟ���v&�e^x�h���m+t����Qn�i�Z�	)]����`�v�W��ؠA���c��[��"�MU �қi��%��Ĳ҇$���H[<;ܐ"l�]��qum�޲t����ü�Z��9�#�rMU9ʛr���QV�ΩD�M�� �[���7)��`��j6�Ku֧c �I@ܔ^BBr�UA�wFoX
RM�
vӅ��l5��@��hຂ��(-Oi㷌M�hvJ�덥Z����j�I@m���T����Ǘq�jxU�#�q��y�ŵ7�8{�Z��Z�j�ۃ��e:\pU�]/(�¨�2���]��P�Pp�h۫d��"v����Ts7UU++Uշ��y�*�U[/k���9G�;����ێHj�)V��Gn���Nk��6���a��[u�6h�� s�$ �8 3��iΆ�#����ӄ�H�e�@�;i2�cm�� �K����I�Kx?��| h���J�RK�$-����3��/�W3m��8�@86���{mŶ�E;mRI]�ܐ�խ��ֹ7Y��Wl9%�U@U[:��fX8I��8�� �5�v�ٺ�ࠢ[��+:	NZ��5ԺM�-�g:��Cp^�nIh'X*�R�ܥ�<;d.��u���7Y`Ueb����-)@ 	j���l��RZ�VV z���ؔ�z�t� 	 lڋ-�@2j�a�Vn���o����O�Wi�l ��N�d��ƭ'L�#8`Hv�H�l�4鍕�z�����UT��e�<��i2o$��a�����`+(�b�� @U%D�购����l������*�NU��_!Ĵr���Uݝv�ދUh� ��'�v�]�]R��=R�q�1��g9�K��`��[nl�LI�.JsZ� j�.整6�i��0 1��8` M4�]t�$lm� 6���KWz݄���  6Y*�-��kl��������VSBѭ�atuUJ�	'n -�mp5��'m��L�֍�I��9m���m�-��e:�$ �vj�����4��k)Ki%����)��AT[5P��t���<���:��YF:��8��D�2lm�Ӿ��d��6�s��:*���8����7UR�6�$s����rI:R�@i-ķ�@H�iҝ:n$�m�-�n��`h���ω  8    �| 6� [v�-���P��w������@G�����@8�'����xbO��(/`)���Bz� �j
`�z�N��%T�G��;P^ �t"p�(�Q��<]�.�Dؚ�f
� ;���+���*x�B z:N 2�v�B�Oi$��@E�
�#Q$B]��D�Q4
� b� ��(�( B&��e�A<DN�ӴJ����U|GH����DO@_ C�Cbb�B����.�W}��`Sl51������ęb�I��Јv���Ҝx >�/ّ���a��""�`����`�UH ��N�v*�J����`JF��!�&X��E�@�S��#�(/���
a�j��RP��] �j/H��HT{ABҁ�#�ࠝ�¤ �������	��P����@FA1D_E���"�������o��������'� �ie ��P�iX�a*��"I �A�� �!(ZT�d&��(J��(J��J��(J����Z��� ��(�	 !@���(*I(��(*E��(��&Jh("(�"e!(J�����*@��@���Z��(H��(J��	��(���Xb��T

@��g����a6��i�̅�hډ��ݪĹ�����    ��m�  h��@   �%�s�m�_M��x  ��`  �    6��   ��Y��"].m��tj�Vp�bd�I琥j�AM4�܎1�f��F�6��;�tD��5�ɜ�0��'���H�悸W0���B轆z��ֻuJ�&�)�<�
Z�T��;�LL�����%u�R���) ʵUgz�I�@��^�5����b�崒N����Xt�֒ �d�m{jUzqҀ�F�0t�OU��[/gЕ�\uz�Rr��ѻQ��u��h�/$�6�7[��D���mʵW`����@T�s�Vd�U۱GV;n5F��=	c��vGj n%�<.�=��m�<�e]<�y�M�6v8��^��\�K0��2�wS�k���:mu;U���bci��eAܗ���<B��=�؎�fU^y���m�-J�n��n����{x�ț�B3KGXZ�n���9�mՓv�d�SRј�Zv�kv��˸Q�èn���USֲ���ѻ[�Ĥ�vU�cgZWO3��3�\l����)l�[�@�f��X]��i�UW+�;\F�,���[s����eلj;���ቛ T�J�=�J��N���BZ1�Ӈ�B��n�[��l^h*��f .-Aq�պ,�3ӎ�ϰ;v���森���h,ciKݺ܃X�b�x��s���C�6��T��ػ9���N�6l֓�]q\x{S���yM���xx�\sb�s�9v��𫳚�T=�XŞb���LޭNlH�=�V����t��n^&ݷ`���UaY���rC',�H�$�	�BV�J��6�����м�Ĩc��]��f9l�K<�E����jA�b�Y�l���kp<��������\9Z�	��d{skUmt�`6��ι��\�T��%�����������P^�C�*��t,"��'��SJ;7�"2ݭg���[��a��yrcq�UT��n�m�[bT�]-���vaWM��^JW���u�z�&{� ����,���[��yV��ۅ�Jv���ۊչ�!q�óu�,��gm�,�Gjѹ����c��ppppo"^u�RM�䞍�jhy�l]�0<�Ԥgs$��M������<&����r��q�Eq��XӺ�ww��B���P�` -�d�$��,����>A�{e9p�{sǗ���ȖԐ)�MU
���zՁ�zP9�v{����+�N����5H�t���O��������oZ�9s4ꢪI��)�9n�'����mq`g��X�,��o�:�t4�5N��mq`g��X�,�o; ����R�6�i��]{zՁ�������3�\X�J�NC�Jm��.����s	ɝ^ۢ�r������A�3�t�X�J���a�(W|�~���2}����{zՁ����eI/fo4e��ַr���=�17Ҏ�S�\��q`{w�X�,�'5(��<�N�N];=�Ł�޵g�B���|X���}4D�*f��N��3�֬��O���������ʮ�MSNe��N���������3�\X��VO���rP�t��U2���v4mX�N�a獼ۍ�[=3�#vz��.�<]nmf�ݖ���+I�/���3�zp���=�Ł��9|�RsM�T�d�;=�Ł�޵`g���2}��7��)h(��m:�E��޵`g����P��	JJ2gz݁����=�����]:��VD%>޿�ӽ�3�\X��V��s��$�SRԕI�E����`g���3�֬�������ۥ0v<�:�m�щ���m��7V/�b�Nf�U��Q����"���{%��Sn�������oZ�3�\X>�vO���(���E:���oZ�3�\X>�v{k���*�5M9���U:V{k�'��ϒQ
g���`{{�V.f�TUI5R�1�-�`d�y��,������	(Oz��'��UI�7HUI����,���7k�'����.�<YHrܸ�t�\�u4�4�v���e��q���J8��X��M��m�uj���*J������n�O�����ŀ{˧�*)�Ժt73T�ݮ,�o;7k�7zՁ����eI5DԵ%R��2wy��\X�֬ݮ,k��2�15R�t�ݮ,��Vn�N�;���h��T�H"�Q`f�Z�5$�}�ZX>f�~��@��8����@��K�T�8�K� ��m�6�;mei.[Ԍ�[i��e����WV���54u܄���?9��\��nzv7Maj-��n�.v9��^�Z`�s�'�HbI�]����[�m�]���9؜���C�.^Ś�U�p�яW]n%����]N��>wX���Nr��9$��:i:!�0uэ�r���i���8�u���6�����׽��t7�|+��؆���ι�<JM�IzV��8㶚�~7>���8{6�y��GV�z]��]������2wy��\X�֬\�:���j�JcM�E������)����`{��Vn�Oh7Ҫ��n���S�3v��3w�X�\X;��=�攴UU6�K���޵`f�q`d��3v��yt�E1UK���j����Ł���������޵�m�?{~~!�kۊ<��r�I�V�����k�
�<J������l!�غ��S�RԕJ[�����`f�q`f�Z�%��p��E	R��H�N�$� �<߷����	���D��ANXLU��Hd���0�ch@Sb��B�*�-X�,��vO���(��rH"�Q`f�Z�3v��2wy��\X^�]bt�6)i�N����Ł���������޵`r�i�ET�U*X�m�,��vn�n��7k�}�2��M)��`�tU�zKV�/J���ۮ��9�=�ln�֛κ:6We�UI�7HUI����\X�֬ݮ,��v��sJZ
*�&�N��`f�Z�3v��2wy��\X��z������P�5J��������e��2IBd�(�2t�=����dK�rj�r�*��E����������޵`f�q`{_m9�ɉ��ۧ`f�q`f�Z�3v��2wy��&9��Y�$��K��=D�>�&�%�gW������쏮WK�mbLm�k|�~��ε`f�q`d���!$�C���`jޕ���T؛T�X�\X;��ݮ,��V.f�TUI5S#��m�`d��3v��3w�X�\X=��J�Ni�B�LuN�脢���,w}j����ÔBQ1�<���{�9�-55I�iԺ,���7k�'���������2s�N��SE
G7]���+���#��N[R㖎۴K����cV��I����n�nһn�{�N��j��\X��V��s��$��U)n�'��������oZ�3v��7_m9�ɉ��ۧ`f�q`g��X�\X>�vO����Q4�D��A���?�͵@}�:P�{"�Y�O����ս+����6:ӥ`f�q`d�y��\X��V���k����R��PU�/n��$$�l�t��e_M�ݶ�3y&�ه\����n]�bp��jܣy�Aح���̰V���h뇢.����Z8�ь�99�œ�%����'�K�M�S�9�u�.'+��-�u�����7��'YG�@ع�ѱ�[&�אgu���M%瀬w@>r�f3����b���<�+���7�$M;�9�6��"�/B�
*�lm!���n`nv��"y���d�5��D;���؎.+�]�:�C�:�F(2s�n����3v��3�\X�\X=��J�Ni�B�LuN�����
"��k� �� ��p;�J�Z�۷I�iԺ,��n�O�����ŀ{w��J�J��tSn]D%����`zw�vn�{k��˹�ʒj�r�*��E����`f�q`g���3v��͞d�cj���TL�Jf�K�f�DbŹ#��q�YT��]��H�>^mY-�r+�!��)15R�t�7w�g����ko8�{�M*UNIS����ŭI,P�CM������w�y{eu	�T؛ ꨋ�޵���^�����#�rӝRMT��4�uko8���Y�|E��Zø%𪓚n���S��޵���^���=�����p��aL��)�"�ڞ��s�NZ��v1�/���䬻I�:��4ܗKEMMRr4�j�g����ko8���n�t�P�TU:n]{�ְ���޵�����H[�}�Ң��ʥ-�/�͆�{�X��I�/����E2fօ(ѐ{$Б����Ht[��t��#@�:ٸ�Df��������&I���Dw�m���2J��4r�x��#��h� �S��h3IGJӸ"(�َL�&6R�f�xo3;�%�����1���ѭLLƝ�h��FPƣ
���%�A�oQj�љ��L���CA�3ZZK6�-奈2\2�k30ц�Y0\�h�v��}1�Ptkp���1ě4u΅sxd뮉�3�4OQ���c8&��I`�#AdD�l��m��pX(�h�C�G1 ��)�I,^���m��n�t�B�'Op浮q  ���3��t g{w�"9ӭF�0ְ���n�!0����Jfa��b�s�>p;v;Q�C�UN�j����G�O�@� *����mE�M��ǲ�u����)I��}���g���6�'ɉ��ۧq"2�36SX́�}�:S2d�3v�X�)�{��┥�~}����F���.s|�ǩJS�}���):�߾��)Jw�����)I�����R���>�Sn.�������X���^�nN|���z�*��I�[����;rۙ��mo{��)JN���=JR����)JRw{�m?�T�JSϾ��R�˰�D�.LH�:�4��d���ߵ�)JN�}��R��~���)J���n�k�3/�p4S0<�Jʋ[޸�)I�����R���w��)JN���=JR����)JRuߟ|jiKEMMRr4���(�!B�u|\B):�߾��)Jw�����	!� ��ĔS	TN ��NrM>��J0�A�����C%QT�m��ԥ):�߾��)@HO~���{��ߩ(���Q��D�ck��J��Ht��z*ڥ)Gqn���Nk;�[�v��˭N��)�̊iU6�eR�Uj>"D/Ow��)I�����R���~��K���n�Rk�3,������P��DLqJR���}�cԥ)߾��)JR_�v�X́�|��́�-_{t�����e�\�9͏R��~��8�)Iמ���JS��ߵ�)JN�}��S"����MSLm��\B���߾��)Jw�����)I�����T��ͪf@́��Նđ.�9�kZ��=JR����)JQ��/���ǹJSϾ��)JRu�}��R�����w�￟��4�$�Θz��-� HN�k��'��+���nu����>;2���L���;��,��:��uhF�ێ�ָ`�i�w
��d�ŷ�u�ƞ@���"r/G�0�ƽ�kd۳��ɇ���!u�Z+n�t\��Gh�E��	�Q��c�\\��Vp�9c���y`��v��gkuZinƠ:����+Yȥd��`V�"b"#
���ST�	L�������\�gn{l����un�t�r6��J��S&��Rc�}�!,;����R���~��)JN���=JR�Ow��D ��߾NiKEMMRr4�o���)Jw�p���'~����JS����┥'w���ǩJR����T�d�*�9l��q"B�ﾵJR����)JRw�y���)N�ͥL��2�n�K���L�(h�Q4��JS��ߵ�)JN��=�Cԥ)߾�ÊR��w��pz��<�~�kF��f�7a����)JN��=�Cԥ�gϾ���)JN����R��y�;�A�F��� |ܒ��S@MT�G�%=r.�s��<�T���ű��u=v皃�-�V4�nI;������Z����w��pz��;�}�\R����ߴ��V��VӚ)�6�
n�� ���>���~G���hnS��ߵ�)JO;�~���R���~��?(�wf@˸էD�.�9�DD�&���<Ͼ��)JRw�y���)N���R���>��ԥ)�}홯�z�f�l��խ�\R��I��ߴ=JR�}��R���>��ԥ)�{����{~�9�-55I��v�ڌ")߾�ÊR�����pz��;�}�\R�����~��)Jy�^�s2�f[��:n���s	��ۡ�q��z8��]ӛm�t�Ҹ�6s�K�f�Jw��I�t�<��~��)Jw�����)I������Y2�3iS2d�sv%���b4N�k{��)Jw�����I�JN�}�cԥ)��~��)JO;�߸=JB�率�|9b�%9t�!B]^}���)N���R�"��=���B��=�� � �T���k�3,}݊f@́�/��TB�#�8ࢦ��5��92d&^��T�R�������)N��~��?��goJk�3,Y�	臒aA�[8�)I�~���JS��ߵ�)JN�>��R��~��)JRw��}�ד[m�Ob�g���:�^K�S�y�	�e�R+��n��{p�u�u��ay]o�ԥ)�{��┥'w���ǩJS�}���)=�߾��)Jw�{fk�S�4�T��� �A���R�")��ÊR�����pz��;�>�\U̓$�ِ2��yC�xD��ʇ!=TUlz��=���8�)I�~���JS���S2d�73e5����͈�*mXn��������)JO{��=JR��}�)JRw}�lz���K���q"B߷�LȦ��h�T���aR��}�)JRw}�lz��<�߸qJR�����R��x}{���fg �	y�]�:���tB����2Z���n�ض.�����'8����{��Rw}�lz��<�߸qJR�����R���k߳�R���}����F���5�s���)J}�p┥'�����)O�׿g�);��߶=JS�|���i��	�t�!B]���R���k߳�S���<�}�퍌��f�*f@́��j�bH�y�3ֵ�R���k߳�R���{���)O���R���'�}���@f^}��8S<�(S*e�^��3 e������R�>�߸qJR�����R���k߳�R��P��>�5�?��[�Ͷ-;I�[A��;�pj권�HVډ9{gb�sv��WL� �6���%�HduwK$�;:m£e��e���57��Rks���)���s��!r8�tq�,�p\��n�nv��9`��:�Z��9�j3R�B +sD���a��מ7I�t���g�d����;g�'S��n��������6ݗixC��a�F6F�[u�do6��.h���feǶгmsM����a�)��e����:���iUUN�I��NiKEMMRr57n�t�)��߸qJR�����R���k߳��JRw}�lz��/���kf�ڰݽ�-�37��R�����pz����{�qJR���=�cԥ)���È�pI�d�����yQ/�L�4��)O3�ߵ�)JN���R�D2S�~�ÊR��y����)O�߳D�|9L���w�$�}��(����~��)JO{��=JR��y���D ��~��*ƚ�m� ��]�z��<�߸qJR�{��=JR��}�)JRw}�lz��>����ӚX�[��Ms״-κ��&�㳰��C�M˺�����ٶ3�g�{�|�<|�i�+lR����>��ԥ)�y��┥'w�{��:��<���qJR�ϯ�o�C��j��M6�Z�"D/N�󴗡/�� 	���Rj���lz���f�́�,�۴�ę2��G��T�4M!U&:�q"B���ԣ�Jy��┣I�~}��JS����D ��o|�ԍMMS���ݻ�Q�A@>y����)I�~���JS����(F���}�cԥ){��kf�ڰݽ���Y���)JO{��=JR/y��k�R���{���)O<�\R������~}CL͎�=��Rf�:=s��
/R���W�i�s�\��Ob��;��x�j�oz���z��;�>�\R�����~��)Jy���)I�~���JS�率�|9L���w�!/w}��?�������\R���Ͽ~��)Jw�}��R���}����F���5�s���)Jy��┥'�����0�QتD7)�{�Z⠈A���D �Z����tSLo[���w�F�����R��y��k�R���{���(?��}���3 f@��rӢH�y�^P�"&�X�R��}�)JQ�(, ���������́�n��)�2Y�n�k����>�ɟ��\�#R^d���e�W����*䳗c]���6X7f4to��{���w�{��BQwD�ɊM�M!U&:�q"2�۽)�f@̽�)�2Y�n�k"D/N��!{��'5#SST�7h�s\�ǩJS�=���## d�'�}���JS����qJR���}�c�*?�%rS�u���m޳�x����n┥'�}���JS����) ?#(�_���ǩJS�~�늂!-���ԓLSRC�cuj0�A ?���^���)JRy~����)O<�\R���(H	�\�h1Lqc�0YA0�ZR$P��~Iw'����R�̹�����%�&)�2_����d	&nHf��♐3 e����)N�Ͼ��)>��r��Z��5��lm&��]\��k��y��ֵ�ۇ��oe�ٗ���#�B�ea�*ƚ�m� ���6=�R����\R����~��ԥ)�y����C%)<�}��R�������%� �3%3 f@�>��M` R��}�)JRw}�lz��;���p�H"B��ˏ��i�9i�޷��R��=��qJR���}�cԥ)��o�R�����pz��/|�־�* ��
eA1L�$܄���v�Jz��?{��)JR{߿}��R�NC&���d�{ټ���rI��A��͏R���{�)JQ�(���I��3.|ފf@́���l������th��I(!��"@����s�!�L�f����:�XY�]�35�f��4����!�%�,2((��
"�#ӆ�X�8a�i�nY�Ξ�]o��¬r���,=�#��0����y��:��CH���I:�1�6:+;-ka�,4l���N%��.��.RKSt�	K BBD���NU����VɆfI�Ri�ab
����[9�x�m'�'��$�H���xt�#�'i	��8R��mNL��a��#��7]�}$t!�3[��mb8�A�}�@�|Ԟ��Eͤ�KpL����@XK��C!)@ݚ*�W�5֍�.18�h0`"F$���0���aR	
IHd�H����V�0w2�)��P�0HKDMl2�ZB�c�h@j0�!)q��AK��`��h
F �(a���"ԗY���	hJZ�dHJ5Ѽ,ĳ���Ѥ��`!��Ѱ�l��Ͱ ��3���^y��&.���݄Gĵov�[��:3F�٭��x	��Ri�Dj�V �n�9&)���9V�*k-n)�+mc)C���ڻF�dH��h  ���m�   �a�a�   Kh�m��l����  @m�    p�p  �[p  �*���
-��.ˤ�̀Zqi�n��ێ-�mڷE�L������d�=�ۜ �5��o�m���y*�s�I�����P]y�%̘�m��f���[10��1Tу�u�@uUU�t&�6^�P�&*ls��h�s[mT� �\[A'	0�ȸ`8
u-�9mr�j�)z��	�Է7P��׬bA����gv�;=9��)f�\��ͻOO�sF��b�|.w��-=��h=a�k��j�ɇP^�=+[��yZ�mGr�DoS#�wh��c�x-�ݰ���p���u��e��5��'�Ɖ�vrJQv�MrJʗ���K���jk�ɹ��v��7Z����U�-����OI����/FltA�]�<��%�"�kd�س)��X����b6�-�0!�����-�h�V؜v��ܶ]�hb��|fް�^u��7��޵mwtܼ���K��ѻ���e�9��r�cY�Ji@����<q��p���e�;g!���Z�0컰:	N	v�awj�n�V8V������];��u��9J�;sg=�N��N�ֲ���%e{��N"�7�13�kBI/�1�a,ݼ.���mn�=Al޻�e{*��ɗ���q����WU�{<�m����m�G�n���N���^�ݘn�[F7���
��|>V8�3��ذ9�c�����Mp�M�NWts��c������Rmk��Wf��$����gs�ՠ��s�s��WE���H���[gFM����8���%9m����4�j�V�O6+�M���rp\貲����ʜ�wW7n&ɸ�vG�7E6�Vɝ2cn�YP^�Wiٜ�S���$mb�m�2���Ŷ�\��7:p�Źn5.��G&NF8=]Q4���
��Y
�~���ܤ
�� #"'j"P�@�tt��mU@D��=��VU|EP^g~g��4oy�T�[�m��n��np�յ@]�-(J�����j�̶˳m?ߔF�� ��u*�x9�����N�Mʓ��-�"M�H�u��gl'<��b%�6jcmϗ5��R N��VB�cZr\8����*�և	�מjN|N��#�V�'m��f�6���m��3n��$�v�&Ѣ]�֜�ctn�/�`g7�ۦT����T��I\(�`�̖�Ӣ`G�u�jh��xn�y3��w�q�@��ɶ{\1oq��J+ֹ�[ѷ7���޷���)JR}���R����k�R���{��T�
)ܥ)�߿p�́�v�D���yq�f���3 f_g����XP�JN��}�cԥ)�߿p┥'�����)O3�s@�ؾs)���.�� �A���BR�y��8� ?��RDrO��Ԛ�d˟7���3 e��0��hݮk,�\�9͏R��	V� !S��~�┥'�}��R����k�P��%	�a�����~��)Jz{������{і�odY��R����}��ԥ
� !B������)I���lz��>�߸qJSow���~g���v70]"Wnby�Z�S��g�@�b��G�pݵq��S�w�����{�����-Y��S4��-4۪�"3.|ފf@́�����Đo�iP�٘�D���C-�M�k�e�پ���B!f�1'Jd8�E��!��ֶ�Z6�2E`���淼����A����4[�Xk�&�30L��4���\ڼ�	�`oh�	�0�8ؙ�/37&0!����@gv���͊�!�%��J3{�!�&bTA	l�ߩP�n݉�s������zl�n�)g�`���L��f���͊��͛2d�ٴ�M�;/�t�v|�Bo0	~ظ\ݏ ����ݓ0	r˭BU,i7��n�\k5��%��GY�,"�j9�fK��̒�֥�J~!	Buv��9��T˗N����M��ͥ@gٛ�HfL��&a�%�?>��=��~�VB!I8(����7ٴ�&d��22N�޻�7��˛���H��v��
��[u�=��~몾�=�\�>A1�8
@G�
w*��(�J�@A#,		
��( C
 4�0���y�����+�v����
��I$�`>��I�2o��fK��~��������T�ɗ$�f���Ӣ:`���
eA1@�d�	36}�@gٝv��b���Բ�E��>�2�t������J�\����L{^5�q���5��Mq�䌚���	�jl}�4}�۰5��ɒ.nǀo��S�ݟ42���� ��˱�2f�o��6�͚I$�����U�>M�7��l\.nǇ�$�voM���{"��u�]��b��a�3�#���;7���ٻv,ɛ&JRImf�P��مd"�Pよ��� �f�ə�;$�{{��?^�ˀw�lX��b�������j�u���h%�n�v��ŭb��/F�r���MHQI%n��ګV&�E����f/� �ؾ�� '�>�miv%MۥI$� �틕�U�)�`���=ݓ0�����"Q|Э���	��;�6, �����f/� �}����m:HUfs�X��Q=#��ɘ�ظ}U��)�`�#T��g���i7�=ݓ0��ꗻ �ذzG�7��}U���V�I�I�k u��o� 9!:(ʵ�z��O;n�Gg�!�!faQ챣T���P�n�muu#h������XhI.\�8E)U��74z2vn�,����vc{�u�k֌�|���Y4��s��^5��ՎGl��Qw�c��m�_<+�9s՝�����^Z:���r!!�6�a���+������I�l[t�V��X���m��:2�m�]+vn����nKVw6�pk��z]�.��Vwb[A\�d�� ���}��Oˀw�lX=#�}�}@{�&`wڕ%�,�!ݫMp�76,L�2�fI�=��@g���|�\��65X*>;
K�� vl|�����+(��$��������\��?���whMP�MЮ�|�?)$��B9�}����=���W^k�~�U����)L�2d!$0�?�zhq�N�"eĩ�t�$�`~ظyM� ;6>����%��i�c��7hT�Vؖ4�[[%��!���-������c#mv��������R�!��h� -��\Y6+e�)�Bmp��?, �������(��U �%BN��=�����ԭجciҤ�3���͏�&Z�%�I�L����`k��P��ؿ�U?�U�	T�����m���Q��w���7;��1��~L��fM�&��f�����������*�&`���1��ލ͋ �sf�&K�ə	0�����v ���<��I������sb�I3s0�$���3��x߶.��w�V]]�n���n�#�U�.�3s��#s8�\F�ls�h�jU��S㰰���q`f��=ݓ0�l\�����ذW�W˻Bj�br�w���f������ٙ�����:~Xٱ��kH���*n�*I'�?�b��ѹ�d��+I�:L�ۛ4}6f/l�_��j���H����2d��ދ �oM�v�f���e+v+�ut�s�Xٱ������9�m�b���i9v�/v���	��n��������=iNVޝ]�/Z4p��;�w{�����9#ZI=ݓ0�l\�Sb�͏�l�q��yP�h��"n���lW2I	�~�3c�~� ���h}���$�vI7��h�����~w�RI��1@f������wd�ov.�ڛ�
��������K�������ou�����_�$��)L�=�8�)C$�6Xĭ-`m<U���ZϿ��������К�X��]����f�� ��lx�#��r��n�e:;s]0����p N��MϢ��]�Н��i�6M*Ē_�		'�,1��n�)55�����͛ �wf���3!&d���9�Ύv�Q0�P�T3��͛��&N���=��`y�6+�@?��%KY{�߿�Y���蘔�!�U6�����7n���lP�M� �)���>h�]�o�U��ɓ	!&&|��]����@|��ٰ3.I0����-��z{y�Gq<�v��6��`�e��M� �)/�{�}���ށ�d:�XL��2ā1IB	�wߟDkY��޳Vŧi0������xp!:	zY M�y�#Vgh5 J鱺�\�A�v�;u�=C�=؀GCs���5)����0�m���|s�u4*ϡ�7b�'0;v2a�ywT)_�4|�ŉ1l����[�`��·[�k�:��2�[׭�#�/7mϤ7
���f�4�^���zwk:7q=�n[�<��7	c��ܱcH����izͷb����s�������շ�؞ѧ�ɺ�U��n!n�n��-��ߝ��$("R��%�TS��l	{?�R_ �wf`�e����1d"Ը<������3Ѻ��33!3&��d��������nl��fI~I	&Pj�ߡ�����C�2�y�zs��`�e��M� �)/�vZD�ۑI*DL݀��s2IgN��>v����z̙��_�L2M�߮��~_��:MU�)�J۾����%�wvf�_ �x�����郵�i�]U>�&b�c�W��Ż��ְsh�n+UN$��%Uy��H�:t�6���}j�����3 �[/�e�lx�M�R�JS��C̽�6���	���cp��������k�h��Fe�.`!��9�ҏ�/`v�~Aa.��|��;zl�n�2d��&Bfp�[ߓ���+j��hM����|/�c���$��r;���n����:4qD)&�"^��%�3!�'���܎�=�f݇�I$�:w���j��!�����MUUM���נ���a�l��W�o�?_ ����	��������h-��^з�]f��h'��tWV��o�z��8P�#�d���whMP�M��x�Oـz-��2�6?��� �)/�v�D�݉1��$���l�}U��_�ǀo���=�٘߬�.��5V�n���[�sf��F�������-_3$�L'L�AkZl��15�l���4�eU��� :���L �	&��L��|N���|��F�66���q�w� $#q����� �Gt(�e�A&&��uM)�5t�Fx�`���ѽ��^w�/U*�;�4�K�	J:#�$ (����J � ��&�.�������/0����j�;�HfZ1�5��d5���h\љ�63�h&+x�ff�TF���8KL�C�#f���h��ON���Q�ڏh�#Ђx���|��@�A6"�"��'�3$�}~����/�f�yrbħS�����fL�>��=���=���̗����|��7#�aK9)J�Bb�n���3 �[/�e�lxnl\���ߟP�3c�qG���Yi�qcq�l��W�^L�+ϴ�Z��l�F���6�"�5���[���+j��hM�MS���M� �����+d�/̐ɒ����v �â�����w�2�6<�l���m���zI&�Bd��嫷�,�D�0.�f��to=�n����z ߻��V�󛙖:hr:�u6
"$�L����r7��=��V�*��@���4	���� �$sM�+.b2P2$b��(��a$�~��l�/��F袓Q3vz3^�f�36v�W�{�~���f��+����.��j��6�v��v���巑��3"��1��|����C3%5/Q
Hx�O L���z ����;���&`��wղ��ۅ2�2�����צM̘L�p�wu�T�| �ݜ�7�F��c�t�/@gۻvz3^�&���9���`{򟯀OVȝݖ�[T|�Bo0�f� nfmXlf�3s�'�wu�~$.�G�E_͵`�� Mݜ�;�������5��ʱ�dX8�P$B����}}�ٳYh��ff��u��v����[���  ����Ԍ4�Lm7��Yqr��rY1Xv�aj�����3��LC=v�=Ony����<۳H�-�Q6���V��]�!r�-L+��_�=��3�lI�i�^� �i:zW��Miq�H��q]hnwо���l`��E�୸MuwIi���x�k)�u�:�1�([	�uh8��h'�6��s��)�"��n�g���,���X����X͸T�+�"�vG�/�{��v��p�M����S ��&j�@�������݁����I������1gt=;�0�r&P����bL�!��9��� v��Xlf�$܆L��v��H�q&1Ҥ�y�M���	���b�|vI��\�����M3�U��3&d�n�U���7�ݻ=����l�n�v�7E7Y���0�p�R�337{���76x��ͫ��ڇFlv�(����Mq\V�]�*r<�8V:M
�D�ɹeʫɆ�w4�}~�۰3�:P�f��d���‛S����Jڣ��y�o�×J�] HL��$�D0�
v*hQ��Ͻ��uWd�@gۛv.d$�86`��]��3PnoU����G��'~�o]�����Ź�B&UL˺�����3/ɥ�M��� ~�����J���eX/��wi�T����8�l��_U|�d�sk� ���>ܝ(�>������nc����I<�1��'n:�E���.�wl�n.�\h��A]F�\-�s�����\8�9�vk�>�����3 %K�S��]:]�� zn�`���7�L�7��ʪ��e+v+���Dʲ�j��'J>�۱�$��&��k� �����X�!�Cm���'d��o�ÀK����p������+j��hM��� U}ݏ ��;$�nYu�J���_Jݧ	q��բ����c���;���<�<]��Y(�M��*i}6Յ�p	{�ٮvI�_`�p�[65����Al���� ��;$�}�_36o�swCӻļ�2�x���wu��(|�ٰ>ܝ({p�rG�O$�DD��s3'Lۛ\P��~�Uw����q8)��
o�$�ה�v7ut�n�i�^�ɰ92^�(�w]���Ҁ�c�}�v,v�9�q��a�{%j��/3��r�ϴku7���q&�ӯ_
u���f��·?�� �[/�N�3 �k�>�	{��R5O�S�0hi���L�7�r��fl���z��fN�{�]�yP��6��`~�p	{��_ ��f Ct��E��v�Ɲp>��{��_ ��f����2�lkCuƂ����q��e�ꯧd��7�r��ݏ ������JbtZLv�I� m���v�p�V�rڹ��=�v��z!�f5(
�s[a�a��HKjܣy��lV����+s#V�tu0W�`S&w@C�Ng�7g;m`�4\	�36W��O���1t�箘}��3�4�H�8��-l��;�u�� ׂ����ҥ�;kz�W��7���˞PV�L�ۧ�Ň�a��{6*��1�btv��$L�Y8���u6#6�^��ۋ��!1�+ѓ�X���Pv�Y�y��DL�"%����`g�iP���̗���΍�=�w8�y��A*)$�`�9\^�ǀz-��'d��d������A$���ԢeDDʠ9�O� �[/�N�3 �I���V�V�y�*Q2�ަ��L̹3!gN����=�J��fL��7w��ݎ�,�0)%��&^�߷v�fI~fL�������I���e�	�"U.�n�4n��r�[��S�v�8�\Z]N�{n,�̼�؝���[i��n��&Л�}'+�}�����>׿g P���,W{���8�B��e�ܘ�@k�f��%BYXN��=t,Y/�M�3 �I��[65����@�]���T���z~�۳�fI�C&LߒI2��e��~�@~~��6�3W����Л�w�'d��vI�����`33%ə��vw���a���դ�:T�o0�9\^�ǀn���'d��zR���ha�؆�
�8�,i�u�m�ьkn�mt�EnW��[d˶է�{��C3J�� �^^D�Q2��$�9�w���[/�N�3 �;^���؇t���<�><ul�W��;$��8p	{�"��X�)�CM� �����������%$ ����E���XB���5H��`@'b�ͮg�u�x�?_ �Vȝݖ�MV�y�wc� ����ղ��0M�����ۺi��K���
��j�|vI�v8p�e�
iYut_�2���tbd{j�YnF�;[.�&}�F������s��畷����wW��ǀ{V���L�>͝)�.C�>���[�N��bn�w�'d��wc� ������zff�38{��)$x�$LD�����K���j���0���	%�a��)�"Jɓ!�7�(����l�����wn��a!�a2H0�*J���S�����W^�k7���(�SoSS`{#u��3�$�!/�����������6��6���r!"R��	���+���m����q��݁9�G�(�i6��c����I;��L�;휮/wc�;����D��Bh
y�"f���J���N���`{#y�	�&`����l���v:��sf��њ��7����`{7�P�v<t�n��Uӻ��|��;���,��J�325�3f�ՙ����/0��2�LK���݁��f�oZ�9�w����{�r��w�� �j�$1)
"�@�D���a�bPAvX��I6��`b.Z5�K��4Σ,��
ң��Ai��lVM���6;�V`� �
�+À�]�E4���4�A�4&�pМӱ��l�1d���Q\��&�nַ-�-�  [@   ��   ml    8���$�t��   H�     �  -�� � .��m��[��gI���m�Ž��m���j�n[�F���D�v�M;t����^���5灻F�Jt���Y�n�P��k՜d�3\	�(�l#kNlEn���K0.��0����&�!���*�Q�T��+]u�L����"�`���焎)KF흁�u�loT�k�-�Ÿ+�m�h�Ce�es�!t��X�dW��6�>����OOg��/O
��Bü���N�MȢm�݌m��\�5��� 6�imּ�k��ӣ�����M�ݶ�9h�U��"7=�zs�U
��v:x��ϒFH�	W8x���n1n������7k�v��9���V����V2uӭ��Zt��+qۜr���q<�;X3U�f��y��57kJ���W\�]J�U��f^f9�ۋv�h��{���t�ծ��v��}���)�^]�e��]xa�}�\Z�9ޚ��m�v�%�������sیg�UV0d.ݖ������S��7�u�Z�8wkٷP݀��bC�p ��,�"�i*v�՘0U�rǬfR�P7r�����}�\�{sݤ3ŷm�T���[�;�:�>�5ًaܘ�4�2�v�C��s��.�3]u�8^��� �s���x�nKV){Ɛ��`��x��Q6�B��g,#�2oWS�6�]ZCx�V�����#�y꜌�����ӹ�Z^�B�0\�Zk!Ʈ�$��=�gwjJ4$�u�-�s�޻!�5vGgN����v��S�t�&O;J�!Ű��\���С��bq�|X��N^�������d�
���D��'oB��۶��B���-�!mrgN�9�qK�7:��p���6�-s��ݗ�؎(����c��1�ٳ��hrʍԽ�w{�U@�|@;@�W��P6���z�/h���zn�N��ulS����dqm��Bt:In�R��{f��ۘ�c�.l�B�/9.W7S�w5*Y3��/c�t����tX�If�ŷe�D>�j�㮋gmyz]K�y�:.��a�����ok��݈�[k6��wmws%�y�k�û=9Wx�x��	���L����P��%j��(S�-c���糳�sP��Yen�c���j��qke�4����H�
�����LRܻ�z���u��<�b�u˝��gNu����*6���L��I�.�M�wg+�K����\9U��N�3 ��t�5E��i7\^�ǀw���'wv���J���!�_�@{���K��*t7O/�� ���;$������v<�-�S��WLv�����f%�(���~����Ԩ|�ٰ>�N���D��hVm�7�}���%��x}�vI���i�E�<��7lk��#%�s�h��c��墠z㉸	�<s�<�jL�3�t:�o"v�yp��`~�'�w���'d��w�9\+fǔ�*��jUL�����7��.dȄD��`�\��p�DLi�� ĦG 	%q���f���$+J���x���{:����ﮨ���+�K���	[�_.�;j�ڶ�.b^�߷v��v�n�wzl��z��Ie2�-&0�i7��NW �����%�	�&`�l-�;M Jy�1*���͛.Y���{��������Eb�:.쿝&�4U�r��R&�q�	�m�^q���8wQŹ�q���x�-�J������=�K��L�=�r��!ßwzl�7��%H�Ԓ���1@oۻw�$��f�R�9�w�����P�����mXU���`�r��}���0����P�|A�$�D�bc��JM�ưL �@�eM	9#>��ɾL��K������v���"���e��bU�ɓ'���:;���n��	~F��=���ܨP��(��]��ǀv䋀OI3 �[/�Kݑ�o���w~~}��G±�o�g�^�/ɺR]|�����Nl�sk����c�dzA&H�C�92��e��������z_3v[�I|���3ܴ].)�&bIS3v��|^� �R_ ��f��](G����ĺ���	S��e������lI|zI���|;^�W�]�S�eM�UM����Os���vdf�����W��� �cT��ϕ��I;��L�7V���v<�I|��ww���o��4����Q엵�T�Rb8Żs�.'&_��]l��q�������/G�ճ����Л������/vG�v)/�OI3 !!t	T�U�ݻ��|�ٱ��3$9���;;��|͊6lx�R�t�*����ۛ ��f o�>/vG�OlW˻M�+�d�	���L�$��;�� �ޚ��Xnl\vV���Lat�o0}��Ų,�6.��3 _}�U[F(�c�F�p�;������v���Rp!�w�V�v���u�w� Hp�vE�ZQ��+��y�7i���R�A"怴�.�Ǜjmqwcld�r��fm4�Ҭ�;6�T�������C�ʝ;�1I��..;v���X��i6y�������:�����#��ү9��A�<�`�.�@�Ļ���w�'��vݸw&�Kv҇7m�I�8y�]�l<��-L�s��,c�[�b�2ő�=��"�P?
��DBS0Pϻ������3��r�Y�����"A�-��<u�����j�k��Չ�+t� ui��o ��'�v���7�&>�!|��4����\�G�&TM��X>��$��3;���w���c3b��%Ҧ6|���U�mp�ɘ�v.��{�p�ȸ�F�Ћ���DU�z36(���>|݊�3'�ow��h�":��e��"&(�3"�;{"�ݓ0^�\{M��X�'*�N�q�֬��}Q�G�1�+p;�+�euAt�t�+m�J��஝���,��.��3 ����;�X�E|���c�rU ������΅	*K�q�}\�/&.طb�;{"�Ҵ�즘�at�o0^�\ynŀv䋀N와J�%�t�t�$�5�'��XnH��ɘ��\;^�W���`7M�|XnH���f���@o��ذ9�L�n�uç�:z<#��SG6+Ga^n/&r��ù�I���h��X3M������l�]1ګ���?n�ـm���'W�XnH��[qJӻv�f�n���خLɝ��gtX~�{�3 !�]U/�6��&����X>���Y'gq'ga0��I�)�!�EX��hcNDj�V���!�*���!y3$�/��o��_7����ٹP��E�K�w���̓?�������1�6(9����9��wKû���;Ó(%�b��{6��cw���FwE�ے.�낅�WWwE��է���]I=B=sUh�&͖��5h�d��f�ur���SMݷh/�� �݋�w��/�]���tP�w]���u�]<ħA*"T�G�b�2I�D��~�3�~�36�;^����Heӡ�o��;rE�;��ݜ﻽J��FwE����u
I���E�mp�&`�9\|�b���*�@!B :�v���r�}%�!�v�P[t�y�n��p�\��@����p�&`r˭BU.��6���.5�ڻV#��vq�v���u�y�0^8��À�]T��6��m� �-ذܛ�n��L̗��Ԩ����B"ER�:�t�SUϻ�\���ou���\|�b�7�Gj��v�ڱ�i��d�wg+�o��XnH��4�즛�N�*�����$���&�?,�$\&ɘ��ZwVӫ�t���eP��ذ?/�?�~���������Tm������(]/-Ur2ܽ͹�H��ڢ�j�N���k��l�V����p�jh�$r�9.���!2՞��z-'*眽�۬����J=�m�i�M�]'rm�v0V�툡��te�9A��}�n�͍V�%E���ͷ"��v�b[r���s��j-�n�.C�6�u�nu��޸�v�ug�(78͔����.��F�us��2�����OF�}�{#]�1Ol֗�8��A�9�;u�����@��/["�9Υ���t����ܑp�&`�9\|�b�;�It���+�4��mp�&g����$n��Tlw~��Fk�����A1.�Ue�I7�}���7�v,�[/�d�3 !���_��m+.ۮ�k���=��8M�0�g+�d�q�)P�qةP�>q`��p�&`��W �-ذv���컻N�����㨹�ٴ�n��i�x7�!0H�d5��T����|��]�nһV7@�f�����;휮�[�`��p��*;)���Պ��{못�߸s� ��;A�/}��b��6t�/sv�&gI3��7�%մ��$�4�p	�O� �Àd�3 �r�v�[W����t�'Ł��������&BfFo_����������7�v,��J���SH�&p�&`��W �-ذ�\8����W��5y�݋�妶�K\�6�qZ ��=�{n,�z��KG����~�����]���2鯮�bo:�~�p	��k� ɲf Cat	T����H�n�z36,����f��{6�s$�d�I��{_��B*UK��$��,f�W����u�<�C��+��`���9L j
H�Li ��3x�.	�{F�4�6��Ÿ[�B`��Z�YXh]�DU�f�<�PD�,%k3�u������fG`�=���w�l	p	q�JsI,�������p�� �"b���zЗ�$�J2��a��l�6�͏VQ΢�*����'-V�#��,�b�b'h��#tI�v��h3[1Pڎ�Ā2;p�p��l�1�t�D��6�a��&68���V�\I	`��fe0�+$��Is����%��h����	N�4 ��bD;S��D���Q�D: USjЙ���$�7�2l�?R�=���`g�u�e��+�V���;�f�l�p�flX~fI��\P��].)��x&T�o0�g+�M[�`��p	�&~��OϿQ�8u��Ρ���QH=�ƹ-�z�m�ݣL�W��Z��.�'En�I:M7\j݋ �Àd�g��=�Ԩ�b��.(�t�ʙ����d�_�&I�����f�*236,�).�1:�l��bL�$��w�9T~d���g��,}�D:�bۦ�������dX|�_Uv���	
""m}�� <wĠm}1S�e�u�7VȰ�l��$�}���?�ϿC��)�k�{f�������}�5��v]��;�;g����K���m��}ۧϢM�@_��;���L�7�9\ul� ��ƕ���+T������&`휮��E�v-��7���즛�DÐ�ff��m*23v,�̓��7���wu���lL'y� �(��Tb�ض_ �f�������b��O L�����>��z��2e���sz���͛�	0���� I�0i  �a�=������2�i�KEUUUŶN ��-�Ӷ���)�ܛ����j�aB��/1�T���P�n��;p��ڦ���U�*a�vVf�ʯ�q۴%`ʹ��s����)��xm�kq����C���e�Y@������5=��$F(1�e��nx�ir����;�� [�v:���n�,L	-�u��"IvK���BH�ww��wg|�dQ�af��	��ie�ވ;v<��\mf[#���7!؍�Ya���ϥ�x����݁�ͥ@y�7g�L�8{�y�����A1#��eLL݁�ͥ@z�dxb�|�$� ���-�WHj��p^�ǀv-��3d��o�r�I.<�*8�0T����ǀv)/�f�3 �����ݏ ��ƕ	�Wi$�
�n�l�0ݜ������%�	�lV�Wm�m��Cn�)n]�=0�r���yy��&���G:����`\��t즛�CV*���wg+�z�v<���$�+p�{��O�z"A�P�T��[��U�{�o�UO�@��L!��	,M2?T�@}��vfm.��m\ubN����'ǀvG�$�wg+�z�v<�.�N�_��cL��L�7vr��wc�;�À{�.)B�t��ۦ��۳��93dn�O�{zx�/7v�u�4 x��Ǉ[�ݱ��T����݃]9xLv�8z���<M�Mi�b�ӏa���H�+�m����`}�:P��|��|᛽J�����y�A����'�<��.�$�۳��={��-�*v��I�!�&b���۰=�����������`v�E�'��G���ջt�o0n�W ���xod\7d�U��۰�ժ-7\����ܑp�ɘfm*�2�â�J�v�LD̢\�e��*s�r�}jw��c�X�WGp��g���7`�����������0��W ��v<�.�N�_��wi���3 �l�p߷c�;sb���S�wAm�m������nǀv���3�&`6�h��CV���AɒO��ޛ���@_�v�>Ik/�@�4+0P@�$&Ṋ$�__W�v�<�)	� !Be�q���p�ɘ�g+�v���m���}G°�3�g�^�5���ov�mI$�^&=RO�(x��n��CK���3ٽ�`g�iP?�v&d��?Oˀ~�ߟ�۴���դ�`휮�����ظ}�fv���W�"�@�t<B�>f��>c�̒I��f���Ԩ���bPD˄�L�����>}�p�d�ڶ_ ���ۗrZ'򿕲�N�w�f�[/�v��*�>��r���I�4J8�JF	�0M�X0��@C��!��c������߿�ߧ��杄��v�[A�i���Bt-�1��^zL����! FZ���\�D����X�z�&v탮^��1[����s��R��lv�;�v�*��:h���Z�9�ޑ��md��Fyn�O��0�,�����wT�l�cEe]�婤��8y9;H�s�i=��l�D�r��C�b�����r�R�f<]��Z�wVɚ:�[��*؛�m���4����Q���*xbB<O�˖i/��k��hqg�m��gOhwAm�m� �-��;}�ǀv)/�g}&`=��K�_ɴ�I� ���ؤ�����n���2M��r�'��L�s���;��3��0�_]ȧ���l��ylv�7b�Zj��۾&L�����v7�����l�lf�&��;nҦ��I&� �-��;}� �[/�w��0���pj�*���邝�n�QvFc���ݎ������e��h5@���C��Лn�N�T*.Ӿ��xb�|����o�������c�TU'���ﺾ.�%�K��w��`�%��}#�;r�K@�����Zw�;�I��l���xf�pmK�P��c��m���7�e��}#�;5Àw��0��K�_ɴ�I� ���<}'+�w��0E������;ꙉ|��v,%ƳZ�IK�4[�G=����)�eu@s맵S����ϛ;<�_9�q��9\��3 �[/�z���-�/��Zi����p�l��3^����ٰ3۴��&fw;;]�Z^e���ʈ���3�y�?�ݛ=i2Ȼ �!��6��!��1!�iX�F`D!�02�B��$�����J���۰1>�6f]�uE����z������;ٳ0E��{�*'���Ĺǀo��p�l��l���xݰ�W��X�:ݑ�]���lV��R�ܙ�=a�:���d����i#�;Z���i+�`����=��}� �I����J5L"It�2L�݁�׮L�I����s����۰=���xxh�J���\� �I���I�����n�])�J)�����ݥ@o�&`�K��/����͘�yli|&��+MUݤ�o�&`�K����'+�{޸(X�uwtYIݍ��ۘ���R��v���;[ttv'f�N4ut�
G���J�j��7����nzG�n����I����6��!�*.۾۞���r���f褾=���Lt
��b\��7d�p����I|�=#�=r�K@�����[u�7ޓ0E%��� ݓ��=�`�J�����m�褾۞ݛ3v������iS������F��p4D�h�8S�L-����~Z!**]2=9�F�@���bfh:�D�K2͚w@kvj�u��fa�B�{���E2�vu����a�ن!$����--�A�IkVXR�Z&ձ�*�i	H��G&X[,Ձ2��A�kA����5����BH`�6�@a��{p�5�2�NE�&a�0��f�0�{�!�Bcae�e@ݜ1�0c�&�z���v�{��p{��{��7V���e��u�zc�{H^ک�m   8@6ٶ�  ml    8���-�-�-��        	   -�� � T�t3�l�R�l�t6���M\���<�	����گ7Wi$�\g��'r�[�6Ɠ��zż��2l����.��ͻ�zQ��I�5([ ��sL�URk
���T�@��y���hJt�䠥Z�U�)��[`	v��R���2 [�s�jI��\���@Vvʰ��jtm��s��n��[�u��K7"޹�X��uK�&ڎ5X�ѴMyyV��v%
c[���� IӍ֝&ҭ]lZ�J/WT�n�s��U�Ԇzum�z��cU����]cBx5�N��v��Z�}f�����nI�D��E�\h1ͥ������tOA˗`� V;6%���t�l��I46c��R��(�t����hmz�tvk�z��VƬ�:��c�.#	w�׆���m@v��v�l�����Z���"���rl��\�4u�cun���zq�S��m���j��L�vӄ���nʵ�+e�<��]�XX*)bs�]��`766'�W!ĆثhĨA-��1�"�ގ����r�I���T�n�� �!�T2���iT�.۠���7blr�gb۷Iس'H�{Nk@�v�Eױ͚�H��� ���hb8�݇.���.Ål�;D����t��nwXv�e�p�U����:6�v�ңQT�&�D9���@������ti�'Q�k�4i�Y��w�Cvڭ�*.;V�=s���1l��۞u��B=�W	���N�J���%��7�윺���:�rg�����`8�ѵ:A#=�>�8�	[n��fܢ��D��u��a�[��t���cY��lA!ַ;�&��xSV�jvʹ�3��!-�gv�=�J\Lv %^���@W�{�����׻�AOP�U�U؋�pЂK�BJ�$�MnuS%�ܧU35S-L�oPn�-��q��Ŵg�I6���ѷ�F��li�VX�kQˎ�;`�Kv�\ݚt�:b8����\��QxGv�x��a㫝���3n�'lX�u��[d��;dn*�g���F�^1��g&&ꀼ��sm�
�m�۱t-ͫ��ۈz�뮡6۲�����'-ǜ����W6�a0\��q�]:���&鍸I�Rt�����������w��ߣ��R݋���k�m8�g���h�{���<�0`�t��\s;aǋTĭ|�WBn�}�<vNW �zm��/�3�����&.�R�
�U><�'+�o�&`�%���?�v{T���I��[j��u�&��ـ{T��;s�<�'+�OM����ĩ����y�{T��;s�<�'+�o�&`�V��ui��Qv���� �R�3�ݻ�Fk�ɾ�؃��y%�m���k3ƨ�l	{q��	�x6�l��0F���n�`����\�����@g��vތ�䒷?gt�����U���:Vn��e���HP`�aaF���M�8̙�=�Z���͛�fҠ=�[�t�ۺ�lv�`��|�=#�;휮����M/�����5`����ń��iP�n݇$�����v��Ճ�p�MT��]`��Ձۿ}�|�_ ��H�|\�����-5V���:�\�<������8CKs����DN|��Tɶ��Iݫ���'\}�3 ������l�p	��6��4տ�o0�l�۞����W �zL�6��ں�I�]�������l����e�a!	Xf��o����tP���b&\Dʋ���L̟7z����`|��̙����6�;�<�˴;C��*��zL�;{"��������utD���{��݋���,�N�m�� �5���=�O:�r.�.-n�h�ʽi�~ v�E�;s�<۳��7ޓ0Igxcb�f �����n��I2w3w�P��vϛ�@n��1t�"�4(������=�����n�I3;��z(?o�� �)_	;�R��]	:��I�Wy��k�w�y�����;P�j�����Ī�I��y�v�Ƞ92d�����<P�n݁����9î۱�Qj��ptvץ��m�;z��T��c:�v�դ�kT�<���2ˀv�x�\8��fۛ ��J��&�Ct�8���p����6.ؽ"�;�Ih��w�T��p����6.ؽ"�7���=�`�t;wWm����6.ؽ$X�(9�&}����4���Q����\ޏe��p��0�ظ���lR��������I ;m�.��8�	�ؐ�k][Id�ӫ��RYE��\ހ����a�z��:��جa)��[vn� �6��[���2�;9+M�m��s���OE�euϦ�O�_�p��%1ӊ�n�T��I��n;s��>݃b�K�Z9⧱��
iu����'9����s;�/n:	tl9��L�Ƹ�&�Ѯ���	)��l7$�Dê�T t�q2=�Z܎ݳqq���J�rX�)0�t�ٹ������1��B��檞�����ۻvϹ��{��|�i|$��J�Ut&���3 �͋�{ޜ���+ꪫ�{9ۥ�bH�0��7`y�z({�ZX�p��0�"�t�ӪHUbMp{Ӑ�7���;�&`��p	�/�@�	��K��`�_%���6.�zr��I˰�k�MYѦ-a'�I�zm/n�8�]����l�R�6Pĝ���e+�5IZg �vL�;sb���!�o�À{��J0E�˸�$<��>��Z\ڼ�>HC!�LRRP`h�fܚt�	���0�)�` �i6&jȴ��X�w����l, ��X��I;B���4Na��<Q���~�U~���\��v��$�w���'�D�Afuq`g�t��fL���w]����7})L�p+�*T���8`�p��0�ظo�G�o��/�݂�i��g ��&`��p�d� �k�}��}����n��U�G2�ny�E��W����"=�κ�p��%�(�z�/+V�i��;sb������zL�6�J\m]+��*�&�o�G�o�Àn와v���7�%D�wEB&T[�T��(�ݻ%bf���.�4�8DSD�i4f
I��!2J�2U���P>�6l�F����$D
&CĔ�&O���X~ފ�$� �k� �mD�[�N�n�7�nl\�$� �k� ��3 ���~}��c��G8�b��H�n�l����hÆ����Z������q��\��HI5�;rH���pݓ?W�W�v����@n��\R��T�/SSS`g�t��$�n�U���>|̊���i|&1R��]	��{ߤ��6.ےG�o�r�}��B�UwM5n��O,�sb���wf��fҠ�d�N̘J".�Jy��{ �������%*��k�v��휮��fۛ ����L}�n�c֖��je��&^�ɶrn�!*;��YҦN9}}��Kt���b��C�Z������&`��pܒ<�����"�T��\wd��6.ےG�o�r��j%"���mݦ� �͋�v��휮��f i!]��R(m!$� ��#�7�9\wd��6.�5L\�Uϒ������W ��3 �͋�v��k�[t!��V�n۫۫� �޾ HN�����ڶ�.�KF���[�6m*YML����Kk�oN��ZG<�=��b'���f�C�2̇iv��:�;k�j���g'3ܗ�"��5q�ι�8+�e���ې,S���sp-�͹�X]���ۧ��c\qˑ-jWY��O�ג5�2�v:��Ĵ��\u��)�6ܹ��k�ػh �8���8�A��{Vڻ���+�>�n�O&��n��Эgw>���4������7ϔ�Żi��i}�B�i��u�?����fۛ ��#�7�9\���!M�iU�v���y�v���;rH���W ��3 ��)q�t�2ЪĚ��$x�g+�n와v���7�%D�Vڢ���\��7�9\wd��6.�RE��#E��Rj���zn��;sb��$X�g+�N��쉦�[w��+�bh�I�x�Ɍ��0�W�[]��8�%B���E���ۻI�ۛ ީ"�7�9\�vf i!]��#ᴄ�\�����k�i�̐��8&!$ʤ��v�m_I2kr�6��6��sb��݊yRW>H;g8����W �ݙ�v���3T�`^R4��Zj���pn���6.��� �l�p�颙�1	���;��݁��lP�2o�{�>sz���۰93,�O�Y0�!;�����v:��U<S6���{6��8���b��uiC�R���t8�,��߿����X�g+�{wf`��p�	Q:���Ct�8���W ����;sb����|��ɝ��wL�q�@�aD<ʠ3wz��sb�Q�x�d��:f@�3U��c�R�8�	m�&��LF�#��: �� 4���# �p3.�]" �AD�V�� @�t�[�a�f&�h^u]3�̌c4��]�N��s��t� �É1b�2	�$�	"�A`���"R+ �YT���;��a�P��ѭk�1t��\s ��I�t;N( ���/ >"��t�|
�b����`+*�(`��}��]s�uW~}�U��)���n�'�nl\5I�����٘���v�%��m!$� �RE�o�r��vfۛ ����w�3��n̈́��kRZ$�3��c{D������}��ϫ<�.����.��Ϝ|X�g+�{wf`��p�$Xה�/��*V���'\ۻ3 �͋�f�"�7�9\���B�TҫV��ݶ� �͋�f�"�7�9\ۻ3 ��)q�t�Ք�V$� �RE�o�r��vf�U_nl\{TN�m��eC�UE��ͥ@rl����<���j�,۶���-�Ae+e
ֺ�M��e�q�-`p;9N��6���l��v�$q�����H��%m� ����;sb��H���W ��%R-�7wVݼD݁��lW$�2w>���77�P�٘���v�%��m!$� �RE�o�r��vfۛ ݑr�0���@��>q�`휮�ݙ�v���2k���)_	�T�5WBN��v]���lP�;�`g�iP��J�%h@b0��$��X�� �X1 b���{�fZ���>_�9٫���Wcq�U@�Bt/M�ۍ��l�jۗ�szWM�ͣb.k��qm�<�C��&�S:�`���P�LG�ʵ\�K�p��rr���7L=\i4C��q�ѷGc�	֜��l�#e�e�wE�[��v��[Y\��E���ɷ]<&���ۊx��s�88��[a�-���9�:܏S�>b�����Z햶��E�����o7f�m��V��"x_��6��=��q[���&�fX���K�j�l������/�ͥ;!��OK�V�ƛ�\� ɮK�7�9\}�f��.6��n��h��&�f�/ �l�p�ɘnl\{BTN�cvS���9x�g+�Ol��v���'��x�4Pݟ?�������&`��p	�r^�����F���v14�y�v>=�K�'��p	�0��u�J�Һn鴘[��ՒW�qͽ��p8ƶ�<�f^:]f�ᝰ����Kᴒ�� ��%��r��ɟϩ�7�n��ݱO*A���	u3SY�_y��9�ЖV��`����i��`H��LH���`�٠>ܝ׾d�����w��1R�l�g �?~� ����r^ݎ���B�TҫV7@�y�ə�'|��=�=�`}�:P�ݻz��m_ɢ�v��Zo�vk���p��0۱�M�"�;�v���Xa�5F��Xݚ8�s���q�5�g��d	�5�m�:iЬn�t7J�9��;�Àg�v�ٛ<��+p�l�=�Ϝt��q�����D�{7n�2I�3w���l�=��l�\�$�foDt���Ze�H���� �ޚ���{)5�$�$��2I%)%/�:P��v����!��w����d̓��������@g�v�9�3;��M����h���Q����p��&`�c��݋ ���������;o�`�7�ыQ�\ȩ��^�p=¼Y��{m�V���Ūo5��=#��%��wu��6hz369�$�p���@g�۸�aLÐ(%�n�=��\�̝����=�<P�ݻ|��m_ɢ���Zo�{�v,�8zI�����	Q:��N��UQ`}�:P�ݻ �f��d�I 0JA0Rĥ2I ���w�b��.4Pݔ�Bj�I�=$� ��|�[�`���=�ut}]��/u�[��E��K1ӝ^��Y�vY(竉�y�1SJ;LT�d�m�k2՘�����2��p��&`ˈ�P�%�ڻI��n̬�8zI�������������O��wc� �I3 =� ��fV>��w�h��%l�[g �M��ݎ��ٛjÙ�������n�L!@7@��n��=�ٕ�wd�p�߿����~?_�@<�(]/-Mե�{�s���m警k��`臛%�W��Ym�&VZ����lB�:����a��ܶ�z۱]e�9J��ݵ�V猚q��cK��2u���L)!�G��:�Kf�:�[��;nsj'26�)�Z�r獜D�uv��@R=ЛV;==�h��q��[Gd���>�9;|�bۃ^��ͻV��n;����<�{���v�#�.�`��qE;]�� �e�x�ľ��� �X��ݗl<�&�*O3�٫��������윮��3 =� ����Xݔ�n����;�r�zl� ��|�ݙX�iq�������Xۮ��3 ;� �wfV������F+��Rv14������;�ٕ�wvr�{�f lԮ­B���j�&���2���W ��3 ;� ･�`��V_ɺCe�w����{nn.;�B��[%l���u����]v+���!�ؓ�`ݜ���f wv?ɓ[��oZ�9�7��x&\""U{�ۿ�&fe-�2Lҙ�
�٠7ٳ+ �r���
mSB��6�`�͚=��Vs2I�ٽJ��������J�m]�W+M���e`��W �eɘ�l|{ī���n�t7M�yX}���2zL��c��l��o���8��kl�>��nӚV�۪��uS����w�7/��2�A�2Zq���yUnۮ��f w� �{fT��{c���Q���'n���y�����nV�l�p��0�R,�P�%S�n�������Y��"!$D$LE(Д�����2�32iw�߮�=��@n�b�T��.��ݫO��w�9\'�f w۳Aɒf}�o|�l��v	�S.����٘�l|{�2��g+�~~���Q��{:���c7.�"��1
�10�[��t�ól&nZ<ާ�>zt;i� w� ��̬������0	4di]1�e]��7�'�L��v{7�P��v��f��x�#fIre9(�S33j��ٴ�o�v���ɝ�f����j�=�fD��h"a<�ʠ7ۻv��f����V��3`��$&	 d�cH:��~���5/�W��cCO0���ݓ+ �r���0�K��v���7l\\U�-��i�\8M�k�j�sچ�����v%�mn_jAk����X}���'������6z޺t[%ӰC����`��W ��f w� ��e`�-���7ai��OI3 ;폀M�2��\8���>mS��T����c�vL���҃�L��;���I:bE1"aݕ��ݓ+ �ÀOI3 ;폀vl�=���L�)�013l&)fH���3[##cD�ش۳C��n04��4�N`N�X؜�7kv�,ػwa�E��'@C���2C�u��y��:C�ȱ�LFl�Y��tlȜC�֕-�y�l]�4Fbj0���tM�ň��̧�X'� S4F��	��Ye6�4=%�HR��'����'��0p���:��i)$N��\l��I!��ZH!���7cRq��=߾9�������l�˒T�B��b�Z]�j�)Y���   �m�m�  �6���   ����pm����m�8        @  d�  ��˴�i�.]��ó ���.�J�
��:ڵp.����/����%����q�9�4�J=.yz7񌖎d��'%�\�1�d�b�=F)��H� 壅eWV6m]�%ej�lJ��s+/-*cs��e�z;[#6��i���H6��n h0N�b�m$��.XY������;�jtmmJ��K��]`u��.:�^�I�W�%������`�P����t� ��SMwK&�-ܺ�VE�����lKn�j�Nvl#۪��3ۅlGW�<��c:��e�;R���G[tգnC$���z5v�gs�������g�����Lk=m�dv����[�� Uv�(��6;t;��Ŵd����,n�'��-�=�=�����pQ�&���]RdUz)淡vNâ�d�<i!7;kZ�Yq�eN{z.�rp���v�痞zv�mU�p������&��)WF��v��\)�<5�P�H�"�A������8zڍ�[G�nኁ@rָ�b%�`�m]��k�M����i�vA�݌�vp!�3�Zo��p��W��N�\�Q�l�c�e`�Ep&��.n��wC�n.����o�|�����z�<�s/H%�����Z�|qZ�3<e=�l��Q���uV�؇=�7Rd%������{z)i6:���a;AЋ�qAn��Ԝ\ktwI-�m�/���/"�o�u7��]m �a67=ӪnH[qŭ1�k"f���$Ĕ���݇��6�F��-,�ζ��$x���ntk]���`���B�6�Rw\&-�4��#L�_n̺���hŶ�s�����Dצ�&� 1e�ۤxg��u�jѵ�g�N7T�]�uՖZP]�A(:�ni��ꃶ'S��sld[���J������{���t��
?��S����aN
�
���x*;�;�F�c�V�,�m �����$'Amv�j�]V^���gn����6��S���N2�ލC�F��ڠ
W%��9b�g&��z`�a��Qh�=�����y�,�TzXF�m�K<p�q�벩i�A� ��%���sAn �n@7A�ݓ�*��=�Wt�ۧ���u���,�9���>vy[�K����Q���5\�X��[�3<-�ڶ��{���{���������L~�ѻ!��-�:��3P�U�;6��O(���O6�r��F���,,�Ct�o�]���p	�&`}��	�&V {�w�'wO䭪N�8�٘�l|o���;�p�=�W����16� ;폀M��X}�zl� �jWt)/���M�	��+ �ÀOM�����6m�t�K�`�we���;�p��f`}��	��+ ���D$�ϛ���R��Wg��/v�8ؓUg����)��n�u�}-;�M�Zl�?o��0����Ik�_8{6x�;5�y�aJ�hS�x����4&L�s۶������۾d�$��g):`�u1	�aݡ�f����V}�zl� �>��B����Ct�o+ �ÀOM�������$��;�V���."%�AD<x����3 ;폀M��X}����3c�qG�f�4q�r�@���nTuX{
Z�۳�x4r٘�Z�����O0����I��w���'���	��w��vR_������+ �Àg�6��f�s33;����K���iX͞(��ݟ�Jm�ɒN�@�	LM	�Cꋥ��dA�q!�S@A�@)���{�@_vm�[њ����pt��7�f`}��	��+�_}�� ���B�T�WJ��ݧ��l|��gw��=����sn��b}"��Q	��707;U�֮uD�0�n,[�5�zc�`\�-v�եs��Yy�C��ͷ���߿��;���٘�l|wb��bwt�ۦ�yX|�_ ��3 ;폀M��X��ҷ`&��%mRi;��f`}��	��+ ���=�W��6�bm� w� ��2��{�r�CY�

(BR�d|��E&��!HS�CB	��>�������k0�Ϸ�ޛm]�� ��2��l�=$� �>m���Ӿ���':Q�6�Y�I!���żkH�݋��$��z�:�g��W]�n�m���m��l�=$� �>7d��%yl��Ze5V��m� ��f w� ��e`��|l��)�N���%�f��f����Vs$��������0	�L�	��]��7�'��X|�_ ��f w� ��BR��N�;t�7��w�e�	�&`}��	�&V=��WI�����}����n�[|8 ��אB���s[g^t�UJ�'���B��]�c�tL�ի��9u`,\�捊�7l(�0�@6���s��W;LW���K�'v]��p�%���L�����y�P�N�VQ�-a%g�=��}y�v��i$������.�<	�V�g��K�I��p�p���r].j��i��f�BVۧ��N����ި�7[�c�r۲s]�b^J��ќ������np��R2C���b'����ڧI[T�N��?~� �>���_�L��do=�n�t���e� j�y����7�L��[/�zl��MJ즾Wi7�7�L��[/�zl�����$��t�%ǘ�Vތנ=��v�f�3&g���#��H�"�O
e��e�nn̙݁��w�����V��@^���6��=��q[�\qB5.�����ѫ]3���N�����$�ԇ����'==�O0����I�[/�zI3 ��������s0۪�:{ﾬ����S$�SU���۹�`fl��lm��;�t����ǀwV���L��32w=��@k�wM�g�b\�yxR�-�M'|�I�������[/�d�J1_��M!��� ;� ���6��t��7��������u�Dw��e�	q�n�=�������qK��M���=>����n���A��>ղ�ͷ�G�wV���L����$����l*0;�>s �=�L�����'0���!e�ڦ��wʼ��몮�������$"3p̓2�I2�>ݭ�27^��/c��-S�]*j�4� ;� 3vN`ղ�wvf=)��;���M]��7��ݫ�&d�����w��>�l������r�+k��gQ��Xa�5F��Xݪ���pvuv���gl�T�p�ј:R����=�<Pff݀}���d�����`����۵Mj����ݙ����2�dx}�n��`���wI�7��l|/vG�w���;��0i#wue�e5@�$��2g�7{���l�@}��v	�$������>7��E���@�q�q��N�ٙ�`{6h|�ٰ9$ɷ��Ͷ����7�ы0;vz���L>E�]�|tmͮ^t:����X�6��&��Oـ���2�dx|�_ �{n�ڧj�7@�y����2�dx|�_ ����'�24't��؋�Zo�e����l��ݙ����'���A����ӷ�q><���}�;����2��<%ٻ8��۵N���4����� �> n��wϋSQ���m��M�T��L�!.�oPn�l�� Hp�ە���VnJ#�6nI[$�DG�,���w�X���c���731f����nm@�z���u�tt/�nx{�C�c��
n�l�{I�^s���+/��%B�įK�s�%��h��v.�fm��9�N�<m����>�s��֝��h���}��˃�xb�k���W.�PN��2��7W:����U4
���5��e��[����i�C	ɝ^ܼۢ�*�9J�y�n�]�*	R���n��i]�� ��π�>��Ӏwwf`�F����E5@�DL�f��̗���������͚�2L���~�R��G ������=�<p��� �> n���ym���c�T���8��3 ;폀�>��Ӏm{n��e�V��m� w� 7�>��Ӏw}�0Q{b�T�:I*�ܽJi:�9,h�[�6�n4�IךA�nL�ݗ�7H�js/�8�5��"`s:�p�Ӝ ��_ �{Uڃ�NiT��uu�{z�.�(R�D
D��l� ���������n��%mRv��;�٘�l| �H�w�N&��`����CV�� �> o�|;� ��f`�F���N�j��I� o�|;� ��f`}��{�\
iYut_ɺCe�v4�ۚ�����5��.���9�f�46�\��@W]�ny@��-q��[/�w}�0���������GŲ�v��|�홀����gW��׶�aM�ZnZ�ASU����;~��Ԧ�!��z! �V9�1]�õ���@��$�	!$M$`����;�L��fXX��bP�A�|a�%�M��0D�FS�KB�RId�ȌJJ�eDV9�H�G}�:D��ޠ+��Vm!M����Zٴ^m	l(,3���É���:$(�GA�[h�h�4h#$�4X:B0�α-A`����"�#+�M��7�sf����l�n���[���'&-!��4�h�a&�Ĉ�LcҦ́	ºځ �Q  ���[�j�I�F�hI$��hh�����`0%#(�gN$3Y�a�0#8�;�C4&](�'��j�*���/�!����_z<Aμ:�A}C���� ��f`ҙ�i}lE��&h9�s�h��@}�λ �ٳ@nz+�*��ӧn������|�홀����ok�W���|ƣ:4��pi��ƒuۯE�!�qA���X�뚐-��բ�CB��w�;�٘�l� �n��p�њ�v�~��yA��5m<��c��G�3��|�홀I��-;���I� o�|:���;�٘o� �׼t�L)JTͷuX���`{���ӽ����@!C�� �*�=wU��FF�<�K�(L̽�{:��ٱ@�٠/��=ə����
Σ��Y���&3p���T�pm)�9���N��y��ٰ;1����M�Q����<���ݚ���������?V��~hNݢ��]"�\ �H�w�N����;~ظ�!v��V��t��q><������;~ظ������n��&���3�w}�0߶. o�|;� �kn0[�[��i������g|���l�+���6,�ڧi1�m'vۦ�L��kn�s���[B���4���N�t9)tYԸ�sp�Xv�@Ex9U��=���&�w���5����u��\��`��l�5�f���L�h�f�^(8�GN��k=�p�7�U��9�����a�ZwM����n�H�g͝��l*��u�h�|ڴ�k�7]q����qG���т-��3�������:ќ6;���.ظ��3kF�n�n:@����kq�4������A�rHNL�"c���/�N�����3|����;���J&@�A��EL���p�f�����mu{K>�Wc�T���8w�3 ��b��G�3�zp�m�L�I!0��o� 7�>��Ӏw}�0	^��Н�E5H�E������홀v��p�e�.N����'�:����z�nͺ�y��G���Kf�OG�7;*]�1U���;u�O� �Àw}�0�ٱ���n�t�����Q0=��kw*��=��[T:EU0PMa����	7_ ����$�ی��yx&bn�����ݚ92fg�����`�F���N�*��k�� ����;�٘o� �׼t�N�J;�%���\8w�3 ��b��G�;�;/�BN�ۿ�j�
�溸�ĩ�{���uK�9��=�����[�������v;�H(i� ���0߶. o�|;� ���l)�N�ZB`6�`�l\ ݑ���3 ��F��1R"�\ ݑ�j��VP �� ��&ja��BY$�BP�I���$Ib�� ���|ǻ�0��p�A%Zj�7�uS`}�(�3n�����2I�������ؕ��4�6X�'i����0߶. n��w�N���#3c�qkq�n�GW,h��[&�GU�`K]�\��Ŝmvb#�䭯�b���`�r��#��=8wvf�"n�ǉrHNL���@��\ɓ;�{'N�'��;휮'�qӡ:(����;�p��٘}���� �﷗Uv��v�-���ݙ�w�8r��~�|��v��J)�G�o8k��~)�N�ZB`6�`��W =�>��Ӏwwf`ݫ����x�����֞t����K�Q3��т8��E�GV�8Rڵ�.y�cvG�3�zp���������%Zj�;u��ǀw���;��0�g+��> w�ԭա�I�Ʃ;L��٘}���� ����&�m��-1$��7a̒d���T��4w�N�����T��Ֆ��Uct�u�� ����;��0�g+�{��~?>�We Z+���
��[|8 ����l�!'I�Dݤ���i���V� :�v��(դ^�-��,�͇F�K�H��H��]v3�|�\j��M��g�x��2µ�R�m�=��]v�/D�V�y���h��ѩ�gq�N��z�
��~5,ə��qӫhӝ'c[Epb�Mu�^L�M�95�xF5�,�p,n��г�^ն���{׽�����|r�i9�[�a.5�Ԓ[�,tx�,�u����+g��U�ۧ<���݅�;�Z�~��wwf`��W 7d|j��WUv+�*�E���;��0�g+��>��Ӏz��[
mS�V��	��}���� ����;�٘���67e�uhT�7\�|�'|��>�N����>�m*�D�LUi�`��_�k� �f`��Հo}�X�!�+4JS2�Nk��)�n}	�Y1�\�f�l�K�i#v{Q3�m�n��&���3�w۳0�g+�� ����&�m��N�LK3{못�߸sj"�*�@u^���ʻ����ݙ�z�H��Yi��V7I7\ ���w�N�n��;휮'�T�DJ�K�<T͇32I?�k��'��;휮����6���]�튬 y������v2L��zՁ���3�zp�ۊ+
�WwAwIݍ�[n����K�۲>v�����S���S���R�mԩ�+HL�������l\;� ��f`�6X�ݖ�աR��p߶.��Ӏg}�0�g+�w�	(�j]9����ݼ���`g���=	%�%$% E � |O�T�_�j�������ҖT��N^$�/�f݁��iP?�b���3��(�\�!-0(���"�n��ٴ�߶.��Ӏg}�0�t]D%R�[�Dݛ��蛵,
qn���+��Z6y��]��K���:�8�q�k�m�g�����=8w�3 �ÀI�t�N�r��ˮZ��;�p��٘}�g{�`r�o�A��Ԃ)�{�f�k� ��b��=8k���Sj�Ҵ��v�`��p_�.��Ӆ����AL�C`�62�E$��˽�f�,DD�o1K6�{ى�R6`N@`�8��.�aN"�K:d�k2f2#o����̓.<˩Li�tX;�;=�Ł���0oT8IHn�A�t�L��5ƫ�.�i���=k�:��3Ӓ�v8��l�k�i0v�b��k� ����;�p�;�; ����R�L�$m:�E���۾fI2gsٳ����@_ޜ+Y&Og����?�);M16����K���3�zp�f�"wue�V�U�*"$��də�3z(����{:�93&f��<�C�!�8�GT�Q`}�(�L�}����͎$��dP�?����?�0?�����"����E?��������TD�QUs�4� +�� ,B"�R�(k�������?�@k����_��}����������ߛ�����Z��_���οg��?7�~��_�x����Q������?�����
*�@
*�����C���?�������W���?���?�����?�������?�����/��?��?�����1P�""���BH� @)(,��+*$ J�(�B0�@������
J	
$�����0�JʉB�	 �,���(���*$�B�((��ʉ
�*�"
$ ��H	*$ʉ(2�@���H)
��H����"�
��B����J�*$�(B� �$���(*$"0�@� $"�@�� HJ� ���� $��"��HH,���!!���(�J��B��@@�!�!
���*0���!"@J���!
�H�*�*2
H�HB�!# B$��H
2��@H$�(�"�
����H J�@B! B�! ���!2��"B�@@) J� H� B�! �� �� ��"�� B!(0"��H@! B� J�H� 2� �� B�*B�JBH0�!) @�!(@�J��
��
	(� H�H+H$
2��H$!"�H���"���B2��*B��J2��J0�,@L�$!+(�H2����� Ҩ�H	 ���Ҡ(����?���TEU������������P�O�z������y����������� 
*��G�������aW�� (���B?׾H
*�����U_������kgF{�a��6~sw��ٰV����������
*��z������o���#���� QU���������q�?��Feџ��?��<�����ه�������xi'�h���o�~��>�@W�F��O6 ��������͟�����R�����d�MeGӀk9f�A@��̟\�۾ �R�*"�   DP��D�� $      J(�! @R�� ��EU)D �RE*�E) 
U ��*TR�� ���J  �  �  P  C, i�	=}�U�5���@�D�{�he�L�Ou ������T7��o����}���q5��A�. =�V ��
�f��s�}  ���	  @E#�P �,�  g� \@ "  �  L� "�1  D
   @   "P    Q�� � �  � � @ x`(`R�� D� { ); ��0�@  P �U� �� D  ����ŅYjK���������ʾ�>�����zyr��P �Jc};�l� ��{nCS� �m�şF�t�m��Nw� =�L���}�v^6ON@o�<      ��  ��c\G�.}����� gA�x�r����N /� ����fx Ðzd�;� }�K�}���o=�*�qL�PM۽�NL���q��ˢ��_ �*T �  ŨG��3Jd��wO ��yu �Ku��{�}�|X����
9�3��r7�  �Ou�X�@�o_p�{x�{n ���ӓ���}ڸ�{�<�Q�    ����R��� ���MR���2`���R�ڔ��  =���(� �*����کJ�� �")���P�<SR�����?ʏ�O�������;[��TD(J!_����* ���
*��TAU��TAU��QV(�����	�ȁ3��SC:�ba��b��"�_�@��X!���aC"V-�I�H� H��A��	1�Y��Is5��+H���%$xp�]A�d�|5�_��"X	�5 E�$#<�of�6q�BB(Q"!O~���=��"�$Ѧ�
HG �J���$R>����4`4����6W�r��������g���X�+B�`D���QiwbA�S��`Qs���cĄ��1jd\8$�"�GA�r�ܺ޵6�4�P��-m�+2D���p�a2��r� �$�͞���K��T��������'�R������Y�	t��n�!��j�$��r?|��J[,'�]�#(a���n��eʐ�錑�����G�B'�
�� A�QHD�(\2y��3�>�m��l�ǚ=1��5�'=a�"�h�E�K �2H��8�I$M��E����w�.���yr�.q�ժD��������k�7xx��k���>!	N�+7U�fi�~�0D�Uxjr��T�z��^w�/t�ʴ�S.�Ϋ�>����́ �"he�'0��8���%
�"�)�W%)����s.�4<0��h>>a�Z0����	�0��	�H
���ѣ`WFh!��F�foZ'9���':H�	$��!���|�5a_��m�t�sy|��3y�����#T��RM.��+Ƈ>��"�KcuU��Ò�J�b��b�K�t&�g	�#�!HGQ(I��/��R����J�j{�AS��e��@�7�m�uf���/<�Ȋ�&�Uc���W{7���*eO�W��Sy���H54a�%4���᎔��@�dd"B_��$�A4�� DH5�7ǵhi���8/"���C�PU�UlHˣ6c���,�Ha�\�4a���.&(ka��p̈́)�6a����	����!��qDj��;՞�Ku����E!V=��`/��g0��0߆g��-��� SD]�2�4��H�aM�)$� ����7��{����L�Mj�\�# F%PԐ�$K"b�]BnL�Ǜ�3��`��0��"�Fl�|<�O��(��9��Wv������'�=H�1��op�\1Ws��]	Nm��]M� �wUs�^n̳=�2��;2�ڝ�Wu9��0��x�^��ԿM�jbT
W����)V��b�sZ�o����/�)��{B E$d�&�l�L]��JD�M#q7������$�oG1���:p6@����!�����X�y�#4xڄk��U��+�VXk\�5�8i�ֳw�ɣx�ķ~��f�/��i`mB�:ws:�	);ؾ�HS�`����9iB��ލ�r]2�͐�0�p��o7�Y��jh1pa���.�M�7��B��@�E�`@J,
?���$����"B�ћ9���ӛ�<�@���L�6s�ĺ0�6W��U�B8�A�����%�12H-�4� B � �H�4h�E���HR(A�A5)@ D�$+�	�@���"HQ�5/�3|�y	�ԊH����0�O��X�`����F)H�b�DZ$
�Pֺq�B4�4�_X�%5L�/��HB�0���H@����琦$�0��6�
h�@��p���4D���ma��#��SϹ~�NF(P~C� 0��%t亥��*�׾L̾���0��`A"� ���F��5�ik8�����Ԣ)��;��I�9�nj􈛫��ɻ̨����n�f��a9*���QԜw�!GA�ț]B�1ٲk^y��;V%H��s����g�Xny}9/��9�7�������MU���(�q�?Zb�!Kt�u,���:W�&��C��*��DZ��j�(BP%4a�7R. 6@�,��J�tc��D�	�,B�
A��$LN)�0" ����	����/Rh�*����˓[���F�~zm�x�+���y��tl<� �qv�U�j�.L��y��R$!��ō�ng8j�>x�1
la���y��s�h7��p<J]�`����l�7R�ӻ���{��6�N:r��^%v�(�1 Q5h�w6� K�.�o�\ٹ�G�9�x�
I�Ѭ�8xC4���h�fȄk�5L��s7�p亙�r�ɇp�DKUuy������L9��N,�ymg{}�ɺ�*Q��Q�*�izĵV�^ۗ'�"R ��T]<^�b�\�Ժ#3�Hy��~�E�8zY�#FR&�R,!�!I�:F:f��0$%tC2n@�42���D�����~}|����V@�X�hA���`cf����0! э!���Q����+�~&n.Ƥ'�b���Ͼ��٩鿰�
�Xf$O���L�R�x^*KQc���HA��ɷ���rDK�W�^ʧYr(	N�&e���jVb5D���Z��x���MD9��s�<���ĺ��j�����l<!8a�~ks�����_0��ʲ�˩%b� R)T�"�E�ƚ��3�!u�ɽn��q�ц6�j��
Eus�ljD)��WyTK���Pz�s�zɘ0� d�����`Mp��{���t��=�g�
B�g���3�u�4�)�A���>!��q���ux}��$
q�����0��>�
l��������Jd�d�)\M����)��#5Tl$KUh3��O�b�Vy{<����M�T5u/	p�ɮ�œfm'>����H���)^m�C���M���YZ]�N�-3|�ZS�K���N�f�k�iŊj̥����mκ�-�gB%�V�s|�L�F��"j��Y���g�'�'Sy�|42�+h�U*c�
K�oӛ9�)�sG��y���xF��w�s��諣FW�!���6$�1T�sس-mQ�3�ݝ��*���qn-�KOח��֭5yB����uN��q��[����f�nB�B����9�P��sA�]Z\6Q���aH�����3����2�FO��tK'ׂ���bj��R��	Mҙ�֐��VL����.�缅)�k6��\"US�W��{6ZD����y�����uc�䈔�-b{�[��! �G�Y��/<���x$���y��y
c�RE����4G̞�.x=ܻ��;J��U��s���˂�B̸����o	)��|�r�A �c�@�5�M5XҚ�v���a�u�F�4ю��ssO$�WD�[�o��������5�ns��<v��3{�77��D�l�4T��ꑚ�1R$�X����v�,a$� �J�d�1 �@�P�B)�TѨq1V��$נ�%	�H�4�hў��H�2<��H��@JA����/���ʣ$q�M�T�f& �{����6A�t����4D�k9f�
{�箈@b�P�!aY����/!�$?!J�����嶧��;�T�#X�v�r%p���	@|�٩A�	|5��`�D��ַ�`iMDSD5
�(A�!#ʗC!&���
Ms��5��B2�sF�S[�4hӉ���e�!��փ��%�aC[#MB��],*�#�2J��d�t��+�4Dji��H��h!D��A��SP`HD!
B�!��B��i�I (�XId�AaM$*ă�bD5�FM�+Ԟh����4���#M&�ڗa!�	��M��CQ�ѥ��۹'�Z@=
]����Bā�E�@qOt������������          l                  ���                 �   p                      [F� �    �`     �   �                p       -�                             ����    -�      �                                 -� 8 ��  ��              	$    p � �m�Ԁ m�m�YBj[�,�l  -v�k[m�H6����i��m��l�R[M�8d�pʸ�N����Ͱ-�m��[[v���@ݶs٧\v�����Wep۵`�u/Ϟ���י�n�Fշ8HIm
Kz$-�F˭m�r�Y�c���J��J�j�m��lm� �0Y� m�$�/�پ/PW:� ��t+Ur��R��Pv�[C��Zl[@	 -�l(��$  jV 8  �Y�q��-�P��UͶ8m�6ٶ�Zl�+Uv��Uj�4�ڮ���iV^�U�o�UVSV���]8�0&�j��+�#kZ
��&�ɻtulضSt<8 *��N��[���Qֹ�YR^�m�   ��I��$6� �;� 5�kn�%�@l�]3t �p�����J���Pm��˲��u�*��[[l/[m$9��  n� l�L�p�A�m��q                          $           �֓l    -�� �t�    8   *NM�@UuUO,���k�cI>�}��t�mk  �m����z�	e)m�9��l��� �p� 6�6�Y����m��-�� m�l sk5-��*��m�u��r���UR� S+Uʠm$ֲ�m ې���]w�$qJh��E�6�V� [���n�E�m��| ְ�sW��[�@p��n�eH9��B��,�1uJ�bz��*۵2���t��p&��W�������vF �S�G�uU�$*q�d����n�c�H��Ӏ�*U�;�[]u[R�m&Ŵ$�e۶6�$��-Q�����U*���������q��6��@V�˲��3U�Y�p�R�K��i ����wL���-�i6^.p�vl��+j�j��[Hp �i�d 
R�g]�X7f�����q���nT S�j�!�F�t��a6�]�dzݳ��
媫� � S�^pSR�y�:�S��iCW78ݮѥ�vj�m� I�ےE��(��
�զ�sn��s��l�շ sm�b�6Ͱ � ����AX43x�6
�� ��3���`  �M��q�_D�+��s�  �hXk���ꪠ����@[!5=l�75�<q�h�-*�na6j��{[V�j-P[�m��m.^��ڱk)h����#t[!&��%����	��3I��`�J۷�e��X��25T�J��M���wϝ��m�E�^�m�    l ���c�Ue�m�������� 6� 6٭���ZMUm-�%�� "6��gk#��ٶ;`B�B�+%��;/��!��l����n��C*�y�Z
N릭�6����u�v��"��᪠�Se,���:x����s�ѱ͹V������xQ�Cg���]k��v3K�şM9wc��\�0���]c���2cXf�*�t2���Q����ꮼ!�O*���e�%UW*���p�2�5U�&�|�5[� �� �6ݭ���޸�km����O�����-򪶨\5dmtG-�� ��$6ذ��M>���]d�m l� ;E.�K( ��-��ӗ���s�� �UU\6�ܛĲ��[kd���CI���m�mW�������¶j���Ŵ-�n����� m��Y�K���hI�����ݮS�jQ���c�6��u*���U�qʁ!�Mn�l5V��$�l�M]Ӷm[ �6�m�$��I�\�Zku��6������u]tv�ۛb���IH�  ��ݷ� d���8��`�b����+��l�͙�� r�e�N��@�N�k�
�6=�*�y`.��gc^Y�Ucv6^�\�h��W��D��3)-UV�F�-ܼ��4mg�j`�Z��Y/-��:I�H�4u㨐�r�,�݆�T����	�*�O#�u�v�j��^D�%�I�r 8�U]u�۵J�ۖ�� �`m����e��
U��*��U^n��he�v��a���j (��NRF���	�rPr�:
�j�`����l�wl��35j�����n��a�	 �s��6����"YN�   -�� p��m� u� 6�  �M�ݕ쨇�yUT�3UQ�-�j���P���N6턵#8�@�M�   ��7m��	  =l�l�@ � z�6S` l[�l@]2��X�V�l�
Ku� ��`�)l�m�xi��gZ[F�-   X�� �nm���� -�� 	   v��@8C����R�� ���z�֐H��p�餎�$  l�p5� HH.�pm���n�%�Iή�'H�Cm$��g��b�f���5��8m�h�Ӕ �Yխ�[֒z��	.�	j��ؕwgq��5/�n�]u{pd�;���P0�l��D�i�gZ��YP�ю�ۨ�����{kjr��ZI����r��O0Sn�W�o� �x�<�$�js�+dv��ܤ»S�s�㗷����soZ�b�oJjm�OmҲ�9�Rհ��Trl
폓�7|�mz4���Ɲ�c猆��%�)�#�7f#B���������ݷ B�Uʫvـ�/rBn` V�k�7]Kv�G���8;j�
�]U�*�m�[v	��LR�Zy�Z
�u�=�6 i6۶� 5�vg���z�USl��vu�lۡ$�Ҝ5��Wگ���y^�7]h��a㱵m��h�u3���r�nE*���p[v�[u��r�Y-Y��4L@4Ur� ���m�� �g:��Un�^�M�禞��p6�m�V�WvI����)M�b裰��eyNwO#';�v�B��u�Y��ܱh!=uk6UU/�9��%y{ 	��U(�zn���f��cs��K&۶:K�cv�h'zmЁ8���� ]-4��ѷH�gr-�C��k��@0c��Zt2�*��K�&L6{�5V�
�*�[���+U[�"�M�c���2���%�n���1b1�Nm�M�,Km\��#���4�V��^�GCb�U����fxw65 ɹ�l� ZpP�V��1c�lq�7�v�S�n��j�ME5��6��3k� -���>���QZ�l�l�UAz� �"��9�I��K��R�5*ʵmJ�P���IҔ�]Uu��㳠 ր-�� Izk��6�5���e[R m� rM�H[շ����K�ě6-��� �`,0�mmm��Ӊ��A�͛b@k�����.�L �ݛ:$khp8      R�    e�d�m�@m�H�6�����I����8 �ր�$�Jlε��2K�-��v�[�	�#ige�Z��]�6i9�\m�8�`ַm�u��I,��A m�#Z��6�$ h�:lڷ`֓��mq���%��;����i�e�z�kn�^��n�� 
�V���o[A�c��v�Հ v������ՀkXq�Npt�ml�0H ��kJ�[m�Cldp
�D�X���ɤW� [�kv�GG2�~>O���L�(�cz}m�I^y]�Z��RکM�%�N̮YѕJ%!Π`m�lm��v���L�
*�vZ����ٰ	 ���i-��U��	��%$�Z�n�� �ʛ`F�Ustԅ�hՓUT��UPgT�-*�@R�5�[u�m��m�     :B@ ��:A���(UUzӂ�  ռl�Q��  ��    ��lsm�p ��          @ m�H���m� 6�     V�� 5�� ��`   �> m���$  �` �$'-�           m�M�6�8t��`  $ m� l([Ki�
��	�U?� *��P��ڢ?� Dq�������*@1�)�h(���/��(z '�#���Q�'���!T=L\> �)���Y�&	�l@6?�!�)@�Pj��' ��8��!�@�B��B,!	$XI$"BHq"��U�ث�8��8�-D��Q>�x�|Q�EM*(��R����SB�DpT�
��������/ �J )8"��0C���h��!�O7V�(HB$
��8�xp����"��P�U�Tv��A�A�"�!HXH˒,B	�Tj��	U���R���Z�TS $�`�b3�  z��1Q('�0� `�� (������z�A4�(s�G���A< ��C_�
���U�4`C�QD
�4��P> @ ��&�H��z&��%QW�;T{�����{�����  m�  l��  @��   &װ  �  �   � ���m�     ��i��  �6ݺJ]i�q�Z���e��2n@7M[�4�G<W��v��-���R��v�a��y�k�8(�tm�����t��78w\�K��OZ��u%�t��Nr�V�E��&��.    m  �6��� -;�"Ѻh{g�\��V���m�u��*�-&k��b��R�ۂF�i�^-Z�[�1���QX�g�ng��h�m�4p�V ;
�G��lv�c����r�d�������iv�sW]/Jʡ�tQH����s�s�h�1�q��{k*��eU�!�� ��@̄���9�`�a2R���x��=��Sv�n����נ�DV��Q�ݟ vD*!��j우w VN��y^��Lv�l�m0��ԍV]'Y�7>L��@u��gAn��,��t�H�m�LaN.˳Y�m��$���KO��*�����=���f�-�����W.�P��v;�J��$��B����޲�R�K*�P�ˢW�`�Q��g���i�ۊjr��59ƞh"Jj����㶺�3��#�TcK��n;v�t���V:����j�&��s6��<�l�z�;d�z����t����j8��yVRe�3��=��t��
��1��t��e���s���zpF�������ɲ�켭��v�M	���(r��nק��<�;<k��ѸS:�y������]m��ۍ��ƛ[Tk���*���WL;0�^z�(V�l�UE\���@�$�e)��k�'E�I�Q�^9з8.C`5���Z�[s��M��Px������[��:i֩�d������h��t�d�'dmj޸i��� �i;h i��h]5��@ ��,�%�f� �w�;����P�
��
PG����{qF��$P*�`���'��k�f��b�5T�mL�B]Q��i��iz1�5YF��d&���}�6��m	s�GI��5��]��Ζ�t��Ĝ�u��.�f�k���C����M��,�ٺ�a��9���&ή�v���Gl��2{^2�j鸺�u����ۀ ��ȳ���ɺ��c��=m.��G��d܄�����j�b��Lոf��F��w�nMj�Y�S�۷	�aɁ�r����l<�v�W<��C�����
4R<�W���p���hwY�wZMl��"��'�_[4z�f�{�4]k�>��5Hَ8�I7$�=�u���9u�@/���R{q$�a 䑚��9u�@/���n�@�1��$(�FF���Z��٠z��h�S@��%@�m8���`��j]����q�jQu�B�;s{#t��{WG�mua�
F���٠z��h�S@�ֽ�����1�&���rX���R�,J"��,N�; ��hQb��I1�&%"4�4�1��������Vv���ǘ6�iAI�N0��@�ֽ ��h�u��;��&�Hԃ�dx��@/���]F�{�4]k�*�T��j�]��Oj�&a�L��f��=�-����nT�]�N��)���,�I�w[��_t���mz}�h�uI�1ēɄ�܁�_t���mz}�h��h�IWq�S#@MQ`y����6�"R�RP�kwn��}Қ��\�&6
F�6	7ٽV�u��������ٰ*�aQ �⑦5$�;���/���<�vl}�V(��nzjdc���g�I'[6 �[\�nָ����n����jk��,�8�tc�j��}�~�'�@� ��4�t4��gX���7$C�����Y�w[��}zS@�:���#RE��N= �fՁ��ag%
!�v�>��՗I1��crM���Җ�w;��B��N����t˵O�d����}zS@� �u���h/B*n4ډ6�RZ�ݳGS��pu�N���	��κE��n������FF���U��{��-�C@������6	�����r= �u���h^��*����s
����#LjI�[n����M�k��Y�E���	�!2E��}zS@���^��m��g��b��ܑ54
��@���F�oO�;��,ە���sd.����U��EYYV�Z�*�s�F�zm��*N$u�:YH��m�p�:j�l��[���pm��fn��kg�ȌK�vm���<L�ŷ(�U\��۟u۷n4��=6�$�؍�[q�)��^ i�ܹ�ro^�d{NU���y��Y]���U}�㝎����kuա�9��շ��]�8�7r՗�����X���W�o�*=�w~�{�-�ݶ����G욺{M�V��M�B-��Υ���V۳mn�R	T�.;�6ߧ��z��h^��*���V]$lƤd�H�#�-�Cٙ���g�@��~��^��x:�� �I�L�i�ץ4
��@��@�� ��*�/�Jdh��h[^���^�m�ץ4�@��X��#�z/uz��h^��*���������u=�ٱ�mӯf����`���Mcq�9qs�:���Nѫ<�M6��@���ҚV���?�AW_�@/�b���ěnd�N���fч��Ōh��h	b� E$�	
�``�F�)R�HP��H4cR�X4�D�e-�!B
�a��TB@���5�������3�PRc�&���U�����ۡ�}zS@���kd�DG#	Ǡr�W�[n����M�k�>�e�F�jFBI �z��X	/v���Os�1�6lf3�k�K#Ǯ}]�8f�Q�;�%�(Η�E�l{#�r�^���`]Y���ץ4��h����t4�$�����FF����}V���^��론}zS@�����&���Ȭ~͛=����?BIyBIU>����;�h���TH6
F�JG�w�\4�JhW�h����,\ˈM��L�E&ץ4��^���K�����`	�#m
H�l�8��\�8mn�sǇ7cXwj�:�`]v�^����܏��䉨�}_U�r�W�w���_�{���;��n]�T�N��E��9{��;�\4�JhWj�>�e�F�jFBI �zwK����M��Z/uz�z����$��U�i	C�m�`{�����6	��Q�s2���{:�)�#FC@��V���^����}zS@��P#GXԐǐy"F68v\�=���t�wNG���g��Xy\��k�]JFcN=������@��������*L�6��@��p�>�)�|��@��^�{���q	��ɒ(��@��M�mz.��� ��3�Prc�&����	$�=�6�ޛ3+Qa�"O����?~/�[$jb�<j4��wY�wt�hu��>Vנvfw\�$IamB�ݖ��-6 U���ȶ�;r<�cVÞ�:S5�Ε� p�T��q1;��S���N�;A���;nѺwNc��额��&ݭaN���x���.�7n�'-�er�]�n��){I�$�S� �3��n'�����v��q6�j�q�q9��ݸ��<\;9�l��BK���$�/W����ڼ�p��]q�"j��vV;����������L�)VM���\ml9���k �ŉ��t@��i7��n�m�o�m4� v�{��E��6��?=ݛ �fՁ�nksrQRۘ�TK��X�kK��P�M�}�6��VfV��3SogS�e8�у��>Vנ�O��[g�4oW�h���d�-�H��M�%�u���m���>�)�|��@��@�
�$L�ɠwt�h�)�|��@=�����}�!(�c�I�]�Tқ\:۲�x���au�y����5��=�N�©u�Ev����_�� ��_�$���5$�wm��H�?�uF��Z�̟ ���������׻��i�MI%��p���ekRIu��k�#SsI���$s�MI%��p���ekRI|��K�,�8�$RI�H�����}�Is���$�v���$s�MI%�^�?��O�d�M�>�$��G�$�v���$������}�������-s�9&�Ůk��e�B�S�v�q�m>x�d�ޜ�[�pq�L� �����_�$��lz�K�����%��=I%��\�#dM
HcN?�I%���$�wm��K��z�K�m}��3�1��;��55
H���߾�}'9m�߳���
 �K h0��ѽhvɄ�	K+(�+��nm��]��Bl�k(*&��n;��rd�l�3ۡ���L�ا#ϭfN�2��l�@E+iu�k��ޱ�e�.������Pw i�HIY���p�t@����WK ٺB���I,M�r�2SXJ���m�Fl��$̺8˲B�����X@�Xn���ù;��WnΕ�n�y���$��-5BQ*�X�k�
�4�(�K�	��5�1�$��_<��fy���u�û���]?/uFv�K]����	v*B�� Fi�t&�� J<�WBi�Si	�a�Dt�h=�H���h
>��A U�ꁰ ����x�<��}�5�[m�^���^�w�� H���I.VQ�I/����$�;cԒ]�ۇ�$��?�v6I�nH����ޯ�Is�=I%��}�Ir��RIu���M�����6{���X��;��e��:c�秭�`�#K�A*��n\AOߠ%���$�{����%��?ٙ����i/?�������w���(=SU�S� ����$�;+Z�K�z��I.n��$���I��F��$na��%��֤��ޯ�K���I%��}�Iq(�x��a��֤��ޯ�K���I[���s��7 �'�"�B�QZQ�KaO;�ss33�x9e���ܨ�R?�I.n��$���~ϾI.vV�$��s�I/��j��7n1�(^u<�NC��C=sv�����ݒs�4�ں���L"��$N7#z�K��p���ekRI|�W����i*����I%�G�����E�}�Is���$�w�����oRIw�n|�E��s��q�nH�kRI|�W��%��ޤ��v�>�$�YbԒ]j����LQ�x�jG��%��ޤ��v�>�$�YbԒ_;���I�e��I㉧R7�$�ݷ��ު���^[m�]���-�߽�3v�k׷}�{�����oߟ:�55R�R�5�m:�l �%������c��lÕ�m�*lPUUY�V�3�Nc��^�˭g<f����Kڢx�eR9�N8��s��ִW���]Cח=v#�x��J�t�����NK��KX�P�E��)����7A;�q�s����n�q��d��u�vպ�ۧ�a��]؝�z�n�v��*�Yź9��i�!$i���;�7[9��jѓSF��WD�/P�wk���63;�g��<_Ϟ>t�2���OVjw�3� >��-��� �o�� }?��ߠ�d�$�ݷ�I%{�ǋ�6���A�I/���������/��J���}�IUҏRI}��$��m�$1��$��W5$���}�IUҏRI|�W��%_bp�#�H�M�5$�{����%WJ=I%�_�$��W5$��s,�<�$���I*�Q�I.J#����6��zj�m���6�%���j�q��z��@f8�E��BwgO���@ֱ�\�U�Bt�Sɱ�)���^����$+��I%��}�IUҏRI^��k�#SsM���%/���ߧb�
\�ݹ�w�s���k����sg��Q2�u5�MJ�s#��8椒�w�|�Ut�Ԓ_;���I
�sRI}�ԟ̄bO�c���?~m�ON�m��=�?�6��6j�Iw�n|�J�%��l##X9�$��g�$��W5$���I*�Q� }���`Y��۳8�	48�=g����)�7�s;sv�n�O��:ڴ�m�$rO�I!^�jI+�n|�Ut�ԒJ���J��
�G��4�jj�m�m�?~�B��|���m��{��$��W5$��YY`x�@�a9�m���Mn�m�߾�r��� ��(�X�E(���˿��n�o��p��^3�YqcRD8��%��GZ�~�s���{�u�����o�s�ފ:?���| ???PO�E�ܸ��ߠ!wW5$���I#��5$��l����o�ݰլ0�̼O!3�k`�1��s��v]�Q詻\��Qՙ�\0ӁsRI^�p��<�SRI+�ϾI!wW5$��֤�d#����H�MI$�[>�$��\ԒVݹ����{��C��g�/6I31|%�����H]��I%l��$��j��K�p\�q�Ғ�'�$�����J�n/�I#��5%s��cn�>�$�� WR<`䉤�sRI[-���$yڦ��V�>�$��\ԒV�I��X�����/[uu��H8��Kګuy�<�(��s�9g��N���z�����D��j��I[l��usRI[-���$��Yլ����"q8���V�>�$��\ԒV�q}�Iv��$���k�Q�̌BNO�I!wW5$��nNr�@kS�w�7m����s��|�)�MG�ln&�㚒J�n/�I#��5���ݯߛ|�/�
�����5o�77%#s��\�v�nՁ�%����v��s��?���;B�ڏm�$����YYV�U����Y�jћ�� �[t���vha.��US��٧x:�q�C�;���RsWY�����2J���p�����fStgv銵*�^ڲ�[q5��͎+���Fε�U8�BN�&�����Mv������q<{q�<5�^3�=�&�S����|��@P.qƌ���\.n�:�zQ62q͛n��U��{���w����% TJۭq�of��{km�a�Ҏڕ��s�1c�g�=�{������9�=ZL�}�~������ffՁ�;��B_���=�e6�q�ҒI�wu��31"���- �wU�绳|���34L:Bܴª��s5V��'`�v����3�ﾛ ���3�MT�%J�
���NÒ�߻��}�6��V	��rv�i,���jLjH�NM�����C�ޯ�n�rv�ݫ�+u�9��[�;�✘�qgi�͸s����0l��Wlg��u��1���wg���8��"�݃�z���N�7۵��}�6f�]Dԡʙ�t悦��ǻ�o�
P���"!tD|�T���U��ﾛ �ͫ�I��w77%S�9�N�sJl���{�6}���>����~�;wq��chp�4H������߿= �o�`f��v�o���n�YM�SS3-�QUUS`��`t(ޮ�� vwU�������Tn&2G�0pQ(ݴ��㛞��� 6�]�Ǜ�mes����=��y����� �D�nO����ش�٠�k�����ᮓ�"IR�����N�7۵(Q舙���>�����N�Cgd�����*uT����ouX�mYiB�
i%�C}�ܞ��߿=�V�["�1I��$����o�z���N���ٰ�I���?u�?Aǂxۊ'94��Z�B��B���������`��`7�l�r�eq�VƎ!�»O�v��qBH-�����ܸ��^��{��L�P�}qNb�˿~zz٠����obQ��chp�5q��f���䡰�ޫ�{��5�vo�DBl��v�,Q��JH6����@��ŧ�	$�<� ����0�r�
��-��Xr��}�ܝ�vwU�nnՇ�lG!B2(�2
��#���B-! B���A!B@��G{�{�ܒt��g*D�!TTURv�ݫ�B��ߧ���4��Z�rT�㑶��u[��ѓG1Gk`�y�	ݫ��X3���W�D(SV�T�C�R��SU����s6���O�G�
!z@�~�������S�R:�LcsU`��|�|BJ&O�~�; �~��sv��(�J!L�oR��x&��i��M����ش�٠��{��=����&�̘�N]Rv�%�wU�n�U�nfՇDBI<��N����OT��S�
���j�3v����
O��W�ߧ��7$�r�7��ӭ$D�# 1� o���,Db�IԹ%qHV�H���zv.&�ӝaw�ͬ�M�Il]�ňT�%�5��(@�甌5��]d���	uǖh1%2sw6ć� �	�%�JkD��T��A��'.Mc��c5&����\2�C�hv\���%��!H�@�b0`,�]#�Zc�A�  r��$��-���f�]nk<�tD�*�D���`�
�X�H"��h�b�B`I��F0�K���"A.�Ig����y�	.�$޷�2P43X�)����I�ֵ�<��%��Øo�
sͲ�Kvhm�Z�bO���3#�=�#�bM�A~K�-n��oz:
T�������H�4�&#7jho-Ҕ"5�Y\�9W��5���kW�[5����9���iɹ��۪�n��9�$��fn�9�2�X @���2 D�A�A�E � D��5��%*A,R5%0�ҙ9��� m�  [Sk�  �   6��� �  �   � ���       �p��  UPq�N�T��FGH�`���vն���eD
�>3�e�����@|��8ue/e��{v�[,�f��J�*4��+�ڪ�oTs6R�m�)b�i�y孱��u��r+�]�h����     [@ 6�u�HH� 8K�A�@ӣk%�gb�-�mJ���\����N+Wkhvm�R{d�����-kt$u��;���0l��0����\��s�۫�4]t5�F�E+�F�ONۊ�8�nqk�jM��!_+�G�rj,I����Xq8_7h�2v���r!��]����M�1���]8X�%P�/n����˷;��F�<��s�c5ˇ�!g��p7l v�.Fa�]D��V�QuF��˵�T�퇝:��;���;,�s��qҮ�ۨ��:��̾]e�����y�.�{<g�5�\ۛe{xq���rm�ٶ[U��kvQ�7j@�ۍ�[gj�L8�9/Lخ2�:6�����n2�X������@^�֕]�	N����n*Yq�ۑ�j�e�t�=��4�ׯMHKd�m��)�4���5��=�˽�^^t�H�N\�/m�#e=gm�1�Y��ܾv1۳��F.Ӷ۰.��gqX��{(x�'���і���uo��1x/l����g.cvV�u�Qד����gA��Av��"�u�������LUÞ��3]6̦��;�:�6�]��&1��{gK�й㵥��6��7��_@an�$D�U����Qn�ݢ#YS�ോ]"�lv��(��<b�y��;�1��ţ��s��Nմmvrs҈N�"�%[C����zd��Y0l�Ҩ��mYK�6�ќ[sj��o(�[l�` 9��L-�l g	�6�m�]5�L� -�Ni=1�� ~w{��׻���w{���D@�C�H�����D�A=LT!�G��i*������d�y��֍e�333.(-�iͳl Wm�E�ÊIT�GCl$;-�f��z@5�lH�v�a�hL�
����<��k��qms�1�ޱ��@:x����Xx7/��7Jr�ٗ��@7��j ۸�z.��Ϋ��q�riM�i(�$K[���\G��l��]�'�|���4����&�筵�um���IN!غٗ�R�p���Jt�+Jܯ
߽۽���ᱦ#���Y�Aʚ�n˚'�T*�:��(����l�l��"e����ww�����Gm) ےp����=]���mrQ����V�	�H[��UU9nf�����w�B�ûz�w��w���VI�	�$�$Š����VrQ	��z���N��Kmb�.��R���â&�{��;���ܝ��9BI7��Vn��.�T��!�75V��V(�Q�]�� �� �l�/[�m4���AL���S����&�c�rZ�C[�4��Q�vH�/~�����Flx&�"m��O��_�ش�ٳ��b^���ӑ,KĽ���ӑ,K���{u�L˫5�as-��.ӑ,KĽ��ͧ!�N��$ac!BYHRg���l%�@E����5���P!�0wk��w�P��6I7����(M�ӑ�3A։�3f�ct2���3p}؉�H��b_|�siȖ%�b_{��ӑ,K��o�v���
ACQ5��������Mh��3Z���fӑ,KĿ���m9ı,K߾�m9�Bı<���]�"X�%�{�{�ND�,KϾ���isY��K��Z�fm9ı@�/~����Kı<���]�"X�%�{�{�ND�,,K߻��r%�bX���Y;�9ul&feպ�fӑ,K��o�v��bX�%��m9ı,K߻��r%�bX��}��r%�bX���g	%�(抝λ��=`X{l�7G;��Jk�l�s�h��N�Y>�����7}����拙�iȖ%�b^���ӑ,KĽ��ͧ"X�%�{��͇�H �Q,K����ND�,K��m:~&��d�3.�k3iȖ%�b^���ӑ�,K�ﻛND�,K�����r%�bX������Kı;��պ�̳2�f�[��ND�,K�ﻛND�,K�����r%�C�\@�m�`)�����1  b��
� "F��FB*���F 0�L�{�?fӑ,KĿ���6��bX�'���s4MkW3&��3Y�ND�,�Q �����?e�r%�bX��߿fӑ,KĽ��ͧ"X�B"�'�}�M�$Sӽ���3.�Ѭ��Yu�˱$D���+ ���sv��	��w{��Ȗ%�by߷ܻND�,K��Ԙ߬JZ��ڻ\�e$��wKm�vݲ�D����8Wf�VD-ָ�e3v���m9ı,K߻��r%�bX�}�y��Kı<���]���bX�%��m9ı,O>�N�e��f��.fMkY���Kı>���i�(%�by߷ܻND�,K���6��bX�%���m9Rı,O}�N�Iya33.��fӑ,K��o�v��bX�%��m9���MD����m9ı,N�����Kı/����Y��Z&d���3.ӑ,K?$CQ5��߳iȖ%�b_���6��bX�'�}�m9İ4�4��@҂�'��}˴�Kı;�KO��r]d�3.��3iȖ%�b^���ӑ,K���D�F� �����M��,K�������9ı,K�{��r%�b����~�BD�U����F�i[=��`�]nm���0�K��s��������Mf�[��ND�,K���"X�%��~�r�9ı,K�{�ڧ�B*@
'�5ı/����ND�,K�v�9�&����Z���iȖ%�by߷ܻND!D�MD�/��~ͧ"X�%�w���r%�bX�}�xm9�,K��k���Vh�Ys,��e�r%�bX������Kı/~�siȖ%�b}����r%�bX�w��.ӑ,K��~-�s5�5�5�̺��fm9ıP���6��bX�'�}�ͧ"X�%��~�r�9ılK�{��r%�bX�}'w;irk-֥�ɭk36��bX�'�}�ND�,K �o�v��bX�%��m9ı,K߻��r%�bX�(�������s2�f[s��̓ys.7e�i�M�$���3���P�q�/e�R��&�URl[1�76Nڞ�T�[���ll0{v�tnul�k�*�h�v�'��:v�x�e��V6d�zn3�[N�����5�`�{v�i��iv�����ݍ>v3��H�w�If������:�"����rX �/b���^��I�f�7mW7�r�dj�69Ȱݩ�;J2�w,��n�L�u��6�hg��ݓWc�=s�N{��ں8�n6.І홙u5sS�%�bw����iȖ%�b_;��ӑ,KĽ��͢�Ȗ%�b}����Kı/���d5�ZkD�332�9ı,K�{��r�bX�%���m9ı,O���6��bX�'��}˴�Kı;�KO��r]d�3.��3iȖ%�b^���ӑ,K����iȖ?�T��Dȟ~��]�"X�%�~���ͧ"X�%�߾�̳Yu�%,�Y�ND�,A�@u��?M�"X�%�����]�"X�%�|��ͧ"X��~Ab.�k�~ͧ"X�%���љM����J���a
HRB����.ӑ,Kľ}��ӑ,KĽ��ͧ"X�%���o�iȖ%�b^�����g�����C�����R��=6q����:SZ�f�f�ɭfj<E �T`��p�53.�Ѭ��Yu�˴�%�bX����ٴ�Kı/~�siȖ%�b{���؂?�c�MD�,Ow��9ı,Oߺ[�ٚԚՙ�f]M\��r%�bX��w���=h���"X�&��}�ND�,K�����r%�bX�ϻ��r'�@�MD�;�?n~��k5u�s2kZ�ͧ"X�%��{��iȖ%�by߷ܻND��� D�K�~ͧ"X�%�w���r%�bX�{�%�ɩY��u5u�iȖ%�by߷ܻND�,K��{�ND�,K���6��bX��'�}�ͧ"X�%�|��vB�MRa���v��bX�%���6��bX����m9ı,O~�}�ND�,K�����r%�w������������^�!��+Kv�N���Nt8{hggW[m5eؽ/T� s�3˖�̺�k3iȖ%�b^���ӑ,K���ٴ�Kı<���]�"X�%�|��ͧ"X�%�߾��5̓S5����fm9ı,O~�}�NC��MD�=���˴�Kı/���6��bX�%���m9ı)��|fSCnj�mҦ�XB���'��}˴�Kı/�w���K��@
�j%�{�{�ND�,K�~�fӑ,K�����e՚5�\�.��v��bY��.�k����ND�,K���ٴ�Kı=���m9İ?MD��y�.ӑ,K��������I�Y�&f�j�fӑ,KĽ��ͧ"X�%�/�}�ͧ"X�%��~�r�9ı,K���m9ı,O5ޗ���Y��6��!BHÉ����Ϡ���pW���k\s������������j��"SMkY���Kı=���m9ı,O;���iȖ%�b_>�siȖ%�b^���ӑ,K��߈Y;�ɩ\��rj�&ӑ,K��o�v���A�&�j%�}��ٴ�Kı/����ND�,K߾�fӑ?(� �MD�/����!rL$ԘfI���iȖ%�b_{��m9ı,K߻��r%�bX����6��bX�'��}˴�Kı;�KO���5���e�kY�ND�,TlK߻��r%�bX����6��bX�'��}˴�K����2D�cH�##	~�!�D�X�����ND�,K�{��S���L�R��u���Kı=���m9ı,O;���iȖ%�b_>�siȖ%�b^���ӑ,K����a%�fL�����\�PʡV��À�����k��ˇSZ�������ww?~�9>�eJ��Ko��"X�%�����]�"X�%�|��ͧ"X�%�{�{�� "j%�b}����r%�bX���\�̺�F�˙eֳ.ӑ,Kľ}��Ӑ�#���b_���6��bX�'���M�"X�%��~�r�9�����z��{��������즨 ����,K�~��ͧ"X�%���o�iȖ?�5Q=���˴�Kı/���6��bX�'�I���R��j˙�Z�fm9ĳ�F*�R�}����r%�bX����e�r%�bX�ϻ��r%�`~b @����߳iȖ%�bw~��Ԯ\̹5u�iȖ%�by߷ܻND�,K��{�ND�,K���6��bX�'�}�ͧ"X�%����#
A��RQa��Ԟ�je35nk33-���`�K�R�T�K1�[����*�8�`�Ϡ�nQ�l�F���8m��ш����(��!��w.���s6/p��Upod�1���9����5rgqvTg�km��\ �ڎ��j�E�{ev���\ms�;��{|��<?;���Fy[r%�����ؓ���6�f�^�<h�Ἆ�(���Z�j�b���J�e�6��f�v����îK�9�O�j��7Qx[�I�3Y2\�冊kY��z*�o\��&jL3$�����Kı/���ٴ�Kı/~�siȖ%�b{����Kı<���]�"X�%��rZ|t�ѭe�3.�Z��r%�bX��w���?�B/���,N����iȖ%�b}���v��bX�%���6����5Q,O���uNf[u3YKK-�fӑ,K�����iȖ%�by߷ܻND�,K��{�ND�,K���6��bX�'���j�4MkW3&��3Y�ӑ,K?0�Ow���9ı,K�~ͧ"X�%�{�{�ND�,�A�O���ND�,K��k���Vh�Ys,��e�r%�bX�ϻ��r%�bX��w���Kı=����r%�bX�w��.ӑ,KĽ�N�oщH�ָ��/\�������M��+˺9���jY�O|��ޗ���]���L��r%�bX��w���Kı=����r%�bX�w��.ӑ,Kľ}��ӑ,K���;��J\��Ys2kZ�ͧ"X�%���w�Ӑ���R��B6��AUD5a�0��B�	)���
��>P�j&�X��7�]�"X�%�}��ͧ"X�%�~��ͧ" X�%����^�ծ\̹5s�"X�%���r�9ı,K���m9���Q5���fӑ,K�����iȖ%�b{�zwY%�1��fd��̻ND�,ElK���m9ı,K���m9ı,O~��6��bX� ���߹�.ӑ,K���KN�����32�5�ͧ"X�%�~��ͧ"X�%���}�ND�,K�{���r%�bX������Kı;�턒�5�h�tN�8�&*Ɨ�]���`LB��%mƻ�����R	� �05���{��%���w�ӑ,K����v��bX�%��mP9ı,K���m9����ow������=�*��5�=�bX�%���r�9ı,K�{��r%�bX����r%�bX�}�xm9ı,OO��jk.���j��5�f]�"X�%�|�{�ND�,K��{�ND��u�(�l]�42�(T����Jh�dMZD
"f����H�@�`�e��*c4�4%�cU�i�D��+�@�,hM+|�m/h�a*���a�"#t�oN�6DSDa�i6�4��4@�.�*�x@�Ib��db�.��WQ5�L�h�]j�\Ա@�F�$��� �ЕXYZ���#~P�/�!) �$l�P ܀Ȃ�(�l6��>pt�ʝ� '�/E`!�G B���v���R��؝��p�r%�bX�{���iȖ%�bw�﹚�5�˙�-5���r%�g� j&��߳iȖ%�bw���iȖ%�by�wܻND�,,K�{��r%�bX��N�vҗ.kV\ֳ̚3iȖ%�b}����Kı<���]�"X�%�|�{�ND�,K��{�ND�,K��oӌ�%�4�q�b	m��p%�%��x3�:�n�`�:�E8�S�:��{��g�=�E�rj�ND�,K�{���r%�bX������Kı/�w���*�&�X�'{��6��bX�'����Y%�1��fd��̻ND�,K���6��bX�%���6��bX�'�}�ND�,K�{���r
6%�bwܖ�34kRa��Yu���Kı/�w���Kı>����r%�bX�{��.ӑ,Kľw�ͧ"X�%���3,�Y�����fӑ,KK���"X�%���r�9ı,K�{��r%�`x:wT�	[B�f�l��
:��Zh� ԉ@�.���nD������q��������r}�ʕez��r%�bX�{��.ӑ,K����6��bX�%���6��bX�'�}�ND�,K���m�d֯�kZ�h֜z�ձ��-�.6-�;v�Gڹ����K��p�b:W������W��Z>{���ou�b_~��ND�,K��{�ND�,K���"X�%���r�9Ǎ�7������/e��c�����d�,K���m9lK����iȖ%�by�wܻND�,K���6���oq�߿�~�ߡ��Wej����ı,O���6��bX�'��}˴�K�T�MD����6��bX�%�~ͧ"X�%���Y/Nj�3Y��\��iȖ%�by�wܻND�,K���6��bX�%���6��bX"X��ߕ��Bd&Bd,���@�*	tʢk32�9ı,K�{��r%�bX����r%�bX�}�xm9ı,O=���iȖ%�bN�� ��@�B"Dѩ�}�����Z�heZ������p
�U]V�����U�άJu�&m�nx���5U�=+��N���Z���c�ۇ�jZ���KY�5t��g�Pb�p5���pٷVu��b�G�0vzn��f�Z9�n�/*u���z؉�n��ƘN�۷
�Ҹb��	-��z��h1�ќ���<u��F� ����..;Fq�n�/Sgu
�.W�f���݃�;l3J�U����k�m��[;�y�؝ڹ=ph�9.�ڽ�r���r*V������U����K���ٴ�Kı>����r%�bX�{��.��U�D�Kľ���6��bX�'�~�n��d��k)ie����Kı>����r
��bX�{��.ӑ,Kľw�ͧ"X�%�~��ͧ"~"�j&�X�>��j�55�\̚֌3Y�ӑ,K������iȖ%�b_;��ӑ,KĿ}��ӑ,K����iȖ%�bz}�MsZ�5�,��5�f]�"X����M{����r%�bX����6��bX�'�}�ND�,K�{���r%�bX�v|S��/#Cj9��������oq�����ND�,Kȱ{����yı,O~���v��bX�%��m9Ļ�ow�������	�^��փ���,Z-��<�us��#�-��gl<��f|m�A��\��jkZ�ͧ"X�%���w�ӑ,K����v��bX�%��l?@�&�X�%�~ͧ"X�%��Ӥ�_�5i�5��ɗXm9ı,O=���i�P8�Z���$`B!�1D@��bX������Kı/{�siȖ%�b}����O�AU5Q,O��B�I��fI�ֳiȖ%�b_~��ND�,K��{�ND������p�r%�bX�������Kı;�1�陭j˙&kY���r%�d�\�����&��	����A$Ny����D��|�{�ND�,K�{�uMs$�W2�[��ND�,K���"X�%��	~��^m<�bX�%���ٴ�Kı/�w���Kı>�����<�[^�6������i1�<����wA�OZx'��w�'�Ǆ벜��J��t�O"X�%��߿k�ND�,K���6��bX�%���6�Ț�bX��p�r%�bX���\֮MkE�32�k5�ND�,K���6��bX�%���6��bX�'�}�ND�,K�{�si�!bX�'ݟ﹚֥�kZ˙Mffm9ı,K���m9ı,O���6��c�U<DQ=���e�r%�bX��~ͧ"X�%�ߤ��[2[�\�MkY���K��.�w����Kı=���e�r%�bX������Kı/�w���Kı<�|K%��Zd�f��e�ND�,K�{���r%�bX%��m9ı,K���m9ı,O���6��bY�7�����w��%9hb�Ĩix��$�<;m���Ƽ�O:SvѮ���q��[n��l̳2Mff]�"X�%�|�{�ND�,K��{�ND�,K���Ȗ%�by�wܻND�,K�����֬��f���ͧ"X�%�~��ͧ"X�%���w�ӑ,K����v��bX�%���6��%�b{����KMf��֍Ks3iȖ%�b{����Kı<���]�"X�%�|��ͧ"X�%�|���ӑ,K�����W���L�ə��a��K�lN���.ӑ,Kľ}��ӑ,Kľ}�siȖ%���H*A��
f�_��fӑ,K����5�j�ִ\�3,ֵ�v��bX�%���6��bX��ﻛND�,K���ͧ"X�%��{���r%�bX��~��wYsS&���_S���s.]�$spM�ݒ0t�����\�t�I��ԮX������ou�b_>����Kı/�}��r%�bX����]�Ȗ%�b_>�siȖ%�bw�:o���-�.f������Kı/�}��r%�bX����]�"X�%�|��ͧ"X�%�|���ӑ?�����b{��Y/㚴ɚ�]f�ffӑ,K�����˴�Kı/�w���Kı/�}��r%�bX�߻��r%�bX��;��f���2��5��v��bX��D����6��bX�%����ND�,K��{�ND�,K��}˴�Kı;�1��u�.d��e�ͧ"X�%�|���ӑ,K��_w���yı,O�~��ND�,K��{�ND�,K�����[x��!Jd[VӖ� �6F�Ɲ���&kͪK�d�76u��ᬩSQ�әI�x\�βMp/:�杣�yzS�[��	]���\�K�#�����۶�crs��9l��nzM�ܠ갼�I�7�n؎A���u�ꓯdv�7K�vݸ�fx����lu�/X<�b�˫�̂Wk2�l�Y���:9�kۭ�*񤱢"�&M�yXBD����tv��Ц����;r[��6��n@t�%�OYٺ2Giz��k%nW��=���7�Ľ��ٴ�Kı;�wܻND�,K��{��0$H'�5ı/����r%�bX�w�5y���\̚�&ffӑ,K���r�9ı,K���m9ı,K��w6��bX�%���6���!H�GU5������ʚڣ+G�w��7���{�����m9ı,K��w6��bX�%���6��bX�'}���iȖ%�b}�������+r����{��7�����$X,"�"g߿fӑ,KĽ����ND�,K��}˴�K��f�k����ND�,K�d�o���[�&�555�ͧ"X�%�}��ͧ"X�%�� 1H�B ��~��O"X�%�~��ٴ�Kı/�}��r%�bX�w��u%��j�5�ˁ�N!LZ�g�W8���mT�	���s�=��OK�tq��cb�t�N��������ow����]�"X�%�}��ͧ"X�%���w����H�R
	<���%�~��ٴ�Kı/���~��$�2��5��v��bX�%���6���v(I ��D!��pP����'��6��bX�%���6��bX�'}���iȖ%�bw�c��2��I��\��r%�bX�}�xm9ı,K���m9��A����H*D!�2'����iȖ%�b^�fӑ,K���횚�KM\ɩ�Y�k0�r%�bX����r%�bX����]�"X�%�}�{�ND�,�b$$Qb,�O{��{���oq�߽����g,43��_�,K���r�9ı,K�{��r%�bX�}�xm9ı,K���m9ı,Ou�{[.�ML�ɣS.�ӗ�o6�kG\T�Nxq�#^�*c.}��Bӽ�}����om���q�o��Y�MmQ�����X�%�~���m9ı,O>��6��bX�%���6��bX�'}���i��7���{�?���ڑY�����,K����i���&�j%�{�߳iȖ%�b~���e�r%�bX������Kı;��7�IL����-�6��bX�%���6��bX�'}���iȖ?	� A+	
�,�e hF-H��(Ab��� �&���E[�/y�6��bX�'��~��Kı<�|K%��[��f�f�ffӑ,K���r�9ı,O5�{��"X�%���w�ӑ,Kľ��siȖ%�b^��!�&MW,̓Y��iȖ%�by�{�m9ı,Ȑ������%�bX���6��bX�B���w�	��	��zɞ���T��{D�[�,5E��;f]̧W�ۡ�������ؽ+���y�f�����}��{��"y����Kı/����r%�bX����]��H��MD�,Ou����r%�bX�~�~�S��M\ɩ�Y�k0�r%�bX��~�m9ı,N���.ӑ,K��^���r%�bX�}�xm9� ���j%��������ֲ�2�4d���ND�,K�߷�.ӑ,K��^���r%�bX�}�xm9ı,K�w6��bX�'���kY�Z��L̳Z�e�r%�g���*H����[ND�,K�߿�m9ı,K�w6��bX�"�B���U�����iȖ%�b~O��"0�F�?=�w���{��Ͼ��"X�%�������w���i�Kı?����ND�,K�{������oq�������"��a�ͻR�f�I��q�k��ٜ��ҹӎ�ڒ�fܮk�5���.Y5���0�r%�bX��~�m9ı,N���.ӑ,K��^���r%�bX�}�xm9ı,N�>%����f�W3S33iȖ%�bw��v�����:���'����m9ı,O{��6��bX�%�߻�ND�,K��u�2h�5\�2Mff]�"X�%���u��Kı<����r%�~F*�!���~���iȖ%�b~���e�r%�bX�����2�̓4Mf]�"X�%���w�ӑ,Kľw��ӑ,K���r�9ıP�5����m9ı���?����H�V�����o%�߻�ND�,K�F?����v�D�,K�}�����bX�'�}�ND�,K��t|��hE$Q"A*�z�c5P�4 �J��52�FP	@��
P"�i�!45)VcE��F$@��!@4���^�;��� ��  -���  �6�   J  �a   l   � ��        m���  oT��6���.Q���bI\aJ�h`�L�Z���i�gK�K�7;+���3��m/n�PB�WI2�N��OU�����ti%�:��e�AAd�㕭�X��rOF�em�h�OSl    � N���6�8�,o'$��l�u���M�9mֻ�N)�v����A..-���J�W4�=YÓp6�3lL�e�ݹ���B�T���<��V���d�/Jn���[�v��W8'���޹ֻ|+�}�6�P��C&fw[l�jv�J7�2+�έe�^x��^Q�3��d�	�
�x8�3�Y6�qY�K���&Bܽ�����9����b�[���ܶM�8��'n��y��;i{��KP3�mY�^j-F�c��bZ;\�������㧦�؈���툹��մ���<x5��7fgG4���:��Y5یg�9���$3��y6u��cT:)�o!ƭƱ=aĽ`�ܭ)tUe7mPI�kt+<\�
�AJ��P�1��Hj\�OA�lNd�$���n�t��j��4�՞��q�ܨ;<�m�`������w.����cm�}�c��L���v3�bۣo8v��RM�0Xy��r����q�� �ɍ�8Q��"�s��.]��)��\��ug[I�F�Uc�m�ۮ����r]vMԐ-a�����mǮ�u��w6�l�nی�d�0��& z�����m*�m۴�KQkT�>cT�f�E�S�՗V� [B,S]�Kh4:�y�+��ЛcSWQ��"���� "��y �n
t�n�]v\ە6�bRݪ��z�����E88�6맠�l���p���	�N�䝙 ې�eB��m� &ۤmnmUUS�.�UWTYWv�H ���$���`�	 )�"tE=�Pt |
 |����0E�]��>DN ��~�33,��fcm�M�j�N�� 8Ii����U�āYۣ����0�����moY9rG=��%��n#-�#ٕ�-۵k��v�G�mt�7V{s�,��u���zgZw8�ۦ�H��.�x�ԝs��ѡ ۳4��`J��I�7\���;��ݙ��s�b�Zzf���Rם<�ؤ4{p���Wn��Y���n�B�,9v���wp����D��;W;fҘ�6��^q�Uv��j0��p��k�{unR�I�s4�R*�z��	��3���9ı,O5�{��"X�%���w��� FyQ,K�}���r%�b]������s�g���Q������o'��{v��bX�'�}�ND�,K�{��iȖ%�bw��v���*�������[�ow�����Z�Y�˴�Kı>����ӑ,K��^���r%�bX����]�"X�%���ݧ"X�%�ߤ��JL�d�fB��iȖ%��
@?�D������"X�%�����e�r%�bX�����r%�bX�}�xm9ı,O���zsV�3Y��k35��Kı;�wܻND�,K�s��ND�,KϾ��"X�%���u��Kı>���ˌf{s�֓K��7�]���y�Z�c�u��rg>��:4nx�������+�?v�Ś噒k32�<�bX�'�g��iȖ%�by����Kı=׽�bX�'}���iȖ%�bw�,>:�MY�f��e�r%�bX�}�xm9Ez�%[B�i	$!ŕT% ��B#2FU%$��!%t��P
��MD�3]��m9ı,O����v��bX�'��{v��bX�'���59��ְ�]j�kY�ӑ,K��^���r%�bX����SiȖ����}��]�"X�%��߿p�r%�bX��}�s5��ֵ�Y�35��Kı=���ӑ,K����nӑ,K�����ӑ,K��^���r%�bX�����f�kY��W2���M�"X�%���ݧ"X�%��>�����Ȗ%�b}��~�ӑ,K���w��ND��ߤ�v��!������.b뺷�qd��^m#�;r��m�����j�a��(���zՁ��ٰ=��'B_(�������_(�UBn�X��f������Y�w;�hz����+�҆G�'UN���[,��*"l(A	� ( �A##V�J��R��,! �$a$�E����G����;���<�zl<%:%é*DMT�D(I�V�=�֬�۳a�O;{��jh˟�<�QŠ}�w4��z�6�=��v�
oR�b�MSd]tN�8�]���Wl���5��eG5۝[q��;]m�����-�)�������ٰ=��%��Nk�?0�oZ�<�E�]KN6�rd�H��u������s@�z׿���gg����7#22E�����h^���ֽ�]f�ު��$���ȢN-��ُ�߿��������%�%�Q�U���U�F,�@�
L�>^��z�4y�v�͵`D(�[�sL�Φi�5S)�g�t��+�d���q�=�;]�Z;��ȧ!9�{��TBWe!���Kt*��T��� ����e���U�}m��>^���˂�'RT��S,ޜ�|�@��&L��h����;��h�ѝ�$Ĥ�-�n���W�w[��>���Z�.hd�*&fIsT�>K�Q(Q
r����ﭖ�Nk�?n���2��m��NL�G��n�@�Ϫ�3��X;�v�b����BJ8J�I%a�zԟfje35�k33K<��� �UO+��Yaץ��q�d�:�D�'M���*��88 H��{u3�n7M���k�wM�
	5�m�f����׶^x(��hm�v���3�H�f�v���b��+�d�Ӝ5<mOD\���ս��V6덜딝��9�iOn��hm���wnKQ�⋶��7"C^ݦ�$�f�δK����n�t�[s2flL 3�~A�@ ��������W*�+�\��6�%�"O[��4q�]���lt���r�t�/2�-:�T�f��z~���vՁ��6�!/�-��Q�[�~Ů9�NFƓ�@��j��#��!(�1�}6w�[,ޜ�`z��R�� rC&h/uzwu�gDL�wu�t@yṮK�.\�D<��̰=���ۻj��K�_�@;*��x�3dfE"4�9������~�7���ݶX�Ukp5J�Q��;�1��c>i�Ś��:S�s�&�;��m��ͣ����V�6�??74�����F���U�^�P�p�Z�&��M]f�r����W���1DB{��3Ϻl��V/x�˶�Q���0�=��F���U��b^��������>η�7#22E�k�M���j�3}�`{��%��t�Z�jD�'���s@>�Y�{��%����`�	%���\�4�r^D�m#�I���jm�����"�Q��!��͇�P��@<� ���$0Rg���h��4����n��v�iAT��ԕUVf��$�=���wv�}�@=��(�@f(�̊Dh��l��V8P���!E�D�$D@`J�նJ��	*Z�I	
�k* �(���ϻ�nI����ܓ�)bŪi9N��SN����!?ww�`��`fn�,:�O�]����̒�LҢfd�5J�=�ڰ>��������������WZ�iL!@�ӣklK`l���Ŝ6�_]x7%I[�cM������i��Q�I1�r|��j4��Z��� �����q�q�r3#$Q�S,ޝ��!$��DL���Z�����uuW��FH��B$��>��V�f՜���X��v�X�Q�ŎH`�� �����F����krb�"�����s�pܓ理@�kJnF�@�Q�~���}���~��s@=�f��vS@BQ����^uؕ/�/$�0�ݸ�����k�����k���:�P���(�̊Dh^��[w,�ݯ�"�����K���)���&����������߾��ﭖ��{�ď��~C5�̃m�93@3;���ݶX~ݛ��ڰ<�%��̺�*���MU��w��,y�6��� ����������fFH�r�`y�vl�#�K>��/ n��X��g�G�o��'��n�h9�(6mҠ5UU \���/�@��N-U#b��8e��Na[�[�A^N�k��M�]1�lnq��=�u���E��ծG�j�ؠ'p����s�.��ܴ(�ݴ��sј6���za���m��n��mu���]p@��+=���7p�s���4�@�Y�;(�K�����ًuπ�����tAJ����V�w{�����|�����s�8��)p��.�Y��z֭�.C��L!���ND��.&n�C2@$��u�s@=�f��n�@���`{5�V��b�����X��W�D/�S'w�[,{��`~��V��0w5��7#rI�w[��<�k�>��h�l��.iR(�1G�8�J?�߾�>��V�nՁ��l�/��;+����@�۹���@�Q�yzנ^�ZQ���Iz֎�Þ�\�Vey���l��	��==&�p��/��w���}���[
�j\�w����`fn�,?ń�wmX[��]�.jYUT�S��=���DF"�S
!D/۳`~��V�n���%�Q	L�����J��QTU:��e����[n�{��޺����rC53.�32I��nO�G���C?����Xw��X����۳`{5�V�,�9 (�h�l�-��<�k�-�s@��T	aN7"��q
'2k	�񍸝��u[/<�bn�/��ں������(J�����-Ъjf�f���}�}l�<�k�-�s@=�f�gUZT���(�2'�yzנ[n�{��w6�B��%2}�X�}4�,*�d�����Հ{۵f�4����('�e����I�LO�n���$�H�0��BH�c�`Hж2�(�sW@�p �YH�CDlXB\j���Abi�B5�VSB�Gq7�JZA"C�=�u|�0��"��D�
�%� E�HA����!�$�k6"B0����i 6F h5��1�jF��hXB$a'"HRi�m��JFk
����{���0e�$�XB	�D�X��\SM>a�J�� � �b0*���X=,~|R
0OO�N@X'�� ��
�ʀqU� v ��}G5���ٸ^���U�	�'2D�x�����X����۳a�B�O�}�����?�O[MD�$�ɠ[�Q�yzנ[n�{����!91��cǠ�ܝEy�@�X:�H������5�<">�
h�n<r)�!"�ȏ��߿=�w4�ݯ����e��ϙsUJ��sSU@UT�����BI6��`wo[,?mz��d���Lx�(�h�l�7sm�|�owM���j���U���F�nI4�Jց��^��n傸��b$�w��v���SR�55%9��`y�vl����~ ��=ҵ�w��6!B4��F�PŅ�����=9����v,�ں۲�b�����͛�$�$z����[4�Jց��@�\�Tȇ2D�x���zٿ�/Y���_�@��s@�/i�i��$��94�Jց��O��%��j�=��`ynj���S4�*J���5�y{��=m���l�;�+Zu�s2����uTMM��ݵ`rJ"!?gu~sk��~͛RP��(I*�*$� �XRy���fe��h��m9i����M�i�[o:�9�z��6��VgleJ�ZP�;g�M٢����mp��v۵���;Wۖ�$����+����8�q�2���b���w�3�;C�CEs�댎�8x�bn� 󇃍�;���v�7���Sƀ�=�ny��&�F��خp��T��l�j��!�S#UH ���{���|�|����LDa@mڐ��6�M�Hu�kX�\խ�/9��ucPX��&��
&1�`����l�3�[.���l�Q��wu���0|��H���&���Z�����z~��s@>��@3�U(�(�"r5�y{��=m���l�;�+Z�Σ�ǋ$�z������{�k@��@�\��ɉ̍8�)&h�l�;�+Z�uz���z߁�l3k�=����T�)���^+�Y�6瞋aCr����=[۫9D�Us���=���<͛ۻk�����4���=n<n)�"I�ց��^�}���$`ŉ#P���X����V˰34z��c�d�$`'��n�}��?bW��ց���@�P�QF�ɏs�� ���wJց��^���s@��+�҂$JF�@��Z�?ffFN�O�3��X�ݫ7)�;521�����^��sp���̼f�[��:�y���7<r�vB5�q3���������nm� ����!%�n�t� ���J7�H�H�^���[4˺��r�PO&Gi��93@3��`{ޮs`�D&�Y�}\��iF���I&0�M��k@��@�빠u�@�/\�ܘ�S�2D�q�˺�׮�}��3+e�	C�c9�T�.�r��J�h�<�u��W]�ݼk#�%8R��ns���K���lX��9LR@�������u�@��Z�<���:�,�Q�2c��*�`��=�W9�6}�v����P���kJ�)�M�?5�ywW�z����٠�sJ�Hb��)�T��B����`gwZ�ٻVO�� �
�lJ`l ;���z��g/�O��$Ƥz����	?ou~rw�l<͛2V�f��0N�8� ��=�����,c��&cq�n7]�k�ݜ0�dQA<�!$$� ���zsfl<͟�%�gwZ�<�qķ����<@�y�oٙ��������}�Ϳ���r6�$�Ci$۠<�6l̥G�D&���X��3`fh�K�$�5I�PMM��C�������@�t�hW��:�d���X<q�s4�l�;ϫz���}��7$ޒDGإb0"
�6�ȭA��@����%x�c�����6�]]HMT R�5�m���F�'F���05�n�:�|��q�s�+UTqù�+�FYu����h��5gpn7a�"�^ �v�8����;����%�x�T�#Ð�;g�c���y��,v3]k�@-�4e���p퇞�������&�v�g��n6F�m;TX�Y�0�[��8�m�P�v^�qׯ�s�]�IRD5I��3 Ή��f%���K��m� E�ױ�'�Lq��۵���iڧ�}�Y�l|�X�4�5XoWK�<�6ln� �nՀgUZV(�Cq�9�<�W�z۹��f���Z����J& L�5S`{wmX{v��/�%3����_����Z�9T�MT��UJ��P���sk��{�6�vՁ�Vkƞ���ԏ9&���Z�?������~����f�^����#m����s���ܹؖۋu���h���v�T�;���`���y#rcqO��I��+����hz٠w�V��+�[c�d�$�L�krO>���
��vU�<�~�����ށ��^�֡d��ŉ�G0Q��>]k�;ϫz�uz����p@��PD��"q�~��z_�����[w4�Z�:��p��1G��˺�����ֽ����}nJ� �mFԑ���d�[�0N��v�lM����d�>����j��U�X/��$��z���˭zy�o��|�����{��C�J��n�A�R�2}��k�7`l�����W��H��)��SI�jG��#�/;��	��ߵ�èE6S��@ E�`K�c!��B�T�A�$��$aĄ�!D}����j�ן}6�櫩��3N����N7�y{��=m��>^���נ^����9LR@#�=m��?�FV���}��`y�6lٺ�������ŜIWf�ڍ%]�1�D��l�×�<<��c����wͷ������˭z��������+�5UNj�����vo�
"1����֬�۳|�`��K颦F�u4���=�_�@��s@�zנr�^�}��u)��d���@��s@�zנz}��%$�D,F��;7ܜ��-R�ڒ0RL�>^���נy{��=m��;�]hci�0��d��@J2���N;|����6��X�'���u����z��\�ȱ4�U���^��[w4��z��͍ɍ�2H��z��������^�˭z�+�[cqd�$ R=�����^�˭z����B�E 6(�
9��ֽ�Z�/uz����ذ�cSH���Ǡr�^���^��n偾~�-\(�B ���B1`q`��@�"���&����O6�
B`tB��D&�0H�`�yhI�m_	FM��y�$�����!tL6!	F�F)p�5e����\	H�ȅi	4���&�]�6�0��h-H[a\ �bP)"K)E��a%Y��n�͐�Y�+��j�05
$du+#4�(F$&�~,E�Q�C���aX�!#�E~ 6l�E�s3 h  jM�   -�m    ]6�l$  m� $  	  m�        �am   ��@6�V�U���$�ƀ,���0{-́������Q�$�˳�y8s[�s��n�jj�WX"z�'VCMM��I�.SR����{ h��1{�N��=F�k*<��h�`      �[E�&� ��u�ƛ�1nSt�W*�@!l��;�Z⋎��Iu��\�JA��oB��]�(c�85�$YXܻ
��{\�,�=���ٶnc�y�Z��%� �ٹ;N��O�<�p�sq=����R�mdvc��TuJHLJwGO%6�n�1ȥ��vܜu�s�/]�����i���Uv�V4;��8��V��v�ڤ.�#<�n��ˮg+��6�(Vs�4�	ݶ@Ӹ��x�oF 4RI�л��W=u�.���%��������R���Gvx�\e�Y,v{�K������XNv�����;+n6��Ǔ�7�FB�7=���nh%�])�˖����Y�8S�r�#��9j�mu�!������U�1�^��,���������Z� ������n����A0�=jE���Q�g��mzXk�\V3�����l�ݸ���-j�7t�`x���x�ٔ�!m۰]X�\s&ki�ޜU%���u;�.b�!�����s���೸��ǃg]��P��B���U����vn�nw.�u��u���g�oA�rlZ�gd3�1us���vKn��qj���l!��Ot)c8Z����3ɞx��S��΄��Pv�*�-BÙ��v�Z����!C�+��n�4���*�hR�.�.���̝n,!d��n<�n^v�wfQ4a�9�A���K���@*켗`�p�0���3jm��X���O=KTnx�� 	��m�l��l6ʹ��lH -���Is-������������S� �@6��(��Uڦ� >�{�����������̫U:�VVU�V��v����/�z�O.�eA�!�㔞Z����E�Zz3��<�g'ZD�;<d�pc[/-h��2�M�4n'sn[kv�����`�]�]Iք�ɝ>G.�7O/H48���1���U����ڑ��
�zgģڤ�ksn�S���sg��c�c�V@�c*��e��n�5��m�Վh��\�+*���W�����{��|z�v�	Nf�/:�J�I�� v9�� �j�ל�����n��Ms�7��I&҈b�c�H������h��h�נ��tS��� 68��=z�h��h�k�>]k��f${��kc��dc$��4��Z/Z��Z�^���s�ǭ���⍸�^��.���w4s���͍ɍ��5"C��.���w4s�^���1^��������/:sl�9'.56p����n1�l�"�E=Y){���6��ɎH �߯�����=;����0���7��W�U2du�%�����~��RDHlQ��բD#�A�����{��wrOo�W�z���-;L���G$Zyڴ����w4��hu\�ر�9�c�-�mz�]��s]�BI�Ws�ѭ�@�*�d�Q��w4��h�j�>Vנ{����c<����^+&�䗎�:���[j�zsl��_B��]�s�v��w>�@�;V��׮��Zf����mŠw��@�[^���s@�}V��^���1��R�l��v��ՙ	B���L���31K^�Z��Z�
����Y1���M�(Q;{�7gy��w]�B��������5\:�)���M+��Z�ڴ����w4�T�Q���c�%�f��q��n
�\�4�2κQ���eއ/^�ӡ�m���s�h+k�=��hϪ��l����Қ��������DD$ٛ�j�ݝ�`{'u�`�N��SA2K��ٻj�̜�g$�o6{���߿=�Z�ǉ���I)&hϪ�'���䜿}��&�@*#�tp3�1����>�@�ԣQ5��n-�;���������Vd�^���7l5�uq��_j��6tdWC��v���tSG�:3�#��Jw�.��Zu�J�_�����f������Z�
���N<�܈��u�@�}V��v��mz�%pɍ�9�9&������Z����l�-�0�AG��H��-��Z���ٻV%	=��v ��K�D�Lsd�h+k�u�@�}V�����I��Ow�?_�����-�HR�ڶ��� $���2v��TmV�1�7��c=\�P8j��E�����0�#��n˷O])�����u��C��t����z�g��onc'����<c�� ������2�����gZ�5�N��S��A������ˉ�d�[�О1�t\"���t;a�bvT�a�hm<�je��bH׷GS��T�Uc#·���ww����{�϶_�����h���Ŧ����ۣ�\,��ݧ<���@�/J�=�r�v��D65#�~�f���� �h+k�>�ekc�!���5��hϪ��ڰ?=ݛ �����BM�]�t��j!�Lm��[���>Vנ����Z��͍ɍ�����9&�� ��hϪ��f�}¸��ӏ#$�Ǡ����Z�l�>Vנ|��P�hQA&�N��+�n�ͯ]����y�5�q��9�X�'�|�1�I?�Q�i�4��hu�@�[^�z�4{.�Q�y"�(��37j���ɷ)�)��H��U3,��1$!��q@�PcG���$�ZIQ�����˩�)a��� �ġy�Λ ��2s]�,ס��Q$��ԕUV绳`�ڳ�D(J�- �����t�0y�Ƥz�l�;�U����mz��j����G�I4��hu�@�[^�z�4��# N8A9��ۭb��[H�
w6�#ɚT ��6�é��z��HpQ4L�LMŠ���ֽ ��h��h��67&7$���rM�ֽ ��h��hu�@��\z�hqF9
G�������l� �:@tĀ�(� �Q�
!���
���V=ݛ7X�iSUD�SJ\�U�BJͭ�`~��u��l�/gat�G���G$Z�l����[f��>�v������e�3=��Zx���oܰ�Ym�[;J�^.Ǉr<�؍��ݒ����%'L������{����OĒQ���M �Y_�0ƈDFԒh���DDL��� f�U�~̚�b�wS�C#k$�?s��l����u�@�^]M$x(��@7��`�uX����V�%�I����fg����������br<nI�wY��f��>�@=���.��c~�9I��u׭q��n�+�Wv�o[-��v�i�ۑ}u����8y�L�僰�����@��U��f�}�f�mB�H����G1�$�>��h�٠u�@=���a��%H��rE��f�}�� �[4s�:���c�qI4�h�٠{�U��f�w9�0bP�����u�@�>�@=�� ������oʀ�55R�E=�|>| �qi���S$9{]�V��ݤ.��&�0�C���mn��v�$�Q�9�g���j�{t򽮗�,��ޥKe�N�x)^�]t#��k; ����=g�,�:9X��ʶ.���\�l\�i�ɺ꓊�g���8�;�7+�7m�8[ф:5���Ê�ڸ�˞�]�&�����\[�(@�ny���c#�n�w��|�n��� ]�qk���]��ϕ���tg�^5mƻ�I&N������f�(��:����l���@=���tQ4L�LM���u�@>�� �[4��h��67&7$ ���h�٠�f���� ��h�*�i�H��a��l�;�U��� ��4B�y'�DsrM��Z�l���@;���U��fa�'<h��,��T��1v:�`������n�{H.��V�L�i���l���@;��s�����F9�Nh�uV��WqP" I(�}D(����B�"@B��(؅q	%
@�۫����=m��H-W��kDm)&�[���;�U��� ����k[)SưRM��� ��h׬��f��tQ4HI1F��@=��`r�ݽ_�7{���Nk�:"o��g)J�K��]q��-�y؀�{qۣڮ�a�Y8�S�vH�/ez�k�b�O�|�����f��}V�z�4�-5�Фm	�a$��l�;�5�{�6�sj�"������*��SJ\�U��;��=��e�P���9�%t��HS@(�
�ݜ	��6 ��Dѣ.eICK� � �b�H��hFl�gl����6��^p8� F @�dR1�E#���Y�bh�L6Bs^!(k%e�h�˩���X��OVW[�_JmB�>��MƌS� �U��T�@_���� �T��G�`�Q�}A��}PC@TH*�m�]���{�f�Ͼ�@���$�O$RB9"�[f�}z� �h��hT�V5���$rh׬��@�>�@>����n �n6�9�2`D�������q�,WN莒��'>[�����q�㒊"6��@;����� ��4��hu�lx�1LxG�94���l��Y��f��tQ4HI1F��@>�� �����h��h^���NnG�I4�� ���`{}֬B�I�w[�;��kM�H�'��hwY�~����}�����^�@��X5��#��vً8"�0hd4�b����l'��d���<p�f�$#ǐjb#��rh�����hwY�[p��Q'�)TT�Ұ?=ݛ��v�X��XU.*Ơc��G�}z� ��4�]��mz�,V��X�Q�����h�����hu�lx�1LxG�94�u�'���3��`�uX�"A(�D�DjԊ������~m�N��&�@R�0R� �UO+������"m�[���c4�1���z^٪��8G���.��g8�/�Y>/�5Î�=��bꎻe��k��q�q��h��k���;��A�\��gF��zyӈ*�촺3۲Q��]m`��q��Xn�ㄒ:����ےŲ� ��̽���9T�:M;$r�R$�]��:��Bm�}�`ca�M�U�+/�����{�����~�~&r�Z����k`�y�l����m����sQ�S�5��:>�/]��l�BLq�&xW��^�@=����s@��1�0m���xܓ@>�f�{��{���ֽ�Mi�RH!8,$�@=����s@�{���Y�w��cx�LD�i�4�]���@>�f�}�@���$��F��m��>^����h��4�]���V���k�qL�LP�K�%8���ع��w/]�<\��s�5ϴ�;PZ9,%&5�= ��������s��B����ޫ �}̩n�2�[���'<��ߛP�X�@!! !E$�EBI+{:ՀowU�g{��Cggt��N�e)EUKC��sz�@>�Y�^�@>�Y�{-�G�U4�uM�+I(~�ޛ �oU�~�Y�w��h�sf9&�4܌�@3��`��=��VN���{zQ���������m��뗞J|I[��+㧡݌v\������ӦF�u	e�z�o��o�Ձ����DFH�U���tI*�t�UD���=�j�!$�<�zlݽV�ٵ}
!6wr�Sh���!s4.���}m�#?���q��4f�Ձ��j�׭�K�7T��u56�D&���`��33mXrJ�7��5k\�*F�*�rڒh��4��^�}m��wwww�����%�!m�tv�َ^.��nIxݳ^��.uՈ%����tt�����>G�dJc�H�
I�?~����>^�����ДD~`{7����C+�ә�&��T�R�??f��P�a�� �oU���s@��vb�`�#M�����l��ͫ>Q	���V�oM��A�]6�I �"�94�u�w]���܆�� �����E~���o�@�,�y�"H4�w]���@>�� ��f�z��9���g��C#��z�b�L�K8�����>�O���}��o�4I��J��]= ��4�u�w]���*��F4I�D��@>�� ��f���s@�{���YUŉm)&�}�@�빠|����٠z�F��dJc�H�
I���[}��_��?n�X}
~��<����4ɚ��"Rf���W�[f�}�@�빠ffr���H��nI&L�i���k�U���h�����ȶ�Q��I���#7b��`&�����m�Il杕x;p��u�zxm.�4�A[�Nw �	Ň&c]
�g��/&�ș�;'n���{t쵹gZn͐f�^��;Be:�k�펺۵{m���>I�.�e�n
��/a�ϸ}��$3���@+�RCl�S�)��i'�\�!wbn��GHt��P�5[�������s�\l�{VN���t	#��\��W�?O�f��w�h��:�Mv(ڒq��������h�w?�ϐyu��݁��7�I)ɠ{��;��h/uz��h��c�<�S$rM�����W��� ��f�װ���#RB6�h?f̀o�j�?{6�:n��`s���s�cQ(���f�}�@��s@�{��-�n�؅"���Qکת7S�ӣ�^���!91v�Xhnv�j��^1��ҘF� �#b�h��4�w4��g�%�ή,���S�2����s3rO����Ѐz�`�G�:�k߾z��~4��4�u�CqML�T�R�??ń���ϔ(l�ޫ���4Zb��pcĔ�q�ִ�{6���V'���;wR�H!H�rf�{�f�{�����@��s@��
��B�	��p�-t.!�#6�v��%����P�|�V5�Թ�;<�!#$rM�]��;V�}n�g���{.�,Q�5$#nf���:?fZ�{v���Wɳ_7��i1K*��u3N���`�mX�(�H0#�HEcE��A�! �H0�U�ID�vZ�3_t���t�)�2����ӥ`��;��Vk��ID�����;��[��0	#X��@�����]���֬�ͫsk[[�vl�n���I��v�Tz�a��\xvt��.Mϳս��Ʀ0ٗ�
�o��נ_t��{�f�|��֘���FԐ�@��M �����Z�ֽ�-66�!Ȑ�QG ��j��Nk��Q�ǿ}6���`g����1DےhϪ�>^��I����ri_���Q � �b�0�"ώ���|�3rO��$��U���9rE�|�k�/�S@=�@�}V�m��6!��x�(�[t�\�a�y�� �A`|���ył7<uO`Bۧ?��&5�=��Z�u���K���V��s��)R�PU"f��{�f�|�� �����Z�����?��5�I4��h޶hϪ�{��=��ɉ�F�ț�C��wU��;��=�ڰ�I>��v~��c��<Q�$��4��h������3{���'�BD$��
Di(�7�&f�V\KbF+�3Zֈ$��ɠ��":b�0���\5�	 ��ՑH�&b	��9u5�]l��HH�0��5����)�Eұ�B,@��!$V�+�H�ą�Ń<ް�L#�kL$X��A�1%�0� !�%�$�7$�ȕ��$��4���1��7�3	IS��Y  H�MR�p�$Jp�BU�@#M�!�C tP�N�w��w{�{�^����?  �`  -���  �m    [��  $      ?�|H �6� ��     -�@  ���D���5P9��X�D� N5;v��a�1�̘L�p��{td��mV8��A�5KHMJO]gb�nBk���km<b�j�,J(��]���:\��r�pY>.�|�fn�W@   � �knHI��M�m:F�� �TD�*�ϝ���R�
�rv�Meݝ�һ F4��nT�WWg�qv2�lݫ��lu�&x#��Wlb�Ί`�&3�M��S�#�s��f�Q#nݝ���/I�n��Ȼ�s��v��J�zwI�(v�䪛n7
�^�܊)S-����9��̨ncD����r�cN�ױO��ۆ���mp���m���&f��J��'M��D%� pݮ�t�̣Q���vz6-%Ӣf]�zc�{/'������.�:^�rb��Usi�jN�	�&�g�sY�����x�'<�7[��d�����I�N�c�\f��/T�,m.1�#�	m����M�a!t�6�צZ��;�W/	��{j���G�L��[Ghx�L����͵u���l�#�����1���/O;��"���\�2Y��^��am��\���Ćݝ�c�������Q���&���<6�Ύ�皪�N�5ź���9��ے�l���7�6ݥ�7g�{R��.�4oJ'W8ɺ��m�q��S7&:����|o��|w��h�G�`� mv�����lr&�Z�d�fv�av=�UuN�$ۊ�ڐ��*�8⁞�<ؚ�mUJ��]���R�������I��(i�kk�q��6Eq���NW����{T\J�v�sǖ�wS]ڂ�x�'d9�lq�b�0���cg$v�2��R^q�ۭY�-��_��� m��T� nJ��ٶ�]5U� ��IK.e�3333332�
� �4"|�|<4)]��}P����z ��{���2��)�-[N�-6��l@�QW��`�csÙJnnf��՗����Ίdm;g�7E�Ӽ�nذ����V.9�g��c3�:���>��g]n:�+��9�Om��=��33�:��j�Ɲ�Q�$t���E�v.V7>������������׉H���]v�gIv,��s`�#e#p1s�Lg=�zs'W;帎��̪�F��[mԚֲ����@��',�ˬ�E'��^�ƞR��m]�ݽ����rK�����gLv����W�,lQ6ߟ���hϪ���hϪ�;���D$b�'"�>W���ď.���y��@�Ϫ�:����F��9#�>^��������z��w���CD��JH�������z���@/�,-�Lx�H`�Z�Nk�?�/OoO�<�l��=+4ݶ���G5ƮH9"ޮv|���㧷j�:�ƻ�[l�AᴼF3{uH �^�@�zנw�U����Zq`����j5�
8���{��٘��}��̝�`~{�7ТCfwsSd��#Db�q����y�Z��z�ֽ��y�@�Q)��>�`~{�6��ٰ�
!�V�7	z�<m��Ȓ�-�z���^��}V��>�@�R�F�8���?�	t�j�V#�7c�q3��y����k�9�Oe2�m��=�t�cl#RA9#�.�����h�������J�G1cQ(����u�����s�2w���(l:5�|��*S�
�9����������nhM�,"0 5�
@R B��
D)�(B�4$MR�FLF�,�C��|�[�{�)�{�MXD"O�$�%4?������|��o��w�Ł�{�%ө%��=��^���̽w���~4����ֆ6�m��45������W9�3���;u�5�#/[u�5�d���ʽ'�M) G���M��M�z���^��M���n R(����t���^����@�t����cC$bn!9�z���^���M��M��.�,m�jH'%;'{����q`n���ơA�BQQ��R�D�)��� b��J%QE����`n�&�U�UcQ(��;�)�{�)�|�W���۔�4�m�r)#1�XD�����ڻx���sz��u�v	ϖ�m��z���x�)�8h�S@�^�@=m�{�4�MXD�I�d������^��mz{�4�)���#���F���2Jn���3����eig�	&�z��<�_�@�������$�����;����^��mzx-66�!8�E4�)�|�W�y[^���M}jвd�#J9$�$�m�-[i��o�Z�[�Ev �T�{LY]l.[��ͤ$ �'�ݻuY�s�W��!�:�/@c��� �zz�9 틻.�c�f�ق�텢��m�.��uŧ����%�v�=��@m���F�H�nm�3��Fd@6q�`��[���]�4��U��^�콯Pn@{
h��W�`�^��xk=��Y�j�V��!3��{�����:o'�1g\��FN���k`��n��×���LϿ��M��|��6��1�Q�k���=��`g���IDG�-�?�� ��Ka�	��绳|ٹ�Ł��Ł��l��u7��d�LJI4�Jh�S@�^�@=m��eU�)�$��Ow��Ϸ��=��a�(P�6��=����SBUKn����ٰ9D.�����~4�)�}ꮴ8�PR�ֱ=�6�e畇pk۴�S���rM{
�'T����}�����b�jc�΂g��f���M��h/Z�w\z8���e���3Y��'�{�M�)Z�@K�C�w��^wM�{wj���t���Ls@:�N��3kK�����	$�����;��h�j��5�1��UE���vlۻV�9���{�|X܀�)�3!R�s5S`�ڰ>P�,����������6�]��,�����R'�^N��0ݺ�^���F{v��v�r_C�I�%��}$��}����e4��z�l��eM\LX�H`�Zu��>^����@��U��H���f%�d������߻��'�}�niXł@@L0�J���_�l�W��D�N��ژ2$�z�l�=��h�S@�zנ{����'"QH�9&��>���DBIn���<� ��Ձ��k�X��sy̏hG�K���,[�7�q���{���d����z2��S��W��ٰn�rJ��2w��������#h�Š|�k���@��U�z��@�p�KxF�nG��f��>�@�}V�������&�R��:���ÔDC̭�`gN�??n͆����!8P�Mۺ��eM\LX�H`�Z���۳`�ڰ=��vDBY�߂�ˠä:֎�0�l�n�|��=y.ț�����݈�\ݒ:W��v�筺��Gݷ������l�=��h���=���M�L1�)�w�������Z�ֽ�nkq��ȔR<�I�{Ϫ�=_U�|�k���@��ԶDȄ�
)�y�Z�ֽ ��h���5U��q���@���`��`n�����`bĒ^�����)<ʵS�)g�VU�j�Wig\]1������n�@�n.��q�u�k%nIњzѳ�����"�n�Q>�m�e֥Z�ط��@1�Z�W;b��mm����݅ӳ�P���ѝڎ`�-vN�����9歞k��ű����π��[7Sl;�gs'ob�6�*���m۵ۈR�`� �y��k@A�R{5c���[-��ن���������{��>���;J2��vK�R]�bl�Ǯ=�Ջ�zK8��8F��2�WG�ՠ�x��܏�>���=�}V�y�Z�ֽ����dM�LJI4{k�7'5���f�7sj��Q�r����jUPL�LӰ;�y���f�-�4{U�}%� c����@�zנ�����h��@��pF�I�2$�zoY�}�}V�k����s���`'&H�Q�ϵ=����37nI�g�M��I�ϟ;�FxUwo�Z��D�ٓK�T��I����D�����}�p��4x8��,q4�
e*���;��lP�5%	)2w���f��y�Z�5U��q���@�{��z����_U�[p�KxF�nG��Ŀ~�����-��h/uz/bT2�ȞLi�94�Ϫ�-}V���W������ؔ! ��4��$E&�k�<h�'E�Q7���R=����p��q' ���>^��޳@�=Қ޹��d�n3"�h/uzoY�}��M����n�"d��T��; ��U��}\Y�*!F��M:��h�+�!����b4˨�a�
FI!��B`B	�aB]h�!BR U`ͳl)5*E! �;R,F]�I+� D�aRz��@�:%������P؇ Yd��
�1!IM�B��P4$+��%MCD�.�kDa�]�C�F�֐SBBU��GhB�
Ɓ
B`�F�
�X`͛�Ӯ&1�D��d �� �� �4�B2�ˢ!!@�f��C@B���=6i�H,X�����0HMj�n���D�,)|f�]$ր��1c���!�$��4�B�M�%
-2�o��&���X$`B,#)��a@Jl�Ag��T*C��`'@��i�?
�=Q
|TC�8��x���P��*�C� �>Zճ��˺������(�y*��9?,������`~~͛ �ͫ�R�8�q�d�4
�W�|����f��{�4��*�hQL�	[s�и�����8�o2ng��;����V5��跶�K�9�%:�~m������`���>�t��U��h6xF9����f��{�4
�W�|�����P˒	�bdnM��Jh^�@�{��z� �VT����8���U����� ���;B(>�*#�G������M�~���y2`7#�>^��w6���ZX�6l��[�@6z���'�[������6�[���!��vyԽ]�.����om�����?p��`~^���׹��
?0���;/٪G'"QH�I&��{�4
�W�|����f������'���A2G��=��@-�4��)�ZcU\H���H��@�{��z���Jh^�@��s`���c����_[4��)�U�^����o{��������:����(�m9�m�JۍZ��tj���B�	�1��ֹ�WYRB+v��6=+i';tWn�^�S�R����o���g?i�F�yz�S��aC�ǆ=�kr�����l��/^����.^��X��th|��:4�c��Kvn5y*ҝ(��0�}�miNr�m�;e�y#b��)�gK؋:��2�����mjzH����[��[���Z8f\c3۝�����N����̑[�QoQtvNG�@N玩�<�ua�S"r|���hwW�|����3>@vwU�r����̢��T!������� ��hg��hu��u,s&q�R= ��f�_[4���{:���?+=�-�$LQ�(A'&�_[4��w4
�����h���GiƔR<�I�}�빠�f�}�@;�� ΡP��ci@O�}]�9f���Wtx�Þ�u!ur�q�;��q���i9q�ɒI���h��V�ݮ�Q���oZ�;E/�&�SEkW3SW5��$���ٴG���CJ�"!�Vo�1nm� ��Ձ��j�%6�LuLm�U�{{�����V|P�1#�_�@/_�@��6��x)��@�/]� ��4��hz٠*ʇp��DHdNf�z����4�l�>��s@���`	�#o��uX�� ��ޯ<�y���nնu���]�m%��3�2`'��h{����@�/]� ��4��l�1)B	94�l�>��s@�^�w���ռ�#�QƑ$Y�@�/]�	��ߵ�ZA����$E�c"H�!$X�X��BB$HBA"�FX"T�$@
(:�h�u��l�=�'���0��j�X=�v��U�{{���(�
'Wu�`v�_>M��i˚�	���̳@;���S@�^�}jh�)�����`\����&wH�om�v��v��yr��k��i�9Z�m���@�-��<�W��f�U�m����T�JsU`~[���(I6c����?<ݛ�l9sG)�'2�U2�U5E��w��33jΆ���l.���-�,�L�H����N_~�[�p���nN�uLA��%�
#BH��_���;P˪�#��:(Iɠ|�נ}��h]��wY������3��Xy2uǮ�ۮ
���{�x:���u��08�[T��^�W��!��G�}��h]��wY�|�נ{�jOa�!�a17˺� ��4�ڴ��M�ƪ����6�@�@;���v��S@��@��.l6��r1�$���������.�����ٰ�ڰ5�)�$#ȜZ�l����^�wu���Z����,�H��#�R��ն�m6 p��g��|����x:q���Ll V�e��6-����g�)�����N�����TRt����Z9�����<N��gѼ�׮��Y$ �=m��`p��ِ�d���J��ň��3�����u���.�pg�q��'v�]oSl�N\qn�Gz��/X6R��m�4a�Xv�z�q[i�{uy ��V��}��������|;���c��;�v��=���5Ǟ0$Lxu��4�+K��F�;^�sM�"C#��9[��wY�}�ՠ}l�h��s&q�I&�[l�>]k�>�X���h�\�F�'1di'&���^���Š�@-�h���4�H�USa�D$�����n�X��X�mz����&�7"�{��m��ֽ�e�@��X5�Ե��v-s]��+���4�gm�r�#��)��.i�dX(�$dl��)&�[l�^�@��b���@��͂��)�������u[�
�$���\g���^�4�f�Wv6��ǊF&F��>�X��l�m���hʰ��$�9"$#�-ى$��uXwuX�6�۵��n�:2��jDMUX��X	$�����~�@;��ڮ�j
Iִv���V.\��=�mk\G듚���mnk�O�5� )�$����NO�;��4�݆�w���Z�{�y�G���,�,�I�}� �[4.���Y�_�=�8�y0��I �_�rO��}��O���OVJa$�DDm�X�ے���z�27�dh�I4
�נ�����a��;���p��$�*�������^�4�� ��hu�@��7��l��2�s�!L[�)嗓��㡞.�l�����n��M;v��n�����<W#���/��4�٠�f�^�4�X\t�)"$�H� ��o�H;{��;w����nKم4N��:@�fI��f�^�4{��@/��qդ���K#I94�Y�n�����	�J:�p��.�fV\�"k�e�(�JCJ$!i@&�1H�H���Q(BXE-�e,e�]a	[I�em�#	�5D~D/>�9��{�kF�f�$b$��h�]f��~�O�:��4�٠ܿ�\S�Lx�xA���q��ŸtGӎ8�={])���GVJ^�F8�y0�rH� ��h�٠�����=Lj��
<Q��(��1���D$�&ó�����73j�(I6{�WC�eD�HL�M�vwM޷Y����Z�
�0l.J%JuR�UV
'���K �ޫn͇$�&�;��7��)�nfJ�d�T���V�I%�����	�{��7$�* ���* ���U�Uh����B�
����*��U�EPG��T��B
T"B
�P�B(�T"�B 0 �P�$
AP��EB
0T" AP��P��AP�
AP��DT""0T ��T �� 0T"*�T T"���$ �B*@T"�U �B(�B
�B���T �B��AP��B"0T 	P�� @T �B*B(U��T  �T"�AP��P��P�B $B �T"P�,EB� �T �P�B B0�@T"�B 0��T 	P��T"�EB �T"$B" DT"AP��P��P��P� @T ��*0 �T"�B	P�P�@T"�$BDT#P�P�P��T"0,B�"��0DX�0��T �P��DX"DT �B �T"P��Q(�B)E��T"�B	E�1��T"�DX ���
�*��
�*��* ��TAU��
�QW�D_�U�TAU��QW��D_�* ��* ���b��L����j�W� � ���fO� ��  ��*�@�(R�����C �!J   ���     �T( �BABT���PEIDU�H   �TH(U$� TE*���QT S�   �$PAA@(Y�i�D��qS�ϰ=g �^�6��NCF��>N��'p��L^�޳�� �9t}�����</��B��LZu�A���tj�ٽ�QP	���k׸� � |�      c0U��g��\ƭ�;t�t<�R�t�������VZ+�s ���������ۗ��ͪ���U�<
$��V[ϱ׎�s�x��|�U�(;��,ULڼ�q�:���zx> �R��(�(R�0���Sͯ���4�6YA@͔�J/� �J3e(J
S;:)sҔ� (�JiI K1�� �,f��biJt � S�vtR��ʊSu��bh�P� )N���J
\Ɣ(1M4���R��9
  A@ ,����(�Х4��Q=ɫ�n�]��9���G��<l=n;��`"|��^}�| y��y�|>؝s���{�!���E�L���͗&����_x�P     N, �>�Sݜ��]���7^����my� ��[nO������^Z.ۙ�� Q�Jb����  �}���wɃ�< ��P��������'�{n!��T}�6r}=�y:�g/</� ��ԓ�*JT 4h ��51JU4�  "x�T�jJ~��� =��#�TH  *����کJT   "$!�*���<S)R�{����U�g���t���2�%U�^O��IR���5��� ���QT�x "��  EW� X����b?��!-`���0Ma
�J�lJD�F���9B�HBBB!!�HB$B����O���]1��0 � �#�@��H�$6@�z����z��dc?ϊ"䙲�q�Ƙ�lhh!@Ő�D��!$W�# ��r,�2\��/5CDC~- H֡ŏ��2y[H�a$��zn:�&�sg�VB"@hB���<�)�==�,�!��G�Hҙ��!�RA8ٰ���I`�ߢ�v�>!���$J	 ��"�Ԣa$ZQ���8y��܁#M!#�6V"�%�H	$`�}�|>X� ��\!5���P� � X�%���Mb�̏%D��q(�^D�5y����4n����qa[�h�~a���	A�<=+͜&8x�jfs+5�Z��ﯾ? �H���RHV���
8k4�!�F����I�$i���dz!
QI�;̵��R�n9����y���1*f�X�h�H��LB Q�`!@Ģ9�|"��ą�����Ҳ	e-�R�^O�+�^���(&)R����#�/�)���k��k�_<�Ņs[S��	�S���h0!L�F�4;xž�yy焐�8F��M�.�ۂv�Զ5t��k�no,�Ӣ��Q�J�OHRL� �/�]���v{Ւӿ5�:�J��*w8�
���(A*p8�sӌ����N<�4n����Y���q<4��h�[�j�f��c8y�Жms|���T�crN�&ҽ�]�AX��W�2Յ*�ң�6$"R��������V��G��«V�����~�r�zz�5:�Ј�W�y�$�U�|����ĳ��`�۽p8���`h��\�6M_rN{<�$`Dd�5�
0V8����3d}���i ������
&��V1q��!�3h�����ןg�<��"w�<�y�Ħ8iwȊ�6�%��6B�ͷ\ru��i��&�8���N��ь�C�!�$�LѲp<=֣�`b��@�a�J`B�B*]�0�)�
�!M>�$4�᫿�x�XB��(�>F%�F��ƌiL1ӣlHŹ�۬�٭l�@�-p��� ���.�#\1�|�x����@�tB�F�l�U�.iѱБ�:��.��7���4�<t<UN��R�#��M��~J����Q�c��Lvyy��4��o[<�sy����͹�Ө`��<Bg&����sIL�-�A���5`�	!/! �$UL` PL@����s��}	_4�"�2HDR���3F�l���l�B4;�J��X� b�a�2�470��%tC���1�a�k$����0��q��&}�u"W��Rwn	�G�؅��7O��\�4x�lJ��Hp��7K��k��Á/.��O�^xx׏���_�;����`R4�f�m�x^r��g3R���+̔����d�T��Zֳ��0��xI �_48
a��8��)�����������vcJ���P�	Mo�����y�h"W�rI7�
��$x�0hc�_
r!L}4U�BJ�6�\* ����6�����	���b�Y꺩�!f�Y^�D�ۙ8���-d�!���Q��ԀŃ��`��p�Q!K����h"\֌wyxa��tS[��a�!LјM�/�.��a�#L�&�O�������@�T�~��^�[J�H����պW��m&�X��g����~�����{�������\@�%�U�Vb�D�%K=�[���5��hѲ�>�lkSA*��@��}*�Zb�Bɗ[���@�+s�R�u<3I�������f��6z��#�ǁ��@���gnDi��F�|IIAt`��Mab�Þ�8�l@��"b� �X�����WF{}�Y�X��i-�F$�Mj����?(&����=�s�Jb��*�D���rJ�k�k˲��J�}�¸nfp���Z`'	 ��Z��5羸�U�U���!'F�I��y����ߗZ�z����"S��c�l����x�;b�Ʋ&�\>�d����@�-������Ly")u>i���؎���&�-6���b�)��3π����Q`���{�)��&b�׷�g�x4`���HaB��q�i�1�	��jm(B$m!��6�aL4���)I��lч<=e�)T��*/��#�><�<&���7����0��=4<5�>9(B�
`Ǝ2�6,i��Ja$a��`}͜a��B����=d5�	G��)�Ç����3^g�-9�B��bQ�D`B��$%3Z��l�C�����|�UW����k����򷾈�orɝ̫k��脯��U�3W�l��Jo{�<�.l0��1���5�=������#�q!@���	 ����"D�D�1Ӡ�<!�%�h4]�4@#,�kM8rIkP0�f� p42�4�����{S|7ō4<[�Ȝ��k���B�[� �>��J�?}�O�x|����B@&�ˣ�����1v�(�(SZ����MD5�����&a}���3f�0�kK�i��aL4xa+��͜�ȵ4}���	L�m��{��Oq��[�NlSs�;+�Z�R��)�)��<���)��S��bmӦb�~HPA4���ה�a
bc-?B�M]�!��i��*��j��:��boަ?Z�$)�j����mb�<�!g(���ӗJ��&���
i���//W�6�Ր,�>v��%	���j�[ږ����,�fN����%;Mשy�o����~��%�V�5�>6�
`f��==���H$�R@�DL+Bۯn߫�(����Gw"��{1�7V�9�.�c����3k��5J	)S�Q�]�^U��ʚ��#=J�X�H��"i-^η^Uw�T�!LU)����ɣ=Xץ����!6�4$!�k۫�l-0���4�[��b"B����'�@�}4l9�Ja�a�>@���j��&o�8M��-Hl�RG��u+i�����!}���7y�3z�A��'&QVZɑ9�Z�6�m�s!��X�0�7�燦��kg2>��H��MӞ{�󏤹���m�
My�����J����MM�Z
D�R���F��@# �D4�c�pt�K��b����D7�8zz�h�����P��ў�$ ��7��IsNÃ���i����C�0�"�s2]�c�6k����$@���p--6�y$$ BS��#HU0�jl@1� @�$bA@�	
2�+��WA�ME(��"�+�M��D�*n(���B�=P�G���)�D�	H�P�d`�I#FX����������!��A�R.���3$H���a3�u�����I!�@�)O	sg#�4�y
a�!\Ԑ��� �X���`@*F�[Z~#>�S�&bd���X�,H\r�r� l�2A!>�%:��L�^ytl��H$\p�$�1"�d"�_Tt���O�ʕ�1��`F1�%���Ja��8��!���I1�U�Y�s�xB4łT�ň�}!���	�D��
0���]3��v��� �5� �z4DH�0E�#�{�HS�o���Y��>�g'��`D�DB� �F�֏�[&8s���dLxA�jc��	��1�0�`aq�,��H�U
�	![*�2e�3��{��=�]��ےFDI$�P 8-�a�v���m@]��Ԉ5�uȵ��!���h                              l                          � �     �   �                   6�               �                     8    [d    @ �>            l   �`   h   �>       t��`        H  �                                       � �|                        ��/ZR�	:@8  n�� ��դ��m�m�	 d�ٶ9n�  6�-�e  n��	�p�   ������P�UUJ���e�  mʐ �6�Θm�`Il�� ��m�[@�d��r>�o>491�6��`�h�8U:�\��G%�B�[��$���5��e�@Z��ꫂ��E�*� � ���8��^p�V�bIKE�-��:F�9��E��m�	 ͮ�Y��ې��
��*�A����]0 [`��6��m�          �          ?A�m�                �`H         �n��c� l�`     	��hm��u�6�6�Hf���3lXk 5���u�lҖ��fհ�  �hA��W-[@  .�� � �iy�Q�V^@�ʯ�ʀ��-���i��  6�v��i�� U*�����%��U����m�mm�   uy���R��U�U��R�|�1:�%,�ٴ�m�-�����$��`' [@��[�������~���Z�MS��j�Wm�(U���z��ҭPY�T,<m ��mfFW:�  6�m���m��    v�   �	��޼Im�6�[@ $����r�R���igKp 	o]��^�`�`[A��m  li�%��:hm[�m�$�8�뜵�ږ����[F�j�Ș�
�k8ر�^^\WQ}-��Y�"�T�,��d.���QPcʯ����R ��Jn�����H@=t� ۶�ݲ�RZ���)��/0T��J�$����2@H4�i�2sZ�Z�lְ �볮֍U]A���)�ԫ*�P�mp�l�d1��v s\��v���[��U� E�ֻ��kXH ;[!Ŵ��BGkg��kxݰ9��-m��jUj��K`-�8�]�v���[gK�M�HH��j�U����ݜ�����[\^�v��m��%�%� 	�����;k��v^@N�M���m�����m���8.�g��*��t���3UR��\lh�ڧB� �"�<���u�`h� R�e�7o%s��ڶ�bb6[g���g�J�6�ŨU�d�U��7�FPR�;tݱ�N7iTe�j��d_T
vH�Y��"
K�>�F�N�ʨu#T�6�����T��m-*�Rnp��fW�淛�S��	�޽��2���ā�9)�	ӍQ���I�9�#U���­J��z(^@jIj�+�� ��0 ���-0,U�M��k-� m�'l�ֽ��cZ�!&����Xl��u����);5W8�m�mU�R�^ݰ��Ql�1����$T���,��.��٪�^f�.�[�Ɂ�7�PUEgll�!2g������΍�7[t��9� ��k��]r��k@	 �6s���[��i�ܖQ�����u����3i���nX�=�� H��d�ʫXL�e���� �Nh�dv��[p8�m� -�n���9o[iAW��v�]p9��kX���}wKPk�k�u����v	ӄ��#�����x�����$Ҷ���t%썐 �sm�]nז� :�ٛm��a,��]�-Y*��NM'�[O,��v�ԫ�
�U�y���Ó�U<�PP�9��z�m�i�Y�Ã�ӗX�#4���-�p  ��sgf�џV2��KS����t��媠&mՍIһ<d����:��屎T�����w���-�J�y����̟�Q�m�
��v8j�'���{m�j��P�6�4�\ ^�V�ք�]��8Y"ҭ�K5�n;��m �I��i�M�� �!v��vݑAn�$5V6��:M�y��#6�L�bF�3	@$�p�]� 	 m�m%���m6,c����m�mz��4��g9,���l�2�   �mvKα�r�`���[@ �`hHְoR��\�h�� -�[Cm� m�H 4� �o$��)k�+VƖ^Hi�� 6�Hrkc ~�>�`�` ]*M�l[@s�-���` H       -�� h  �bZ m  �kn�Ye� � �m����L�zkb�Im -�p\��;�m��   	�h�a'c� A��g �[%qm,�j� @�am$m�  p.��!#m&��ݰ��  ���l�Y7T�0*C�m����[�@UUR�J����ʺ�c(�T�8�nU���s�́&�i�޻��m�:�@UUM����(�����Rv� :��n�;�$ְյ� *���S.��ٸ{6bHƥ�����m�B��/6�+cs�I��.��:��'X�+VS�Ã=ʡ��۔ l��]qr��σM�ThV�Wf�y� 5
�+�˓�j�WB��l,�&j9�z��s�%�벎�ێ�+��[�X����x	���f��m�M�S����t���mb9��U*�Ue�j��-�� ��A\��X�F���jP m�m��[[\���Ͼ��I���dwgu�����'���;rF�Ʋ.��V�x35[Y�6��v�t�ult�r1��4]��yr��x�,�7ϟ67��qy,�-�̵%ěmK@WuUUR���<+�#�z�  Ɔo[:ثdM����m�<�����Y� �Ԧ��Y�����M׬����[mN�,`�j9�L�l;�S�ؠ:�"�#E��Ƕv&BM�j�6YX
�Zٵ�ۅ��F�]uUP@��ʃ��j�$^�H�d-�m����f#U�[v�F0Q�j� ��C��뭸�jN5���U�h㦚j�}}��H�K'T�(��d�ٲ�rAm;m��� ��-�5�N�ۛqHn��22��+m��m@m���m� ������v�Mm	�*�C�9i��n8��H�lI���  kn  �n'8�n�v��V�� �` �Duyo\]6�`�`m�����'>��z����mv��6�[�m�ۀ-� ޮ�`8��k��[f�s��m�k�*|����jL�!��T9I9�e��Y7m�qΥ�-���(nC5mWG	�P��4�o%�R��r��j9p�nڹj��ui;��^�$	��K']�IkH��[B�Ӡf��t��� �R �WK�tW-���SST ���ڒt�  $�;Y��  ev떰6���µ�[A�m��6e��  � ���v�hׯ0�N���b8 ��n���^� m��m��s9^ɹy�
V��X�j��Xk�^��l-p-�"�4���Y�����<�a�۴��5�x�ȥkX�aѷ��5��1J Y+tݰ�{h�ڪU�U{phݤr�� 	�^��fӴ� ^�K��m�� �V7k'YF����C��b���`  �钵PմS�)V��[����/��� ���\xN.y�Cc=]V� �t���Ji�7����`�r�m� -�S�gj�
��n��� ͠%Z�(�/�ʵ��a�^UN�@yvZ�������e*�q���u���۳�[]m�`  m���ƶ�Z� p��H �m���I�Mn���R�uU(�jU^Z�V����ѱ�p��ʭÖ�eB	햪���8� V� ��ni� -�Q�l�!����|��HmmlB� �&E6p���7Z�n� lB�� ;m��n��$[A�� I��  �l ��
T�h   m� �  ㄀����m��&vZ�-�U���.�p���8�ݍ`�[@ �vM]CZֿ�*����"�!���� �"� �z����(� q���H� +��z�z*�U��Q1E�����'��ɰ\9## �Њi_ � ��_Q@�x#�A�Pt�At�A�����H�I%��a�c  Hŉ$�`H)6*�}P[��S�]D@�6(�� �b��� ��x
 8����.�h�� �0~P6��*��������O@^!@Z��@^*��IO�ā��`���R�IU��!� �_x |��$R/_�j��AdP�XA$I��"@�*�d`@�>(�@��E`��( ��OAv ��A� �"H# �D��T��><E6�������@����x�����S��-T]!� x�Abz��
:E>�E���)@1S@�D��j��|@H�iW
�qD�m�������u  'PD()c��{����wvO�4f�yX     � �  ��[B�    ��  ��[A&�   Hl ���$     h ��    �i� Ŵ[R��vyn�Hs�P
��F�Nn�g�Wc��y�!�M�%d)�N�KM�l�I=��l   �Ѷ���[��[E��p컆��iV�M��+B֣J�U �]p5+[N��1�����	�gP�TS��Rtb�v�K�v/5q�p�T�Xb�ƃu��/7X� �{l�ηK��Ž�<��i��N�hip&u����5�(�A�ɽLs	�='&�m=���9�6՛\fC����]��{۰sYY�
�!�؊bM��n�u�����2ݬ8E��'=-���B���N��U�8�d�;=p��b^m���<��T9a���v<�MMֺu�WX븠3�2L�ǆ�h'3v��:�nh��a��O��;/\��cZ�Ų��a�n��Dp�2���(;k\�zyz�Z^:�Z��۳�9kH䄍���m#�ўb� �2�m[L��Ѻn[fUBj��ayMM*���I��p[�cZت���[*��q��E��zwc�-ۻ:1;�K�-�A/'i9]�����̖��Ǭ�;%ї�%�]8�v�.㮝�u���]��z'�kYWמ5���n��#v.		���=b�Cb�]�<m=��� ����֞��'���LW3�M��бe�D�`�6��{��	.�+1�s��ӔA��Xt�����c��;�.�q��=N��\U�	t���ɓ=�t�q�t�x햫�M/���%�\Ig�狥w�k�E��Wu�v�a������5Kq�.�*����[l@��Sq����qs{eͥ��M�n5Ա�k9� ��Z�^�Y"҇m���e�عf�� �F���dP��֭�:Ax$���]��������⃵4�@<��T�D>@HL@�"D~����$�8�ޭ��vͶ��nʕ�ͥ����]t�� lԼ�́F�JŬ�F�'S�F蛍����\v@���]��\\h���!X�wi4�ڷj��t����9���phqv�b�v�bڀ�	W����9���\�j^^h�z�#��;p붎�Fvs�ų��{=�.�ɀ�ɤK�(��]r��cn���qQ3U�]jMd�(��P1G��fe�[���/��1����9Wnx򋱸�{`=�*9Eێv{s��y�ڴ�����@:���bx�)��"c 9"�>����uz{��>�j�>�c�H����䠜�˺� ��hs�hR�� �n�	�$�"nG����v��[��ywW�}��s�?��0�M�v��[��ywW��� �}���X�]��O=fN+���ƫ/v���V���5�ne4=��
7�В6��3�E"�>����uz]��s�h.�D�J3"M8�4.��g�EBQ�9B��*{�03k�X㹦��ג1�?��q�wW�}�1��ƒo���\�3o�יvH
��L2G�@���@���h]��wW�}�'����1��hR��˺�����ڴ�W��m����aK�uX5�b�7���s�݆ݷ="6��3��nJ��f�Xn���ޯ@����v��u����݇�O�ǆE�@��^��;V��:�h]����֘a	�q$z�]����3�!(��RP�%	����m��UZp�NG&E�C�BI)ώ�Ɂ���0��`{6�`yw\j%�&�@#��|����Y�}��>�]��W��rF�Lm������z �n����v䰶a�m����m�8B����-v�,ٙ��o����@��)�}N����^�_+[�#8��I"�h{�4��s@�{���@��O� c����7�`zsz��I%2}���3z�����,��s�(ә�|�����@�m��rIB���i�r�D�rU5u�E�@/����M���h/u~m��~�}�R�8{H4X���d��r���v��㝭nc���>���W[M2O6�Z�t�+�8�$��=�~4�+��|�����@��NEb�8�%4�+��|�����@��)�|��5�ȓO D�h/uz}l�>�Jh^Ws@��Z�F7&J'z}l�>�Jh^Ws@�{���ո�-,�RH��ݘp*J������.���_[4{���$� @ԂG-�m$����G[A�'�I���h�M3D�9��i����L��nN�����`��;<=�B�<=u7�F�6�1�q�k���[pf�8�g�y�*qt��\v���%�����i�u���m�`��\�����\�9���-Y]fE|��:V����۠r�Q|�zE�Z�����8".�����5J�{������w����n1�{f"f�j�]U�vʓ���V�u�.�z`���ع:&���Q9eE��~�Ǽ\��@/����M�:cQőSr���>���R�������N��w4�v	����q�G#��cٷ�ݳ�0=9�LS�;S�@<C��I4�Қו��>^���٠yuU�"�19��ו��>^���٠}��[d��*n
��#��sq!�-k���ú�<����ܭ��q܇L��]� ��#�������0��`{6��������?~y����pqǠ�����e���%�)d#�, k�ck�������HąZ�P"� ]�&��$�a4��U�������ަ�;\�1��&$�I�}��>�����W����<tg��;������ަ��lf�vX�7E�9��i��>^���٠}��/u�hn*=DN'"q
rz:Ř͹ݶ���b��#a�����{WX�m�{t��g�O�ǆE�@/[4{�4�u�ֽ�r\�L'�qI&��t��{��@�zנ��˪�9A���Ȕp�/u�h/^�$�/%��DU�큙��ӻ�q��k"M<���>^���f��t��{��@��Z�''�F��@/[4{�4�u�ֽ�}�>���6{��3a�Kի�rZi�WD�Ҭ����U�D�.F�`���fu۪����|0;w��NwWВK����{��O1�?� C@��Q�|�k�����M�:c��E��󉸍��^�^�h�Jh��g 1w��,�wW-
9w/��I$��ݜ�ɧ ��8�R�IZ�T��������f�8�$�@��S@��Q�|�k�����چ4�qX6�F�|k�ؽ��5�%��'�5:E�:�xt�t����̒,\�i��m�������4��zz٠{�)�|��5mA<�N#@�zנ����M׮�@��Z�7'�F��@;���Қ�]F����@;�W"�Z.Y���8�����4���3�|�f_j�Sy���w6;W��J�@����Q�|�k��f��t��fe�q5T�H I�&D����'ͶB��/Z��Y8x4�c�m��U����X[��������̼�ᗲ�Ǒ�G\�c�p�����A�Ӗ�=�v�9�N{���:ސ��fp_��>C�ݲ�n��h���jY��P��5�9+)\gt�z/]s�9��g�����Q�^g��r�u֞j��ӄ���gu뢳�;�6��f�-�;8�;����wf.�V��Y���ױ������)��ݨ�K	���=].�y�W��2�[�g�#q�߿= �h�Jh�us����7�"�Ǡ���f%M��M8w7��?ٗ�1>��x��"x���h�Jh��4����^w��?+���*�M�1�$�QÁ�*T�3~g ��k���|��À|��5ƞL��h��*�^���M�]F�޲�ki$��7M���3N�u�%��%״�sn�N�a��b�x��l\���-���o������Jh��4����*]c����Z.軹`{6�i+P�%2v�9��h��@��O1�?� X���r0=��,���o��X�6���s���F���U�^v��t��{��@.we�`��x�%$Z�j�>�Jh��4������U��]V��f[�����/Ml�D�T�N:�{v��;����E"�>�Jh��4����h]Ui��?䜑�j8h��7�f&�Ϲ��7/u��va�IU6~y�������4�dN#@������K�٘� �� iL<z M�"l����R�3���p�$��p�����l`�o6p(20��<�9�A���!�q�,0�G�M_4B�&�$�`B`A&ZD!3^mҍh�F��H�!R�چ��4�,Xp7)����H�$6Mj�a��#�(.�aO!F(j����W	LޚZ�Z9�a�h�!L��ʒ�Փ͉�4B�	�������n$nA�0�H1B���#*��0��[�r\��l�n�S��	� r����ѻ�p��À5Cm�m���/����o������f�NJM�ٽg4ԛ�����.9�j�ۣd$a	p�S3#(B,c�*d!R`Ĝ�؁�t�����W���Ȥ��!L@!���A� hA��<b x��b��X���!�@�i�/��}�y�������4���I�����yڴ�Қ��@�ʗX�cj3&2H��Қ��@��Z}ͤ��iH��X�%猉svm�4z�.�˫l�.���gܦ��<�S��2 �4�u��^�y���UU��ɧ ��/Er����q��h/uz�j�>�Jh��4�p&_��7�"�G�^v��t��{��@�{��;$�V�2'�q�ܰ=�|0;w��NoS��H@z
�(��@�(�Qy��@�x�W#�NH�4�uؽ����@��2�tx��i=�����Zuس���i}��ig*Q��r�����vd�B9^��6�O�r�v� ��f����g ���n�I��D��@��Z��M�]F���W�yeK�rcr(�`�$�����ۼ�`zsz���,m.O��d8h��4����h{�4���#o���s���F���ܾ��V����4����?;��{���N��{����t ��!n$��^�流mH�6٬�d����`
��W�	��K%h!5�3����q�Q	vo<ն�[�y��s��m/jܝ2��wh�������G]M�&��\i�k<�3e�a�v�V���%���]��]�_d�9�zN
�4����.�CRr�m���,�\�n���礋ce����YUԜ'����Gm�T�
���9���[u�3L�l4���N'���K��w;��z��q����J�����F�dQ��W���t��z���@�\�f���q��va�*���� ���|�y��yuU��C�I�6�������@��Z��M�mX8Ԁ�x�Ȉ�h/uzWj�>�Jhm��>疸F9&&���=��h���w9��f��8��r��_sd����h{^�{Gnv׫�$:5���Ec���$GI�B��(�����]Q���g�@�n�����@��Z��M<@�TW����s*���������tUq*���|6� ���m*I�;��]�\��V������]�@��S@�n��\������B�]��m%T�f���M8s3����بr��dOP�ŠwYM���l�:�V�{�����e���Y���[x�.a�vv�мcVۙMd�oВ-9�5<�Ɓ�� ��h]�@��h�nD2Z��. ?fd��U$�/����-�?[t4���I�iD�ɠu�M��h���3>33\# H1H2�F&�O{�ۡ��f�VT��&'�E��rJ��o4��� ~���ڥI��4����z����'r����[f�ץ4�)�wu{	1<cm���
]s��N1W���v�ソ�\���F����~���/:��Cm������=�Jh�S@��C@.we���n�r_ ��sj�36i�;����e�ԕU6u={v!Giہm����z���<��@�YM��7#�NH�4^�����)��������@�֬jL6�"8����)�wYM׮��}�Hى���̟��!�� K���2&{n�v-]Mv���8F2������s�&(��8����;�����C@���uNLILb��;���׮���mz^��:���b�J��w!�;�� ��2�j��W������z�`d��d�D��'@��Jh�SC�+���4�%�-���!@�5#��=e&�����7�?~m�y��m�י��ͷID�ӻ�����O�jD��2GHv�;h㭠[R 3q����u�.`�
���G@:�g5��`.Y",N�V$a�Ǝ�6��Q��E;��V�m/c�N����pV����<q����R�{�2�϶wk+�S��۵�rG��u��y���'��?#|ɞ�t�H=��vsl{q��'^�9�� w	���^��1��q���n�h��Wi�ӗ���n��w���|�R�dy���u�tP�ۜ�&�]�����Wn�r6q���[�.��S\������jNHJ�K�����K�]���^f^Ҥ��]�m���q��_���ܖ]�Wn\>�����檤��F���_�6ٞ�'m���>�RT��T.�G���%v4�� �������?d�q�UIz�B�&���ov��6> �۾�m9�Èj�����K�"�^{����}�|�}���K�P�L�������o|�DZ�5�ې�m���0���ڥ�J�y���6����|�g�N6���i�11��y#-�g
]mD�7,]�v���N]\�̜Ǝӥv��骽H���_;O�ʕ��C�m�����������?d�m%�/�6�}�|�?��ۨ^cq���l| ?�߿^s���mX%$ ���_�D�ќ����m�{����6�{y�|�Uwm�Y��ڰ��Bܗ�Ͷwf������|��W��v��|m���z�����o�X)v2�-ܐ�m�	I���>���o����3/�~�J^{�����o��>�K�M�? ?���͏����w�9�z���3���m��9��6��}�%ج �]����&9��]��Z���ǎy��"#m��w'2S��w�|�|;2V�<�D0?�m��v�����0�m���0Ԓ������c������z�U�5L��m�y�s�����)#{�現m�z��|m���2��R�������r"ԑ��vI�m���|�y����$�iU(�*Z���9������ͽ�8�o�]���*+�܇�6��$�vo���o����Ͷe�9�ު���3~��o�f�R;�q��+D����^f_�6ߒ�Kʒ��%T�����u�߽����o2���o������41\S����(����m�{nx�.���\-�3ۍY�L�kZ�,5#�gE�n�'*��n&Bܗ޶�����m��9��6ծ�-I%�m|��*Z��F�8�r�K�m��9��mR���{�x7��}ٺ����^d�m%UWv�oLۻ�,��v�ܸ}�m����m�ɘ���*J������m���|���4\�q�Wv�r�g{T���w���m����m����9�m"$az�iFB!E�K*����+"�a5��H�� _�ߟ��o���߿��*��f?? o/2_m�J�3~������>3���dϧ����<}{x�6{��3a������Y�-uH�s�ɳ���D�.F����ܼ�ϋLH�,�&�$$����>�$�]Z�M��&c�UK��m���|m��;OP7*A��m��q��UJ������Ͷ��e��{��ﶩ$����l#�Ln5s�� ������ >�~����>�$�J���I\����x%�$��6����ٻ/���7�}�m�f>Y���UW}�n��m�OC_-X)v2�-˹/�����|��T���K����?;m���~��߳ﵛ�ۂ�����0"�0��?1��3j�"D��,A�1��xR�m ��4�\<�qc��\CF�a���t�B	�s�B��a5p�y3�%`l��<ٶ.x�����~\�|6b�@��	q�IBl��Lj�$D�+�`A# @�c�����(`B�Đ!3.����Q�X�� �1f!�$"bD"����!按ㄧ�.�F_����.��փG0�<�<<y�D�#��0 ������٤ۡ5����H�lY�!!��y���Z����p:�����(M*7��o�&����jWc0�HI�`�5�l,��sNb���	3! <}aQ�5a�a��SA<'�����9�3�K�"Be�9�<޼����0�],H_����ZB*&��=V����)!�ib��szw�p��l����3 DH��� ��0�&���@X�FAY 0�EbA@�y���y�y��I�#P���p"7�y]>�[w�:H�LI�p     	 ��   mh$  � -���  ��v��  rC��  � [xp     [@ $     )�Xc#!L+�ʵ��j6��ST�c�p9��E��ؤ��i3��H���䝶�a	�D$��e8��UCm� [@  J�U(
�|j��m[[��M]�q:g���� Vmª� �id�d��ѝZx�� �Yx�V�^�� ����V��Z��W�N�8�N��H椱�Jx�עnܻ8جl��.q��1�3uv�v5�T�`������Y�d�J�v�y�	q]�'�nn��)�<�\�=n�G�*�[��-�s�JpOB������a1������w=�n���̯>*P\���+:�ӹP�b�as�$;��΢�����ݮ���=l��lq;��K��˴lL�磉N��ײ����m�x��pz��uSŇ�x���$�7V;/�y<�Їm�_���t���N���ݞ�l�r�m�0kj�K�au�]�k	�/`\�,t	eWgX!��XYZ�����[H�z`ے�
��a&]N�jN��W4��Y�q�6�cX��ǇTb}��3��n�۷��\���=Z'Eyͮe#'\"��7l���ۯ�;N��O�iQ�a�-�k{;��{�s��8�Jã�6�Z�`�J��.,�p�{j\p6]�a���"��	�vܼ0�/%q��.n��95��ij�L�y�4�pˬ��/B2q�Ֆ�W�ݪN3���d�V����?:�r����vW6�M��L���C��v.]ˁ�k��`��m�E/������Ԃu���t��W.���`�$p=d��0�vS�`$MkM9C	�x�g�Q�u��YwL��)��
Y2k]�v�l����v�n�Q�'�9���:���j����	^��[<6	����|�P?
�Q��@�N�l�PH�z":A�*4U� >֥��ִ$H���}mI�#�Ѷ�N�p��B�F�x�I|�g�D�[UJg��ѣ ��q-$�f�ny+ٱj�����j�[.툙��8p�0��f� �6��ko8��s�-e�O6t쎜��Ӯ�*��r�욝8��
u�vR擶�nk=�c��X��<\�Ƥۃ���۳��o&v�Q�l\=7+q;$訪�Q��/���y�S��9j�L~���w�~|�� `�Ԗ�\~�}�L������sqv�v0���n�z;dH�������o���ޗ�쟿��ݞ|����d�|�o/2^�T�ԊJ�H���<}�m�y�廈nZ��q�8�o�L��ڕR�P�������m�������%�*�jI/�e��$�DPR\������d�m���0�紩%�H��I�<�gm秼������r1�"n�K�q��U/UURn����m����86�왏�z�R�$UR�7޹��{��~@ܨ�\N�>������|m���W�)Ug���z�c���6��s�}�m�����r˳V���I�Ȃ]�Ց<z�<�n��T���5�p����w{��嵬����(���I.�?~_|�B�jI.����:���^�v&_��2���/�}���2$ѯ	s@�a� �Ȱ!m$	TsF�S0(�h�ѫBYL��i ����u��ة�Y�����HXLM쑗Dn:�q��"@0!�nk�* u 3|��;�>���/_��왏��UyRU$z����V
]���mܹ��{�現m�ݼ|W����Wwݛ��ly�s���Z��Y]>�Muo��?{��?߷������u��m��˜m�$�]�o�}�m��kC�9�Q�o"J)�RIz�W�$�����K��>�$�έǩ$��lƌi$:)s/,n-QU�丘��VU�n����gq��/��{�|z�؝W��)��~m��m�6��s�}�m����RU�U_�����������F
�\T�6��s�}��J�ݾ���6�����ͤ.�&���3��p�� 9��}�J�ɻm�}�����-T��b�];��EbA@�� P �E�A!P�b�P%ߖ�����m�߷�s�����H]�q��+rܳ���J�z�II���|�m��N6��s�}�o�����ߙm��Si�ԭ�;�P$����u�m���K�ϰ���������o�L���߷ߊ�����x�Z���һ�\�B	��ɣ��;�����Y�b^]�yۥ��I�5$�u�}�I{�[�RIzݦ�*_�[ly�s���k�����r)�>�����R��IUݷ����ly�s���fs��T����y�-�Cr��˷"���y��>������7ꪻ���w���z~ �۾�lN���M�m�K�J�\���6��{�>�����S7m1 =�;�}�;9�m����,�7 �M��%�6����8�RU�]�{��w�� 3���~˶�Ew.�;^���<��&z�h�hu�.���a.}�jl�y�`�z���m�������L8�̚�U���8�����S�]ˉ��&Ԓ��svp��8v���$��Si�ԭ�;��Ґ����z�M���e4�01�Ղ�c.2�rN�I>��N�{���&�J��ݜZ��nE.�r\�Gw�����*��������?fL8侪�UiU$�����9 ��G-�ޒ��o5�j�)���vm�vy`���`�%���8�ݘ۠��]8�g<�iJ�v�mht,Y�F�pk\n�Sm���<��mۣ���N���r|�gf��GG�x�O:��5t��6��;f��i�7�p��rv�gah�ܮ�VG�V�m�%��z7v�lt��L��%�H���l���!�mP�T�]\�\Vg�v�;-�i�7�B]�8�pVGvZD�p���*�m���/p[Lvdn9^��?�o�߶� ��N�2a�J��a�{���kv�.ܒ�H�R�8�̜�T�M�ݟ���?a�wYM⫕jF%!�&��8�ɇ ���p���z�$����I)=���p���Ӏ~��v�9b��L֦����Q��G?w�?rO�������J�J�*��URU���+��(�1cq��LmI���e4��@�.zװ����,�M��4v"�K�"<`v��ӱ�v�=7�].��5?!�@R
���Jg*#��-���zp�&;y����%I�_�3ޞ8/x<�j�n�s5f[u�nI�k�U"(�Sj�!�|�>�dÀ����K����TP�����Kr)t;��Q˸p�_��|�dÇ�R�RJ��JC���Ӏ{����e�4�6�6�Šz�M ��h�L8UUO{7S��k6���NqK��w2p�J�R���?�y-��h�Y"x�ۍ��E��! v�Q��ͳ���mA�/9�.��=�RsD%!�	7#�@�n-ٓ�I|��ݜ�x;W�VJ��!�3���?�*����zx��ޜ��hb���b��1�	�1h�� gs'U$��%Z�UI�٧ �^�| �؛Md*�	vԱ�p=J��RJ���N���go1>��0���Z��0c�i)&������7S���8�̜ ��i�ܷ�P��p�٣��s	)q��鱻gV۩]d�L��_ÿ�>��R�qH��p����ش[)���.��W�`�w,dj�Իr'�?fL9����T���@�����~������_?�%K�%_ʤ3m{��.ܸSR7� o��� ��e�]�z���=��Tr!)pJ�I'�T��R/f���:�|_ ��0ܚI���`�"�#�F	 #���I$�!	,eX��"��Y�������ֿ���+"�r��Ͻ���e4��h�נ}���� ���.��`-����GX�ソ�\�5�X{A��*��*j�>d��;�U�w�{�� ?w�8_s/�IW�#��^���ͦ�
�c�]�m�p�{��ԒI�n� ��4��2aͤ��UJ��%D����[嫍�,��mܜ�����>}����$���Ӏ���;���܊]ȥ�d�|$�_�I{��p��� ~���jJ��^����g�|�p�Y6�dn@�v� ��4]nnI=�ߦ�$�7��a�H6 HVD��	B�A&}��Zֵ�j�Ă�2D���z��m�������;�];$]l��� @�yT�[n�7*[�������l����6������ݸ]c�1t���0N�5�-��u\-�6��g����/Ykzh�f�:�;*�kn�e�W+�.��䞵�+ۋcSً@v{:l�vX9��x���죦rv�#��m˖��ې˧�+Y�:0��Va��ٶ3�-�G���䧶e���Zi���v�3�ۜn�Ԫ��*>�.}p�n\)�)$~ ����4]k��Rh�ՠ{.Tr!�pn�I' ��e���*�U�H�=��' ����| ���ͤ��$]�����1� 8��������Z��h���=�֢A��7���%J�UJ�����> o��� ��r�ԩ/U*K������� {����*ݎ9w����^�@��^���G�}]�v�������Y.��ѻtX�Y)�,��ݭ��$$�E^�������r'nKv�T��UT���<pL�I���������G�}]�@=z��α�2?�rdxԎ$����7� ��B)!
JE��HհVIM$�FEķ	���T^��.V��^	����{}8{ه6�$��vg�|�p��ڍ]ڊ]�p��� ?grp�UUU7��N gsI�?~�ܸ9d�S�R�8I*_�
�=��wg� w��8ʪ������ǥ������$��{0��T���s�=_��@=z���.xb1K14�'A���WK]\�N��6���n�N��m���`)��@Q�C@;���}ט��;�j���̚p���HXӒ�]����c檥M�w6p�OƀwuS@/T�e��LD�ddqi$��~��{��Qt*ECȢk�s��0Ѧ%�.<>��0�KWWi-p�J"�aE!��H$K��d�0��L��T��Sfa��KB��eee��Q���a�xx���zB����)�
I��!,H� �6l��,&�-F1�kc2��W	p�����-ܒ�����#,Cd\� @AX����	� `�Y���o�j!�������l���(>�'��E=@�J `@�+E)�ڥIn�3�p��|?��˲7ae�[n��z�����i���8Ϲ���J����ݵ�-ȥ�\�Z�#��wuS@�u�@=z��Қ�����܁�Vk��r=�\W#�y�g���g��Nˈ�J�p��^�$��98�p��(,i�ȜS�_ߦ�z����=T�W��I��`y�����\�H�� �jI��f��Қ���@;�2sUU*����O^�#�W��I�_���4^���f�z���k�c�U���R���*�+ٞ��}�� �����O�4��RC ��	&+,��b\e�BT!��Ip�H��(J�#K����  g|��rN�{f�cq��.
I/����IRO��>���r��@�qq1�"qIErz:�3�w=��8���!0��]�i��z�&�o'�z��#i�����-��|�͜3�4s�޳@�vPk[�d����3;0檪�I�ٛ{��{��h�l�<�֍I���#Ƥp�?v�������%^UIR))��������4W�`��iAcO!�@-� ����fva�ڪ�!*��o� ̼��pQ��(�rh�l�-�M�y�{�ܓ���f�T�B�Lh��+ ��֕�W���wo��I�D�� ��h�I'a,����"@�Nk(@��umK�� *��ѵ6c�yk�H�v-��[�ɴIc�ɭ,󷞓�F��]:ql�n����'�o;9�Q"k�u�;�Ͷ�<v���7k3(��/'oY&%9S��e�Zc�9Ox���kٺ����;މt�����|�4r\�����<J��ٺ�s�wnG��ȪCM��kun���&�{�wm��=[�@��]�������랑7���z�{�������?3F
���4���� ���>�;���UK��ݜ6�]�P9W,r�o���_Ȫ��<��� w}��3;0椩y
���O=�\V���G�<��� }��ޔ�=Ϫ�ʷ���D��G%�6�%�UI]�}��=�8�}V�U���e������$����pI%䊪�Y��?�y�}| �����j�B��9?�[����]C	R���=����`z���oG-���+%d��QcR8|W-����l�U�����a�l��3׾h�]�n[�SW5w$���ټ7��5	-$�F �,�Ą �l� 86ϭ����6����~(!%Gu-�����;������ ��Ç����������>O�ǅ��r
A��$��J�J��*�?��������]� o����|6?����0Q
C@���>��RK�R��z� w}��3���m���?���5G��.���ю�\rvV�'��mFa�&c���s��򱛝��U`]\�;+�Xou�;v��"#�:�ߖ�~��x���H�A��{���g{0��y��g��|Ԫ�3MZkq!�Iɠ~�~4s�i���$��Uf��_ 3{��u����.��jZ�%Á���u��� ~�d��S@�}VƖE���R-�� ԓ�nπ�ɧ ���|�ݖ�n@�gE.e�Ū�Q�.&8��c:ۓ�0'��һ�Qs#kײ�D��3{��۷�6���IzC��b��~$�JB$ܒM�Jh�j�/��@=������ѱ��S�̘(�!�u�-�ڴ�l�/t� ����\V�����mU=��| �n���ÀRI5I$�T$���	��S7��rI�}�0�7N[�mB����̜R[��>�{��g��@�u��<q#�$��SrF���һ�կg��vN�s�]r���F,۴��;!2fdi'&�{�4.������3�svp�[mީt�Rչ.��^�|�Z�h�Sf$w�,��,i�	#�?s��h�٠^�M˭z���F�,qa)	"�j���n���N��2�~���?b�A%!�nI&�{�4ٙ������� ~�d�*��~���$��H$H$r�-�:��s��	h�[�8�{o&���F��UF��ԃK!0�+A��m��<ԫ��e����rvӚS;q�<9�8�nۈw`�{v����
�5��݇���������m��R�Sm�`,
b���&��On�����b;D�ג�I���5�ʣ�/]&�N@]�ʡS�����a�Kڢ9[f�\ʚ�e�L<���v6��	� =x ���[s��Ce����G>�
l���?�ɂ�R�����ՠ��=J��72i�:�wYqY�Z��D��/��@=���Jh]k�ٕM��m�j�ʶ䶡r��svp��<�נ_;V�ԹA��40e��w'�%䪗�!O�{���5����~�����T�}���7mm�z��;�KV�pϽ���J��R*�������@�Қ�W��'�p$�����QೋNFl6՗!kj�F�����	��4�q��ՠu�@��a��R�EU~�ǻ�����K��� �.BH��s'2�QH��E*B(U$���URUd̜8ݾ��ޔ�>��U�%!�nI&�}e8������I*�$���$UT����8����&��tlt1O�2�R��Zw� }���ڤ��$���pO=�9���1�$�@�Қ�[4�)�{�U�wZ�bbD
H�v˲��[���z���ܨ�9w1��ͫ�N�.#���Is�r�5t�[r[Pw!��ݜ?d���}V�{������1��w' ��0�I6w/5���. }���/	;��bqA�r8h���I����s��yH�H*B��
�����-�*�*��<�J�*��9���?fM8��E�8ډ<�N-�]� ��������u�������� �D�� ����yUW�W��x����;�����ߵVV����v����hK ^[�O��Y��.��t'I�B���4Z�wwlξn��;w��Q�,�7�zp��]��NU��� ?w�8w�����8~ɇ<�W�f'��#�I%Ze�7$��� >�d��&��4�V�c�S���y������$����=��8��O��ܜ�UOȱR>���Ws�}�'�O����%�ae��w' ��0�ʒ�*��I	)������� ������i�q��/:zĜ&6h����0��ƻ:�;gV��m��͛nr�Á��͞Zm�l{���]��v���h�����;q�ݨ�rp�s��UKʪ������π{=<p�{��~�}ˀ�ڄ���.�o1����%�T$������� ��fc�n���\�������l��}9��������z	ʸ�8�����' �I*�f���^��w& �J��EU!%�}M�� 9�(D�&�||}b�Bh�Ɣ@�b0!HD��^4ijBl�h0I
��m�j��R3R2����@�(ɧ{�������ŗ�p�U4�     $ �    [A     m�[@  ���	   �� � [xp     [@ $     :�<��*��jV�c[MFlM�����N˧����a���5�t#,��f"ti9n
-����h
�  �   �M����K�	�.C9{;x�� ^�!�v�d�i�
S����Ŧv�N�@Wen�M�� �F�	.�Z�
U��i}V��#`W�Uݮ��7��a��x�;[P�g�[ΏR��8�����oG@Q�í
er�WWnh��f�]�m��R��Z�<K�%ڽ�	���]���-�����`�-��� ��::�x5oc��X4���j�!�/0ݐv	�Uv�n���'
�,jn�="�vh�Lvz�	�sv��2t�HKd��<\dS����*�S� �2l�v������ݧ��G]Z:�������x���v6��u��D�nWnl�=7b��imT�G$K�#B-#�q��ei��%]��k#���:V�@U�=lW�q[NװPl���V���嫩V�#N�k����9F��b�j���S�i�p�(��CQ�j�ɩ�m�U�q��\���ک�N�1�bs��E�//g�y�I�.zN�r\q�4e��z�z1-�顶�`�1��n��'֢t�*#�#�����FEk��"�E���kqۮ�:�x��F4]��;bY�ݺ���8�i���мE�6`ծ��[�Rzۀ[�h�[� qi9�qq��.��#��:7R��-I�k���AW`��X�Tܻ!�3��H�c�u�_3t��������O�k��#x��x�Y��� F��J�:d��8�L�����=b���c��(�}��ҽ�#e�t�H�*M�8g�����ѥŁn]{4*L��Q͜-69jn�k/ZnU�=]t�k���>�{����_�_@B����> qA~U"+�8�TM*lG��=�߿w���߮�����$#�! ��/Cy�`[R6i��rPi�,�� �R���[[R��� ���B�l�3/m�ر���[��l��=�� z:<:��Gq�;[�8���.�F���P�hK�m	��-��i%�污4v6Һ�7c���M���v��t+�r�;�����ő-�}����k�m�v���j��s��Y���Y�N՝I�2C����B�{��1I��v��W`��^-���N���n��Ƴ�r]�-T�:�@��5�3w~sy���������G���h[��X���iH�A73@�u�@��0���' ���<�R^Uvo�^mll��F$��;��� �u������^�嗄���!��8��UJ��]�� ��qp�s/�}ܘpW�`�n	D���G&��빠yu�@����{�����16�����������̸�l��g��:簖��l�p�Kԕ/����Km]�(�$���=����YM �[4w]��ȵ9n�hw.I|��Ô��UH;T���!,%n �1
2�XA�lI �I 3��=A_�RKʗz����� ���|����t1O�2�9 �[4�������꫼{�_ 3���;�}��P�pM2�rh�)�yu�@=z� �[4�ռX���MHh]k�?�UKʯ=���3}��;�&<�)2���?s�K%�x�6�,Y��b�����u�vl�Gnֵ�J�oK��ɆÝ86��bX�%��w[ND�,K��{��"X�%����f�3șı2�޾R���L��[y�w�Zc.\-[�ֵ��Kı/�}�m9� �DȖ'~���iȖ%�b{���6��b2�)>�l�/�L��L�ݙ�.��[3Y�m9ı,O���6��bX�'��{�ND���"�������K���*+2��B���	 b���x�� �L�u�;��"X�%�|���ӑ,K���w��5�����jk%�M�"X�~�w���r%�bX������"X�%�}���ӑ,K �&D�߹�m9Ļ�ow����C��j~{�7���ľ���iȖ%�b_~�u��Kı>����r%�bX����m9�e&R�J�/{�=�&&0��KrHRp�֊��h���T�-=��<��E�U�뀜���rO�~)2�)2����)r%�bX�{��m9ı,Os��6��&D�,K����ӑ,K��Mw�j(\�&�p��9K�)2�)gw�6��bX�'��{�ND�,K�߻��"X�%�}���iȟ�C�U5Ľ���0�Xhɚ��5r�SiȖ%�b}����iȖ%�b_{�u��Kı/�}�m9ı,O���6��bX���n����bv\e�ܾR���L��3�����"X�%�~�kiȖ%�b}�wٴ�K��8�L���m9ı,O3ߥ��0���ja��Z�ӑ,Kľ��u��Kı>����r%�bX�g��m9ı,K�~�bX�'�����Z�d2�,��5��I��������b�[]�c�MXW��9n�o��T꿕/���4\��6F˵$�R�I��K�u��v��bX�'��{�ND�,K�߻��"X�%�}���iȖ%)2�vn�	m��B˸�K�)X�'��{�N@ G"dK������Kı/���m9ı,O��{v���oq����F�(����Ȗ%�b_{�u��Kı/�}�m9ı,O��{v��bX�'��{�W�&Re&R�b۱�'*�����ıP? 2&}���ӑ,K������9ı,O3��6��bX�������)2�)2�b�����pM�Z��Z�ӑ,K���w�iȖ%�by�w���Kı/����r%�bX�߾�bX�$�0�HI"�'I'����I#mHF(� m�t��8��ڐ �g[m�N�fh�m2� @�y��N�J����F�)�j\wmmm��n�h���r9�3u��th�m���Cc���W]m`�/=����X��óv�i8�Z8���r7�;s=�ۇ��v��y�Ǻ�N���]f�Ү�Q�C� i6��mpz�k�y�e�z��`S�m�M=�5�m�j4���7�?)�1BV�������~p~�Ks�=a��k�mڻ��qx{`t/W�pP�u��,;�S�K�&띚��5sY���%�bX�~��m9ı,K�~�bX�%�ﻭ��ȖRe&R��<r��&Re&R��-���nL�2Lֶ��bX�%��w[N@�DȖ%�����"X�%�߿o��r%�bX�}��iȖ%�b}��-��i��p�u.I�_�I��I�3g)r%�bX�{��m9Ƌ����I�R
H���U T����'m��m�u�4��H�b}�{�iȖ%�b{�{ͧ"X�%�}���ӑ,K�A�y���/�L��L��=�-�v��I��Z6��bX�'�w��r%�bX%��w[ND�,K��{��"X�%�����"X�%��{�蹄	,�\��[/&�ڶ'�j3x�1;������v������2���l��D9.�r��&Re&R}�ٴ�Kı/�}�m9ı,O��xm9ı,O>�y��Kı=�Gs�����rNR���L��O��9G!胃��Av:�Ȗ'��6��bX�'���ͧ"X�%�|���)|Re&Re,�3cQKr���nMm9ı,O���6��bX�'��{�ND�ľw��iȖ%�b_~���r%�bX�߾�aL�ѓ5u�j��ND�,K���ͧ"X�%�|�{��"X�%�}���iȖ%�b}�{�iȖ%�b}�ޓ,��ƙ�FKsY��Kı/��u��Kİ�&}����Ȗ%�bw��p�r%�bX�g��m9ı,O�P�w��e�2�75�v�k�W�Ϝ7h�2��v9�{�Q�n�bC<Hn��9���k �󌖞}U=���2X�%�����r%�bX�}���r%�bX�g��m9ı,K�{�m9�L��]ٚ�r��Ӄ.�D�r��'ı>����?�c�2%��w���r%�bX�~���iȖ%�b_~��ھ)2�)2�vnڊ[j�A��w�,K��>�siȖ%�b{�w�iȖ<>8K$����p�@�)I*��++	Kd��*@�J���~ Q8dO"\���ӑ,K����iȖ%�by�}�]K����D9$��K�)3�*��{���r%�bX�������bX�'�w�6��bX�	�=�~ͧ"X�%�͋�c�'*��$���)2�)2��ﻭ�"X�%���w�ӑ,K��>�siȖ%�by�w���Kı����,��87�iv�.�ֈ�g��y;v��������Tg]�i�c��[9��u�m9ı,O~��6��bX�'��{�ND�,K���ͧ"X�%��s6r��&Re&Ry��i�b��$�j��ND�,K���ͧ!�Pc�2%��w���r%�bX�������bX�'���6��bX�'ݝ�2˜�i�td�5�ND�,K���ͧ"X�%�}���iȖ%�b{��iȖ%�by�w���Kı<�~��5p��pp���K�)2�)>�l�/�N%�b{�}۴�Kı<ϻ��r%�`t�DP��m6.�N�|�m>)2�)2�l�h�wpjZeڈ�NQȖ%�b{�}۴�Kı<ϻ��r%�bX�g��m9ı,K��w[W�&Re&R��姢��v��dr]��;t�Yjz��c�H1���p'�l��]�hdѬ��5	�SYs5v��bX�'��{�ND�,K���ͧ"X�%�}���a�Eg�2%�b}���6��bX�{�����$5��U?=ߛ�oq��'��{�NC���,K�{�[ND�,K���ٴ�Kı<ϻ��r'��J�L�����R�!�%��/�LKĿw����Kı=����r%�bX�ϻ�m9ı,O���6��e&Re,�3cQKrJHF䜥�I�X�'��ݻND�,K��{��"X�%��{��ӑ,Kľ��u��K�L��3n�V��ImFI)|RbX�%���[ND�,K���ͧ"X�%�}���iȖ%�b{�����K=�{��}����K��"D�ڐH�m�����Gm�Ҫ�"�j��>�l9�-�H͓���� ��!f��l�Z!xah���[�=�ˡV�F҆S�ъ�.�gGv뚒��g
��Ŵ�=���`ҫ:{�d�Շ6��P:��Ɨ�:���ßb��e^���J=�$��ۍJe�t�[1��7�v�S�z_YeEt^í픓;_{�������yk㗎`�������t9ۆ���UfM���{�\�h;\Gi]��j�rdі�ּObX�%��{��ӑ,Kľ��u��Kı=���r%�bX�ϻ�m9ı,Osߥ���Ye�8Z��|��I��I��_so���"dK���ٴ�Kı/�w����bX�'��{�ND�,K����\��5-2�K��_�I��K�����Kı/���m9ı,O���6��bX�'���ͧ"X�%���^�C���OJ��������v���g�w����bX�'s�߳iȖ%�by����r%�bX��~�m9ı,O�����$5���_=ߛ�oq����{��ӑ,K��=����Kı=����r%�bX��~�bX�<~����n�h�M��S��]nDׁƷ=�u�N�����at�ɉr�k?q"s6o2^Hk!�j��ֳY��%�bX�����ND�,K���ͧ"X�%�|���a�șı;�~��ND�,K�5�ڦ�eִ��S5���r%�bX��~�m9
�A �W��iț�b_��5��Kı>ϻ��r%�bX�g�w6���*��S"X����kF�ѓ5�M]]k6��bX�%����ӑ,K���w�iȖ%�by����r%�bX���w6��bX�'��2[��nL�2ۚ�ӑ,K?��T*�`j'߹��v��bX�'���ٴ�Kı=���m9ı,K�w[ND�L��Y}���Z��pp����&%�by����r%�bX����6��bX�%�߻��"X�%���nӑ,��L��ݴ�Am�.DH�5.4З%�:n��s��p��nzݩYy��/p_��{�ߞ�19�RsY��SXY�k%ֳ��Kı>���6��bX�%�߻��"X�%���nӑ,K��=����K��K�����ڻQ��.��/�L�bX��~�bX�'�뽻ND�,K����ӑ,K���}۴�O�{ۻ{����q��������D��6kZ�r%�bX���߮ӑ,K��=����K/<� � `����N�\�ƎP��8b�F��*��0�S@�X�k!
����a��d�$�B�s�Ysi(�`�е$�!$��0�P����h@�"��BM��
B�Y� �0$FKS����ѣ����@�FI[Y9�L���f�%̖�<R���K�F�(\ &f���������, �ޚiH$3F�.�+$�`�X��2�*��K���`F$�f���#GAb[�1!\00"T�$��`�Q W��J� �	(A�Fhn ��|�1����l�*�(����F(�}�1��JpW� *��Q6�P ?
��z>�=�bw�s�iȖ%�b^�6r��&Re&R�b۱�)b�49f�WiȖ%�by����r%�bX����v��bX�%�߻��"X��$�E�����)|Re&Re-�7Ѩ�q�J�S5���r%�bX����v��bX�%�߻��"X�%���nӑ,FRe/����/�L��L���BD�cۣjM]���eӜ���7pN�N�(,�����R�sѺ�4��w��,K����ӑ,K���w�iȖ%�by����~Y�L�bX�}���N�I��Ku{ȱ�����q]�rr�"X�%���nӐ�T�L�b{�w�m9ı,O��]�"X�%�w6r��&Re&R���]��j84�u���Kı<�~�m9ı,Os߻�ND�,K����ӑ,K��u��&Re&R��6]�R�.��u��r%�bX��w6��bX�%�߻��"X�%���nӑ,K�1DW2'���ͧ"X�%����h���4MMa�e�fӑ,Kľ{�u��Kı<�]��r%�bX�g�w6��bX�%�߻��"X�%��{~��<9YT{>�7a� 
�����nֱ�s�q�t'I�B�j�$5l:ֶ��bX�'�뽻ND�,K����ӑ,Kľ��u��Kı/���R���L��]�[v=,RF�,����Kı<�~�m9ı,K�w[ND�,K����ӑ,K���n�R���L��Y�fƢdR4:��y��r%�bX��~�bX�%�߻��"X��DȞ��߮ӑ,K��y��R���L��Os6H�F(��-5��k[ND�,��������r%�bX���߮ӑ,K��=����Kı/���m9ı,O�;�d�9tY2�2�ֶ��bX�'�뽻ND�,K����_w�m<�bX�%����ӑ,Kľ{�u��Kı6P�"U"YQa�`HQ�����߿��L�Ҫ����궺 [�P�流m[@�3�l�݌=W=[llҽ8ӭ�+�'��iД0�(�5��3�k�͍�u�}-Nx:��=���ݶϭ<��m��m�%� �}a\v���LN����mٸ��i����B-ཉ��	lͮ�[=plcg���g�v��<�SoU��s�g��Ҵ5=vE���#vu�'�ƶ�F�Q�g�-~�����w�{���⟙��/:zĜ&6��{a�p�b��.��[d��O�����[F�s���iuu��r%�bX��~�m9ı,K�w[ND�,K������<��,Kߵ���r%�bX�gݤ����)�,�5��Y��Kı/���m9ʑșľ����r%�bX���߮ӑ,K��=����ı=�_wV��SXj��Z�r%�bX��~�bX�'�뽻ND�,K����ӑ,Kľ���iȖ%�by���'R�$�_=ߛ�oq����{v��bX�'���ͧ"X�%�}���ӑ,Kľ{�u��Kı<�KnǠ��H����/�L��L����siȖ%�b_{�u��Kı/���m9ı,O��{v��bX�'�����یcl���
\^+�[s��[��؝tvX۬�3�r��-T�:��qz_6k6��bX�%��w[ND�,K����ӑ,K���w�a�D'�2%�e.�o���)2�)2��金�b��֭5��k[ND�,K����Ӑ�� F"$ ��R1�1�MD�;�~��r%�bX�����ND�,FR}���_�I��K1n����љnk[ND�,K�u�ݧ"X�%��{�siȖ?�"_�w����b�I��s}9K�)2�)v�Y.�je�ե�֮ӑ,K��=����Kı/����r%�bX��~�bX�'�뽻ND�,K���N�35
k,3e���r%�bX����m9ı,? $s߻�[O"X�%�ߵ���r%�bX�{��v��bX�'��s�R�!U�Ÿ��[�5�6�R�{A��kV�ۯ\�v������e7/]=��ӑ,Kľ}�u��Kı>�]��r%�bX�}��v�y"X�Ry���/�L��L�ݞ�p�m�r�r�r��&Re&R����_�I�by����r%�bX����m9Ĳ�)<�l�/�L��L��"۱�)b�T�Y5��ND�,K���ݧ"X�%�}���ӑ,~Uh8j&D��}�ӑ,K���w�iȖ%�b{�_v5�K�ԅ�q��&Re&R}����Kı/���m9ı,O��w6��bX�'��ݻND�,K��wZ��b�ˑ�%ܓ��)2�)2���ͧ"X�%��w��ӑ,K����iȖ%�b_��u��Kı?"g�����R�vW7'��Y�V�tN���$���'NU�_۬���0������w/_;s��ۙ�333Z�{ı,O����6��bX�'��ݻND�,K�߻��"X�)��w6r��&Re&R���]��l֭,�k6��bX�'��ݻND�,K�߻��"X�%�~���iȖ%�b}�����P�,K��>�L�)���5��WiȖ%�b_��u��Kı/���m9ı,O��w6��bX�'��ݻND�,K�~��̰�$l�G$���)2�?�R���=��_D�,K�����r%�bX��_v�9İ ���T�����)}��Ӕ�)2�)2��{c��mK�z�WY5�kiȖ%�b}߻ͧ"X�%��_v�9ı,K�~�bX�%��bX�'}���!ae�6*�\��Q�\fd	�ۯLn�Q|�Q�6�(;G�eŷN�ă|�~oq����ߵ�nӑ,KĿw��iȖ%�b^���a�	�L�bX�����r%��L��SލD��u!n\|��I��K�߻��"6%�b^���iȖ%�b}߻ͧ"X�%�ߵ�nӑ ��"w�w0�X[�i��i7�I�{���*AK�ܔ�$��*)x�����Kı/w����bX�'�-;��`��	.䜥�I���e,�߶��bX�'~�}�ND�,K�߻��"X�%�{�{��"X�%��}���j�E�Fӹ')|Re&Re-��ND�,K�߻��"X�%�{�{��"X�%��~�6��bX�'�p��I%d	X�T�6�)@e$�H�4%#%�d�h���N�Zֵ�[x�Y�H�6�ïCsZ���v5��l��d��D9�*^Ws!�hGP��-��i8��t�5[�%�:�A��mѬ�=��Uz��:��[Y`�����I2�cn�tuˬ��{6q���٤#r�h998Z�pPl=q<-�v��y�Aƽ��ܶɜ3v��si;��1<�m�cä[s��4]��j玶�c��s��"\V��V�V�-R�@7�A�؆{\����f��rf]ч�r'l�rT�d�kW&j�Xfˬ��<�bX�%�w[ND�,K���[ND�,K���ͧ"X�%����iȖ%�b}�ߧ�e7/Ph覾{�7���{��?���m9ı,O��w6��bX�'���ݧ"X�%�~���ӑ,K����ش��-�N������{��7��w��ӑ,K���}۴�K���/w����bX�%����ӑ,K��d��,RF�.]��/�L��$�������Kı/w����bX�%�߻��"X�%��w��ӑ,��L�ީ���%ի$\|��I�bX����m9ı,K�w[ND�,K���ͧ"X�%����iȖ{��7�������e��Ğ��De�ǝ�ڻ�=//�����-��M�ӛ�6^ӯ�v�왭ZkY�ֶ��bX�%�߻��"X�%��w��ӑ,K���}۰�<��,K��kiȖ%�b~�~?\�i0�\��w')|Re&Re,�;R�P<D<@x!�l�Ȗ&��ݻND�,K�ﻭ�"X�%�|���i�I��I��y�����[$m2�R�Kı<�_v�9ı,K���bX�%�߻��"X�%����nӑ,K��;�5�Zi���55sWiȖ%�b_~���r%�bX�g�w6��bX�'�k��ND�,K�u�nӒ�)2�)w3_їlWp�#Q˹9K�%�by���r%�bX�{���9ı,O=�ݻND�,K����Ӆ&Re&R��6'v�cZ�K�a��11�^m���v�p�k�0�{7n]�\���"�Ӗ��fh��5���r%�bX�{���9ı,O=�ݻND�,K������<��,Kߵ��iȖ%�bw�~����$`�#�/�L��L���5�D�,K����ӑ,K���}۴�Kı<�]��r'�@ʙ����Q9$��d�K���)2�)2�����ӑ,K���}۴�KP<���!JB��:4�`I#�
�HF+E�A(��q5_k��ND�,K�u�nӑ,FRe'��$V�V\��-�9K�(�,O=�ݻND�,K�u�ݧ"X�%����iȖ%�b_O��bX�'zt��f�&C5��u��ND�,K���ͧ"X�%����iȖ%�b_O{�m9ı,O=�ݻND7���{��o��-�a�l�#AW�ږ��%�t�mcLg�ۻY�����4�L&Y�ZIsY��Kı<�_v�9ı,K��{��"X�%����iȖ%�b{�����Kı<n�֚k,3M\��r%�bX����[NC��"dKߵ��iȖ%�b}�~��ND�,K�u�nӑ?*�TȦR�o��Wl�E[Q�w')|Re'���w��r%�bX���m9ı,O=�ݻND�,K�{��iȖ!���o��iC�[���>{�7��,K���ͧ"X�%����iȖ%�b_O{�m9İ8��G7���|��I��I��f�e�)b�0r��k6��bX�'���ݧ"X�%�}=�u��Kı<�_v�9ı,N�wo��)2�)2��˶��w.˒F�ݻK�ݮ��ˋt���.�GJԎW���w;��/&�	#/����Y��b_N��m9ı,O=�ݻND�,K���ͧ"X�%����iȖ%�e'��$V�V\��-9')|Re'���}۴�Kı=�{��r%�bX�{��v��bX�%����ӑ,K��N���3E�!��5n�WiȖ%�b}�����Kı<�_v�9ı,K�߻��"X�%����iȖRe&R���Z�al�����&%�by���r%�bX�ӿw[ND�,K�u�nӑ,K��=�siȔ��L��b�n7%4�vZ�r>R���X�%����ӑ,K���}۴�Kı>�{��r%�bX�{��v��bX�&��j: 0b�a�Tfg�0� ��R��&ijα� �[%6�BT��))�a3N�f��Y�;�)a�\�"��H�Djċ5kM�r0B�ތ֋����봗	R1%ҚH@2����y��g1d�T�hI5����HK��aFP����!	$��Z!	�Y,��[a���D�[
���F!0�2с	K�� z�TH�� >B$��x�w�5��L��K�m�L     @ $    h��@    �`��l  ����� �  m     � 	     gI-1��i�����[i.�]J����ʚ���l�m	��R�'FR�ج�j&���ԷtE� m�    6�`-�6�qՒQ�i�5ܧ�dˡ٩yb�im��9�v���U�A�ŴP�ێX��6t��'XiA�Ŵ6غr-R�g�nn���BuJ��҇i��s4����m-˶�c�Q�j�،<�0�K���0n[r���;9�V�)�]��>"v�Lbx�7	�碣 p��]����#��nݹ89dqv}����Ō�u�b6�q�{8���#��޸&�%._(�m�َr��c�@
�x��{l/��^:��]��t�OH��<{@��,��㦬v�=m���l��F۴��o��V��t4B�u�2��c[\�,�Vp �������㲮��D4X�����W�M��cLjM#��Y�2+��R�,��U��#)���:�IK�*m�݀6�a�8�Xm����6/����m�+h��[�[5KӐ�jL:��{a�8wko��6z&��j|u�t�Z�N:�[�8�ジݓ\:u�t�
�����7!c���i�L�,��y,v=[&}m�q��hyj�{�p�9��y���n}a!ݹ+q��m���N��<��9�]Q�7�l�d��4���vE�'�3Y��[�25j��C��e�6�q��BUV�s�`C��u���5g��{t�^㝷������$���/
�6�J�u'nP˺��%��]�s�V]�sq�jg[%�K���t�3�p�--��jvu�����ksƶ���H�&��ܦ,\�nzu���6�'��Q뗀�cq+YK�$�V]{4�R0��mWKj������:F�5i�WuGj�te�j�K�(� Z*�(?���.���\�E��{�^���~��O�$H-�9mv����:�� l��q n��K����i @��q5/Qn�s�U[z\i����\I�ݎ.ͷ���>��U�����yXͥ�pu���[��NN�I�{c������.���ŋ��)�,��ptulx��q4�˦�It�u������l�����K
����`�m�]t���˷`�;K�u]+h��Y����y�y���r =�tSD1ۋ7KS�n�t����Q<sɎ�<{'Nj�LZ�3��L�����S�%�b{�}۴�Kı>�{��r%�bX�}��6��bYI��V��R���L��[�68K�Թ��jhֵ���Kı>�{��r%�bX�}��6��bX�%����ӑ,K���nӑ?eL�b{��nL�!����$��_�I��Kwy㔾)1,K�w��iȖ%�by�w�iȖ%�b}�����Kı<��{�h�֫�2k%�Z�ND�,K�{��iȖ%�by�w�iȖ%�b{�����FRe&R��i�_�I��I�n���&kV���kiȖ%�by�w�iȖ%�b}�����Kı>���m9ı,K�߻��"X�%�������ǘ7r�'K[��s�ڻx3��4�N^����k����؂ݥ燞�����*�O"X�%������r%�bX�}��6��bX�%�ӽ����"dK�識�K�)2�)e��d�v��#d�5�ND�,K��fӐڜ�,��,(A�}A:���8�q�O"X��<涜�bX�'�k�ݧ"X�%��{�siȖ%��K�kq�)��Է.��I���%�ӽ�ӑ,K���nӑ,K��=����Kı>���m9ĥ&R��i��mq\���I�X�'��{v��bX�'���ͧ"X�%���o�iȖ%��RdL����m?7���{������ZP��k���9ı,Os߻�ND�,K��fӑ,Kľzw��r%�bX�g{�߻�{��7��������]2��M��S��kr&�	񃮢wq;����9�Să��$M9rI|��I��I��3�r��X�%�|��u��Kı<�����Kı=�~�m9ı,O=5��.�����m֦ӑ,Kľzw��r%�bX�g{��r%�bX��w6��bX�'�}�ͧ"X�%�~��ִa�9�զja�kiȖ%�by��siȖ%�b{����r%��2��AFm�"j'{���ND�,S)<���)|Re&Re,��ݧ󉅆kP��kY��K��������r%�bX��w�m9ı,K�{��"X��P��~��6��bX�'ٞ����d��w/��)2�)2�fsNR���L��O�V��|�����}���z׊�DJ`�Ƣ��8�!t��k�u\۝���	��+��9���� �I1�j8h��f����^��Қ�U���L��
c�@�[o��I&ξ�� �ɧ >��' ̾�p�������@��W�wt���$���vp�7o�|����r!;���`f���=�����	(V���Q�ߺ�7$��>�T�u�WXd�� }�fN��K��m�r�_ ��S@�������B��LblMι�c�=�ֽgͱ�����ЋZ��ر�j���1�D�A�@�wW�{�U�}�)�v[4�q'�T��!�H��=Ϫ�>���-�˺���J��������t��}�l�>]����h]�D��X�n#Q�@=����ަmoK�(��������ǋSY&Aa1ɠ|���=ϱ��ه :�2pUT*��0v�rHH� � ��h���'��`$-�bE�חi�nz!��ڪ��:*RU�-�lˍ��̼Ԏ�8���n��������Ӷ�1�zv��PR{:����ۊ�Yn{a��'�Sr��v�Ҥ'`�p�LWm����HE�:�b�n��,B��]�\���K�O7a��uV��=vmty�T�9�Y;[�C�t���ѻ�����y��R��9YT{>�7#� �tǑ�kc�;BNݵ�v�t'I�B�j-(Y��k��������@��S@;-�@�wW�yz��C�ra�5$Z�Қ�m�˻/�u�2��UI6w�ƢrGRՒ���`���`zwz�;�Ln���&<�Ɍr%�<�M�ֽ�Z�wJh��4�q'�T��2I#�9u�@�t��{-�@�u���~�x��AK��@c�X��Ɔ�7w8[��\=�<gV��qk�oK�`�vC(q	Ǡ{�S@=�٠|�נr�^���H�O�x�H��m��!=���8%-(&��ƺF2�	rYt��F`J����m*��e�D$�JIS���2&���aX@�HĻ�^?"�y{ϳrO/}�ny�Z�U���L�ib��$�>yܾ���᪩Ro;y��[�8쳬L��'�&7#�9u�@�>�@=�٠|�W�yz�����ra�9$zy�Z���z��Z����?l���8(3s��%�9�պ;9j.���+"��zCL�wqQ��Fqh��4��z.������&<�Ɍr%�<rM��^��ֽ�}V�{:٠[n$�j���Z������3+zYHP��$���W$0@0+� b���}�m�.��.�V�`�e;�p5U%O�����6p����^�@�}R"�jD���he�4��z׬�=��h.��#f
�����dz5�����k*h�C�#V���뷐��p�0'<But8��_6ߏ�e��ܜ���=T�W�[�8v��&(�'�&9#��f�~�����_� \�M�ܠ_roFc�H��@����Қ�ֽ ��hy�LNC�cd`G��_U�zs������	Bi$���%
�U���1�FLc�,��h/Z���N��� ���>�J�����nOGX�'S۷h�M�3Z�N�h�'�^�|�2����ޔ+��.vs��-?�ߟ~[2�����zX��N�<�LCC��NI�^�M���@�ֽ ��h��DNG�)�"M�@쯪�*��@:����;�V<Z��2	��L�ŠU�^�u�4�)�vW�h�jb�P�'�&9#��f�{�4����Z�'���� ��q�8[���ְ-�h
m3�ى4=�X*�u  Pt�hMm�]�֎1նMN:J�7B�{m�<ʝk��&�C�'Q�ҮD��_0�i���9���d:��m���ڶ��<t�z�Pi7cQ�����B��3�m�	�۹�Dz�ʈ�A�x�>䛦�6�����n-N���=�_
��m�,9��{�ѷV���&
���yR�j�4�fqdnܻ�=��V�f	m҃�yKŷN���͏��Ɓ�]�@�ֽ �l�>�,����ǌ�iHh�ڴ
�k����Jh�d��##1ȖE�8�
�k����Jh�ڴ�jc2d"nG�m���;+�hzנ|��[��Hhq��4�)�vWj�*�^�u�h�?~�n@7�A�؆{\����JCcu��W ��8[`�;�����`��@��M�@�ՠ�� �l�/t�������I�M,Rdr- �����"�(FH{(BEcB%!D� �F@��"��)%�"#01���]]��!6c7u��
�jYrN f����4��ZoY�rⷊ�)���&��-�M��V�[�h[f��;bɉ�Lx�Ɣ���]�@�I$�sg����fva�5R_���?:YYcp���Z�[�yݹ��c�Gɻp��G:1K��;b�����,�mMyz�_ ~�������)�vWj�;��O5���d$qɠm��S@���| �̜�T�M��`��;l�\e;�pݚp����.~K�RH(Q��4�Q�=Ip�s�b����H�H�%e20�G� @�cp�����,�B	��պk�I�)-+]x@4B�d ��)�AFM��h�HSk	VsD������ @��Yu�30��]��h�ˢ`Ma��0H�|�ټ&�D��P�� ���<�x���D����D��8� ����<P>ClO<OD�E}PB�1"h]�iH.y<�|���=�[�{]�9�'�)�"M�@�ՠ�4��@��h�-Md���L�E��4��@��h�ڴ�Y��?���	$��4Lbcv����ӹu�{:��<���[;�m='�"�nM �l�-��ev� �٠r��C�r`�rh�M��V�[l�����&'?���iHh�ڴ�f�u�h�M ���1�FLmDcX��@-�h[f�m�����FWj�;��OZQXYd��r��s2pUU����.~�- �٠w;Q��F	̎	A�'Ϗ�nm�eY3�ǩ:�Oh�&���{Z����n&!��'$�߿OƁ�]�@-�4��@���D�D��bȕ�8V_q�ʕ*l7sg 3sg �즁�����I�b�#qh�f�u�4zS@�)�r-ʘ�2	�Q�I�z�ޔ�;/Jh�f���7��)���&��-�F���wo[ �޶D(p��!x�  ��R)  ���HQ��� �-��T��U$
�~��rI$�� I���nӦ��6�Ԃ�����s:�k�͠��Z@��au�BF1$�!R����l�÷b{%pH�3���V��T\�4�r�g��s�������My���ڰқ���4�#��p{tp-Φ�:�zlv�r�#k�g��u�ۤ{��ўA4oog�`�+L��eF竮�];��>m�n���\�J�+���fqT���5�f[y�3Y�ZֵIBr/*K�v�N�N-�n�ru�v��ą����/r���LNAL�qP>���wY�r�^��>�@;���Ǒ1��b��u�+��s��Қ\�z�)�b#26�+��y�Ze�M ��f���%[�4�I�!���������}�@�z���H�D�xE1diH��Қ�?�͟�so�}����}��Om���V� �ś����f|hޭ��sŬ�n�5w�9�����t6��ߟ����:�|���z�UK��&��Z�r�
��wd�p��_,��$�X�� �@$R&��֧�}��>Y� }��9�U��5�ڿ)����Ǡu��@�)�{��9^�@��زbs�
`��#�C���B�_s�`���6{z��ޖ�ِ.�Wn1[NHp����=K/s_�{����Қ�]cx��HĢ�{N�K[���a��^�r�����ֻ\��k��k'�8�& DfF�@�z����_�a䪫��͜��ƭ�۸�\��>��5RTً�4��͜����RIz����RR�����r7�DԶ�|�����ܜ"II(Q	8�M��z��ޖ����SY&m�&CC�fffb^���9�m��}��ڪ��wy� �wV��C�'�69&��z��}V���)�w�8�T�=��h���v�ڶ(�v�������8'�E��z��;r���9�S���{ޤ"�9�˴��\�d%ܾ���>՝�p��'���6����N�A��,D��VvaͥT�ٛ8_��}Ϫ�;���pK'�j#��8�{��~yܾ�%�H)*�wݽ������Ř��+p,�).I8OoS�[��՝�0�*!j"A		XFH�� /��=:��T�qc�m���z������h��hW����Ƃ��$b�1��c{^+���&��&1��s)���;��ww����o��4�O1qѥ"����ۚ�u������Z{�ǋSY dm�&�����<�W�}Ϫ�;=n���ʘ�?��6���<�W�{�U�vz�� ��N |gm<w."�K�|�Kʄ�^o7πj����w2p?�RI��m����bs�
Q�G��z�h�l�9^�@�>�@������$�$H�[R	����v�imD�4Y��%UK{F�%l��Ԁ�\�]N�R�B����yiL�"Ϊ���S��ɛ�ꇄ���xZf�X��X��,��S����y�ۊ�f������v����X�4�a�n�9���2i"���Wj�;�f�պ�Ŕ��/\�:�,��\�vyĥ�WR9�E^�y�#h�Ym�zut8��tY��n^�wo{�ikW1��Rj�]�.���=��^�s`�f7a��zUkg�^.ň�ۊ�lyHܜM�ͱ���ם���}�����I/��������ؔ�"LMdn94W��=Ϫ�;/]� �����n,x��B�@�>�@�w4�h�W�w��"9�$SF��@�w4��Nם��o���7���77�Z|Md��RdNf�}�����s���s@���"x�ۍ������ ���=�B]�}��=�S�z�n����=�S�=&(��<���4W��=Ϫ�;3����I|�������OA]���Mfk7$���뿈⫰D�S��8E�}���zp��_ ���'r��+r�K��ugs��w2p�IU6f�������Ζc���҈ƱG3@>�f�u�4s���s@.wen8a$M�n94�Y�{�U�v[w4�Z��^*8�M���6���'	���xR��8.������$��y
sm�z4qc�m��19&��}V��m��>]k��mp���G"Q�c�ґh�� ����f��}V���cf���|v�H]��
]��:�޾ w3�nh>I A��aXB$�!"AC�����˹'��f�����1C��6����ݾ��Y����T�T�^n� :n�z��ʸ�H����}��?�Ż�/���= �l�-����! ĤHs�
]!��.ۚ:���dj�d��n3VT�tHC���'?�D�(�#�@��h.��[f��}V��Ζ����bR.��e�ԛ���;���Vfqp�vT��7�H�������J���I������1����ϧ[˸�m���4s��n���sr�H� F0�QIbZ�T�{��gvm�K��jG�ґh����ֽ �l�=Ϫ�������w
��]q�2=�ݦ�y��y#�n�x�m����t���R� �273@�u�@:�4s��ff���a��� �g��r�h�Ww/�m���Ze�s@�wW�-x�S ��7&�}�f��m��>]��[f���\ND��(NMRKԒ�^��.׻��s2p?�R��o�^�?@p�ƔF5�I�˷��ow[ ��[Ww4��<�D4��8.�a�k��$��6�m�I�KH�i#�)M!C	&�����0$H�٤��pR�IĀFB
�I�����9) &�CH	��-��b�	A"@9(�������p��	J1�Ja1���	rf��3���5KCa�@��c�a�HM�c3�kd�$&�4\$�D��!�X�:6��*�0(����$��I@���,y:��
�e�;w��     8 	    �$�   m��� m �-��� ��!� � [D�    �  ��   �E����kn�e[�@:):�"_���+���NwQ����7UƘ����m�ua�RėrA��}�"� 6� �  &�6��-�n��کG��rV' �JR��k6r�v��5��[�ek�`��-ƣ,D�\苲�v+���6j�+J��U��ө�H4qr�*�4��������4��(r�]۝&�<ܖw�k�X:AW��3s !��#�sE��<dN�M��k��P�5��ݲVʟ���7�`=\��>�W\�<��P��nQ�\�1�rU��v�n��M�5���9S�(��� �`)�n�tح�Y���P��;]�y��j��R��3����+f��[�6rq���p0�+��h��p�c��F7M;��x��O2�R��!yԅ��@�G8qGa�8�y�n��mHNӺ �͓n��<��'3��@�ڶ�j�kU�A����vW�ȵV�# �����7�ڪ�$,(�l
kf�����6�%��m�ۮ�Pz�ۑt�v�r3̋���&]�ֻ m�qٵ�����e�9���.�T岑��曟g%@�[V9۪�����2��e��oN)J�B�Bm����۟i3i�X<�Q�b@9tm��+�����:+u����4�mE&��PZ�T����Y���8�{wD/��uR�G�d����-���upl���n�3��]��7+��+����V\��-�L��%�l����J�l�|���+�̉��jz֓aM<��2�b�W=n����r�gvy�J`� �@R�:���ݹ�l	��l1�[t�1��䁠��$#����A׭՞Ͼ�۾�7n��5�Ў �j �"�Pt��0A>zz!8 �A<E}A ���2��Zֵ&�I�D�G-�ޒ�B�}��` @UT!��@a���TW[llҬ�jt��v.��h�����:��.�=q�-�q�v�'a]X'`������wv�m�gsp�t�`��z�f^���㎷;t��T�����A	�d��U�������5Ϝ�I���; ��cxLW]�E�qS��d:n6:�!"�N�$붃Cd����3F�&��z�3|/&j�WV�D�.OGX�;�ݻt	�݂u7m�A��|��$Xz�����fݗ������o߿�����h�����@�㒭��.���'rN }�����R�5{}��:����^�@��Dy"��cRM����>]��^�@>�@�uLZڄ�hN��|����f�}���y%�W���ˀk3�v9c�B���z׬����;/]���^�}��B<IR7 �7��=qə�Is���s�i�2��A��/nn�0���4��4��s@�wW�z��y�������)&��z�o)RI�����?w' >�rs�UT�%�IT��z@�K��یVӗ ��_ :�����e빠-¸��x��I#��f�}�f���w4?�US��6�<1�w ���X��8����i�������u03+��܀n+��؆{\���jk� m[�ٞ�ݎA��wGS��w|�����4�=u]��[�4����`zs��������[P��M	��h]��/f_ >�d����=I*M��;�v���d�6Z���N��0ou������B���m"M�L�'�ZƂ��jD�tJ0 /�!(ٕ�Ƙ=�Lr{���+�d�!w/���vp���pϽ��/Z���e���X�&�BI4g��h]��/Z��hZ�Kr7��z:����y:v{J�ɶ�htu������z�孛C�R7'Kwͷ��r���e���OUR�U/��}��/y����˖(����e��ٓ@�{����@�|�NE $cr�*�����y�NoSӝ���5H�<��@�{����߳rN_>�7'A҂DY�C�R�T�%�[K��ٽ����|�p���MX��L�ަ�;��{;���7����wy�;�Sm���R�-I�v;C,�W$,����wLݝr�b�q�gx��e�qISe����;���=���ś�0<���yZ��&AL!2'�}��`b��9�LNwS���2d��?s�,�&@��h�nh^���fU7��v�����~��d��M]��r���'7�����`��`b���p�(`�!�dRH���z�w[o4����`8Imf�������Ąq�$�����ְ-� �V��k/gm�#�YP� @�yT���l��h]mգI��:�?���;r���y�^���m�Iېa�Ol���mV��\�Dn� a��`�����ݧ�gv��Ū�t�˺c9;)�̚�t]�+��[��t���b�6�N��{�ų��6�]�81sr�M���r爸�j��L�e��{��cy�p7U�v�R��_�ݛA�i@;I��>�����2;vݭE�9��s��܎!Yw,R�������� ��w/�UJ�������m�J(��ELrI�{=�sf$r������z٠{֦-mBA��8"��';��{;��fw[o4���
���CP�iǡ��K�����vp��s���I$�}ݾ g^��t��E�d�� �������=����l�մ���l�H�Y�1yu=�v+N����A��J�gj۠��ϧ�^�52�s�,�&@��h�u��<�k��l�z٠{�e��Ōp1���ܓ���f��@��z#�����{��}��1f�L�r:�lER���swWL��l3���	DJ���s@�߿=��UI	�1�̕wl3���y�NwSș���`^���X����"y1I&���]����%��}^ ���`����uҞT��n�KNܺ݋,�!��f|[Yӆ�&��in�5w�9#1t��6�7|�';��{;��fw[o4�̤OuTa!�D4���l�z٠{=���??ٗ�*T�g^��-A�BBj�n���1f�L�B�^I�	)		x��5�\��ܒ{�k@���9��F� BI4g��h^��޶h^���Y`8F�c.���\���|Ԓ��wv|_wo@�{��zװ�����&��1٠q�b�c�N��sڄ��{A��An����|��p�0o�2) {�~���z����䪕|ï���3/�$"#i�drM�ֽ���z���z�bQLq�q���=���z�����z�jƵ(���"\\�T���ɞ����NI<�}�n@�|P2�߶nI�K�x�1c�G�}�f����s��w��|ʩ*{��2�e�����}n����û^��[��9�C�l�79Om�4��s� ��NO���-��w4s�޶h.TW��Y��G�?/ٜ\�U&��� w���}�ՠ{�e��Ōp1����=Ϫ�z٠}�ՠ{=n�\낰��fAI�{���v���w4^���䪒$m��@�V��1gsL�ަ��l'�����䟠$H,�$r�6�'amu�j@�εT{7�.�ڗ;0K�n�=)M�k�H��A+$E��!'[�p��Cn	�ix4%m��zv8t+`[����ۚ���;��Ϝ�Iu�������>��/d���N��Ggs:����o�Ɲ�<bh�{nƸ�Z�9��G���l5���w�6��n=\�C���sc����t���=������w{������Ǐ池�5��ř8�J+oF�>ٽ�f� c�2���a��lRpS��O$jE@������r�W���@���@��X֡�1A0N)3@������&ýݜ��k����.j�J������0�bI��z����>���=��s@��@;���dy0���8I'�fk�]������z٠}�S�AO�?�9�����/uz��hW�h���I��6ъM^˰��1Y��W�s�1�1;����V#���b=v�m�ix�7����m�uP��M��@7;�s@/\�f75a��kY�$��~��@��Ҋ�	E���`b��9�L�ٞ���a#m��94���۹��3?������@�H�I�<�9R����>�� ;���e� �ڱ�C�"$�8`����������{󿖁�[w4�s�Hى�@��7#� ��t'��]�<�Q�v��۰�N7A�p�1s6�p͒��m���~�����[��r�W����dy0��94���n���^�^�4��x�
)��	ȴ���7$���ٹ��$��hn�����C$�L&d�3LB*A,�ap��q��BҤH�	5*K��P�i	a��k.$��BF)H�(�*	@���-B�d9(�"B���	��A� �.�X�D!`�#	� �"�r�f�:�g�s7�ByC,4�0�h���!Ad)�ZP�Bff74RX�!��H_!��c��������laC��,dfx�K6H$�Z��Bd(FfE�)3P"C2�.M:XU�d�H��04��/h�
�Q=a�C�g�'���%!�W��^�������(pડ�p\��ꨘ�TS�U�U���Ky��gӀf���b�x�]���V��.�*y}; nf��_q��n�\�v���Ȥ���@���@���h�����Q��I��@��Ĝ&���SnWu�l���Z<gV�'m%4�<ۡj����d��I���>��\��r�K��l��6�(�y&F�(�ZԷs@��@/u���Z�Սj$Q�&	�%Z`l��0��`{�zX�y���^H�1%88���@��V��{���C�b1H�4 ��/�!�/�o��nI9���fh�� �$�I�}]�@��w4]��~�N�J�ng.�И���l�g
]l��]�,[um�-��d��o\����}3
p�����~�7��u��| ��ɵT�|������l�p��V\�����uz{��>�ՠ}Kw4�\���ra�G#��f��v��[��r�@�y.VB`bM��I4��hR���uz{��uu��Ģ� �Dԋ@���h;�L�z���IEDDDfw��"D�ڐH�m����7;m������^U$��a���R�r��Z��Z�4vm=�GQ�f-��ݲ�6y�v(���ќs��cs��P�W���`��ŷ�`y����yzc���&��g���詻 �V�Z9���E�/6�g�w�k1��� x�ۇ�0Z�X�v�ѵ�m�R��c�ts�d��Lii�{����N ��q�r= ���.9��]aއ^�a1��nwq�df�D��k���6���N�^c�$������ן�8F(�(����^�4��hR���uzyZ�G�S�G$�e�>��\6��7�3o�o�}Χ����)������-��9wW����e4�X郄�1�栜���� ��hyڴ�n�����8��b���Yy�;��;=�s7m��#���|�{2Yz����쵽���
9$��73g ���>��^UU_0��m�ϭ����N�I'	9�}��a<D4(�"��.��s@��^�^�4���N`�I-ڗ��}�g ��w/��IRl���@�?ߖ���cZ�a�
L�2sz�n��=��,q��2�s�b������@��ՠ}Kw4/uzu�xb���2]�j�\rfiRW,����^�R[(����=l�,�)�I"�hyڴ�n���@/u��u<T�s�O�$���;�`d��0��`{+�X��郑G���PNf���@/u�OI!	`�!BH�� ��Ȭ`�� ��M��s�.���]� �n�	�90Ȥ����`{+�X㹦$�B�;[�S%W�	�BbjI�}�j�>������ ��h�i$��)`�9��ӻ^R����V񺗭{q�-����sN��5���I��hR����^�^�4��Z�Սj$Q�L�p�p��r���6���~���-��=疸F)&!
H���8߯1��o���\�����̵na�$Ja�H���v��[��yy�ٹ0@�`ւ<Q|�y�w��}����r�S�q�H��fqp/uz{��>�hԪ[��ܒX����N]�s	����U�m��-ц^�q�u[��^Vݚ��3y,7|�����{��>�hR�� �n�	�$�"rG����;V��:�h^��b�]ca	��I&����@��w4/Z����9z�Ԙ��BZ�9R�I��7��:��| ��4yڴ���H�"LI��L�<�k��f��;V���w4�w~w����p$rA#��Xk}B�7���m5i�����;|�k�
�@4@<�F���m��l]b3�V2	��M���8z���ͬv�J6���wl����۳�h�mɀ����y۞���쉔�n�v��i��7Y�!/uɷ,�^�nm��o&^��*����8+nr��$賹z��^�mQ�Pƕ����v�Y��*8�s����y��w{���rv���)��k�sY�7�3I{OG%�srpb�9񋆹�&9�N*��7u�߾��������9�L�ux��H��$�I4��Zו��<�����@��'����)��$����8����|=UTٽݜ�ou��d�rK�i�*ܷqp5%I=�懲}�}lewKݳ�0]Ȫ���I�D�@/���v����h^����q#s$�Fe�K���nv��읎��5��[��>�Z�v�:�݉yA��BbjI�����>�����@/��.��&9��ȣȢ֮������8��؁��.��4޳@��ՠ}�q�MD�"L���y{���f����@���ֳ-Ie��p�%�<������6��X�i�����;'z�U�5q�
I��}�� �IR�������z}l���J�n7��<Ð�Iy�0�:#rh��Xێ�j�n��k�n�56��S���?�D�-�u��<����Y�}�j�>�c�H�����A��9�L�z�����i�r�v�x�0Ȝ���Y�}�jрz/��*A���/��t?4����`b��޺(e���E���]����02sz�}
3����*����01IyR-�u��<����Y�}�j�/�x�� �[��2n9��I[fΞ +S�uv��5<�n�i��	���M��ަٽlewK�o4�̥��rO䒃�R= ��4��Z�빠y{���kc�c�0�$Wv��Wt�=��L�ަٽlnGj����\d�>�U?�f��^f� 3�rp':ꛪI5W����ASAB���t��T�Z�!!�W!!	SI��
Kad���\�,�,
A��X�Cj��w�}w$秺ϡ3Z�3�m�w ��ܾ�=�����_ ��.}�����q��O7��4��+.9����P�����y���\����b�%svZ��ή2&�z{��>�j�>����u|��7ܖ]���$�v�5UUSg�7x�^f� 3���T��:�^ۓ��$q�QH�~?~��<����f��;V��uƵ5�ț�)j�$�o3o����}��|��'�Mߗ �mnڒ˒Sm��r��;ܜm*���������o�y$�����T_���
��쪠�⪂��ʪ
���*��UPU�D@��"�	P�E�@T! `�$
�,B$Q0DX�U@	E�DX�DX�@T"�E��DXDYE�UQ$�Q T"1DX0D@" ��UAU� U�P EW��
�UPUx��*�� ��� "��� ����*�� ����
���
���(+$�k+�� �C�B,���������(<��;B�� �LAZ A$2�B��5Q@�π      J �Q �IJ%R�TUA QA
��H
$�QH�R�*���x  ���@ 
(
�=˜���@�y�gd
��0$	>x )��{�v1��}o�>���es��מ����#���s�:���� Mi��  $ �q��{}k���1��aޜ�'����������;������|��y_g/��{��W�������� =�֜��O^q�-��)��/�}}��h=�w��f� > �   �s�=>���C�0z�`{|�����7��_,r��J�瀣��A��GA� n��o ��`���:d�E�2!�d���� $ )@唆�M���@z\�� ���l � �=�)s4��΀l{is�t ��C�s /8+��� h,� D� ����t�ٽ N��,�}v� ��  ���t�zɥd�X�e�o :\+�w�9{W �@�������  iCY�(i���#!���[/C'�C��     ) �  H�P��di���6S��=S�mC�<Pi����D�& ��0���2 44"x�U%S�4@       ��U*�� �     )�����J� 4�  �i�4 JT� �F�4 aC d����W�֋Q쩖�^b=��ި�p�$
�3�A���� ��?�$��<	DP��*+�������� 
���%������w����;d��Ⱦ�������w�N���~Pc��f[öW���61�KBB-ށ$��F*��j���Q�v[���I X�I�x�H6�(9	wLv8�d�J�����yH** �i$];�[�|�����Gu���鯯�i���㯱�v��o�s���a�Q�f,3a�a�b�:f,x��
Ù�>Ȱ�+
��0�0�+̙�y��řww���3R�4��1f#�fds�8j�
�UZ@M���˻�ߑDr
*��Q�"�>��=����DL����,TOb*
{ �;E	��'��i�=��|�I���y�n�Vd?"m���V�d�2�\�vw������N�'�$��M_�������+����k�Q�3�"}]�qf>tG�Z����������ۘ�B9�;�3�l$JW���D��A)#���$�T���9:���:�X�i�(ҧ��:�اD ��
�n�S������N�y:��S�9����-��`�C���.~!
�k����8�8tF����k�7�D��7����$������E&�8X}T�lu�ya��Rᛇ7�8�,�N�����H��N���7;��v�Чh���B��^:l���#��
F�:!�G���9�XD2���(��w���"��;�Ylnpd`�` � ��NW`�������D	|/�:3�'Һ.@�DG).\b.][�V�H�qw��q�{�����0
K-�,���v��'�	�΋�	paB:�,Jb�\#�ư�9���,c�L`a�=���)�ﾼ��a��$$]1�H��Ma�{�F7���Ð�
�3��7��e�N���)��p�8]8��N�
c�9�F�d�05�0��Jx ��[����;z��j�2JbD��f�p7��k$�0+���]y<�(��tB#�1`"d�����a#�23/3��9���B\�7�S�s�@�9H]w��X��@��`�����7��0Ӷ#i��)��	�wNö��0C�V�S�w�b� <a�}�6Py��(0S{AA)�d���{�.�@�����������e�a�`) $���u@�S���'@�6����D���|�9!т���@ѣAF1���:�S�q ������LHhP��Б�$Ȑ��Lzi�9�B��MI�Xa� �u�aөĂb@a(D�0׉�^H���hCNt��%�y�$�P�Cd���7!�F�L9�s�;ӹ��U��.!p�d޴�S�7��8f��h�L���pÎ��qt`\ٷ���x:���ps���9����ѣ@�(�#w��$M�8Ct�{e�s��օʐET�Ύ�-
aS%��ŉ;�lVX�D�j�X�@"H1p`�1`E�Y �VJ@q$�����h�щ�E�$$�;b�Ԅ,(A��"C� �{����t�$�a�Y�s4 Q{"�P!�o.��|���OGpa
&H�X���d��t	-C�(Y"IX�1�BL����1c%�����JÊE�*`�Ǝo��n�����@�88H�b�B|�����¾�X���ˆ�r�K��5�!L�^HV��K�h0H�"jW��5���N��S%�T�W
oS�����iǪvJcM�/]�#6p�+�ƘSx���	����:/d*B��t�
��)�����A$��������%9�-�S�;{H�qLD�Qd# � V`D�ԑbX�$C%��Q����H��@�� 4� �Ԛ=LJ'1�/���f2\&8	�A�(S�9�4K\ �.dLȏ6���v��{��A�����=�w�s�v�!��{�o����(󣇊g:.�Qpfa�/:�ӡ�
nS�KӽKݬp��ÿ^����B�u�àJXaq�.�A��!��^�6����*�s��;�!9�ۖ�d9\�18G4Ύ�4�!LX�D1�0���N��@�
a���Ji�
�0 �/H��^�H�	ƾ��X�S2k4
.�YV(��1�%RuiӾ0�sF$u 4��J��-le���)����a#�0<|u{�Lӄ��S�Wj��#��X�B�z�󝘂ڡIdy/�Odm�����P9˵ԈR�P�0j�C����/�Lp˳D������0�޺5�;T*	��!��]�I���7�I��1s���$#�<�C[tID!|]��d D�]���C}��X��XC�Qk�țM�/K%��2
"7�9�ȸls�/,ErS���xu����1nCXX��aB��&�
a5,$
��5�F.��<=�� s�� U�R,�R.ƹ+}	7!�CF!C&�!�����$&�zq��p3C�ۄ�}�Oxy�E�D��+���e:�Hî%r@4�������o8����{o��H�U)F�P�}�D��8zzGo�=*=�Ö�yT
v:8;�h�F����p*�"h�@�����P@>Ns@C�{*`lJ9�'���j��(Į:��<	q���`0ap�Js�k)�^)Ѳ@�2ᬺ�La�a��D��-��N�W�(	:�!!9ޝ8��`P�Y�=��\7<:��М���:lX\	HaB3����	H���j�:{z�|�Qk�2H2��VWf�8$�eu�$	G7�3�!�;'�]0��Ӥt���CԸ
��S������d��Ȼ]��|utz�������4�l	9k��0tٺ#LE�˻��.�!D*)�	�9؉&�N!N2W9�q�q_T�
�:hc�XG��������E2s'\*t0FfI
�����T�p�9<��C�.vt [s�+���u�� ���z\c�tw=�K���_q��ñ���9O���`:��	(�`�6Yh�`�p&�t8�q��^�_8���B\��\a�9y��,v���� ��r��}�4������:5l�h
�@A�Lv�0@E�`���A�@�TC��� �I��O�~���	�8�jbi�88't]J!�RU�� Y�8	CO{4��0�δ�D!�I����(�#7���������Z0�t�a��\0J��o4�s��gk
X�;��םkN>,+paa�e�BS�;�;ÄXa�ᆈB�$�]�+��8��V� ��$�VB�ٜ���DBr&F	� I$F�Q���C�R��h�$
F�8GLx����0#"F�kV(�i��R8jD�:G&+
f�aP�&�@k���70���=,)��9^��˯�t��L�N�xt0��/\�И0��0�:S0��z� �g��r��L�
 ��[�p�s *�6Y	���d��ھ�9;��(>ql�Xa9b���ޛj`dP�X�M.j�
����qgE��9��5j*E���{v�	��bv�]=��h{y��86�e��a|�Φ���7�RR�Gӻڃ����i�O��Q����Ж�3ǯ�$��>}����O;=�q>�/����{����w�w���__@ �     -�  �     m�           ��  � h              p$   �`                 ��       ~�|                  8          >��         	kdnq�h[@-�km��J��m[m��me�h�` kY�l"���8��r]�`               �  �                                                     ��                0                                                           �|                                    ^�����o�>����-���Qf����hp�`  I�n$���H\��  �`��Y��%�p!��UPU]O)�v�4�m�l�M�� lշm�YZʮ����I[�� �[f�-U��%�����Y�"�7u+�מ��6�`���'�۾	�C�vز�+�UU��)�+���8Z�lbB�[�������Hr �jU���@u��6��V�`����U�^B�IN�  r��[k�����M�)�kV�t��I�btg.�H���d�.[�Nk2�\mU��a�J�t��뎜+]M��6�5�i6�����U]*�s���7�U��R�ۻ#�W���*Z�"qe �5AKR��C�5�C��}$K�d ��f�6����l]Զ��a�	$n�H ܵW����m�Ē$  '������[bj��@��hփm�lӮ  ��a�2�-���<��ƫ��Zv��a���ߟ�`6�+%�:��k�6ڀ���'A�ʵTq��l:B�rAk���I!��X֞�{�$�M֛=!a�i5���UJ��4)��V��{�v%�#�1�p*��L�q� ;/�ah�X6�cp����|p�[����X�S�C�n�q�/lIcpgb��{=�5�
����أ\� x6wPx�<V�ln�K,V�Ҳ�[B�]����,���d�U�0  '[��
�[]U/�I���V]��L���s��U�b*����jv�cg&t`m��m�kz�m8��Ým�vvN)ɑM�uUU�X6��i�Lr��  	m!i��p[���f�ު��m��p��XL[P-[lpm�n����ۀ6�`$8 $6Z[I)t�X�5�Z��Sm�ZM�u^��q#m&�v퀺��l۶(���� �$������V�9'+.i�� ��𼭫n���j�Ηi^e[�c����IŻ�N��[@H�+�R�R��&�E��E�Ij�m:]�А�%J�u���EUʠ/,-��e��U[�5a�@$z�����[[d�3=TmU&��+�@mV�]���ر��tJ<��ݖ{Pơ�t*�,*�*��s�G5�f�x�V�TFm�/5JKR��I'mïn�q�k�[%H$��v�E�'��g\3����~��[/*���Kz� ݤ�a�K4�m$��Il��7lf�T[O8��
��U��J��uUuK��7;b�$���'����`-���ۖ�J�9j����Ul�Wm�$m��rt[@�^�U*�W�Z�W;hԛ�ӣ�ۘ[]%�gm��`  9�lM1�� �87m�b�%����h ��	    �� ]!5@9L�p�UM�.�Z��EU��Jl �m�/i%�i�.�    � ڴ{Y0 � ��۶�  �m�l��� �uf�+�M}3
���T�UJ�dVU�&�\k� �M*���`�m���H��	6��-�����lpX*�Ij�� g���I*�����l�m�@��[�I�� ��kZ��	6�[K�&Xj��.�%���\�J�:R@�� ����f�U�۲մ��dΦ��y���U�$��ݖܧ*�ݸT�bZe�;i�Է>�8�I^8��]6�$�-�K�r�lÍ����-9{N�l��ܺ3���˜p��m\�kj���>�Ы�l�\U�Ý���8�̷i΀���G9�=vj�����c=nH軪�@l�\k�ک��Wv.Lf�뭽�æ��眴���^٦��u�-��r����� �Y�4PYĩw%��K,�5I �m� ���[u��	$��ͱ6�Y�]�X`Hm�  �)$���d����h��NѢ�5*RK&��%�[�`���|4�6al�Od��(��j�l�;A����|��Um.y,�OB��ln���[a�N����t�MВNoE^njqz�;K�T�p� /n���cn�[[[u]��PUZ��8(��j�u�.�U@H�gҽ��5V��3*���t.:�H��r�)m�z�o�7Peu�@t��^P�n�����8��=�v��e]�q��e���eN��uM�k��i�
UM��GH7=�*w��Z�=���W ��q+�V���1mR9� ��jH�l�{;Of8N�N�vml�o ��l�H��Pa���UUR�=��R�UU*˲�*u�3MŔ�#N�G��[dŲI%(m����p��t��`    K5�i8�� �m����m ]�7K��[ri5�l 5��&�O[R�p 6�`�� [[l	 6ҵmT�IV�b�_U;am��ij�i����   	 �am 6��auޝ��ʴ��uJ��J�T f٫u���h�$;m���H]3l�'z���౏�	��G�I�ӵ�J�U���B�U@UW���mշT�4�e^�f����/@,�`�_��Z�����V����m&� H[� mJUN�,�kM�   ���m[B@��nqm���;m!U),�4�J�;kn��  ,� @M�m��M@6�`��w��m_5Ԫ��6h �� 6Z�[%䅳�A&��*�P����g�}*���l@:(
�ڥvj�\É!��u�h	9m�dІ�@ZE;I�d�,�� �-�A#FV�"r�R�]]��ȗS$��l pm[ۯ�*dm���(�R��w ;����&ն��S����� 1����,�9qHa�T��p�@q�U~/�R����X���h��p��t��`��:�iM��	V��q���(��ض�g�zj���Kt�4��@^�z�]I�
[sq`�P9��<�Tue� �8Km��T��y��h�u�tPk+�ܑ�:l�g[čY�G����٢��u+*��myM��T�u�\������w�Ϫ�����s��$�$��f���^��֐��$����GǑt�,����wg��������2K���GC�����ս��w�|�6��<}������s��g����������{������������wwwwwwws3333wwwwwvI&���������������������AB�
� ��z���5G�� |TS�<ȁ��S�R�r��(�8�X�=��"u�P<�_|x�����G*���^�d��8��3� ��r G�C�*��`!�!�@�� VD�!��,"H0b^q'� ��!��v�s���\� ^� )�;�B�ׂ� ���hj��EA=Q{*�t.�x+�T�QJ u׼D0�;�ΐN
�E�D�=
v�| 1�L��� <뮶�k��$��*���A��-Z��<U<���@ �W�_E��T;��a	$@�C��B��CU4�j> )�"���*�|@��A� �1�F,'h;؞z >���UE;����U ���P{�T��P�� �:;��n �(�4<=}��n"��*��Qb�߽
���<�]z�AK�#���P��"H�)�������EE&����B]���H��T����
������@�ή�(�A4ڡ?����'�-�!,��Yw��=�����m�� m  m�I�  �6��   � �`[@m�� �UxYL2�b����i8  	�         ��              l      u�D���ݻg��C���[!Ю9�c�������rl*��͸���2���Ჸx�.��6�%9��!n^^z۵8vM��\p7h�!m���ڸ܄]gt!&�v�-v��.�@g7q�C�f�����&�x`�c��rő�҉��d�,^�b^�k�8���Ԧ�vd�cnɰT�ڢ^ێ(�uvV��c�Y��v%�V��s�N��2tp��Kp��p"ڴ�������;������n�����]��n�������*:������CA�d�m�77�wnR^�R���k���v�K��[�ET�7c6wj˭����23�نF�����U�ֺ؉�x;�('k`�շZ14���v��d<f���e"Mm���nn�{CQ!�T����8�kd��4m%<�ݥKK�U����G8�i^���K�rc�v�$k]���ܤk���>��\k]�qu��(un���k�j��p�2�r�M\�t "��&�Y�c
���+�7�!�n1cͲ�'k*g'ntw\ە�\]�8�����⥓���Z���V��.ݙjUUYY��Θ�Fиgt�h�����mw�6H����[�/;�Ҏ��b�La��͛']H�:�b.��c��M�q�Vr�Mą��=�G:�yw���|�r�S�ʧB<"�hOUC�*�����"��7�:G�~� v�uB�;,��[��H����sl�; �Gk, m� m�4�L�k�Uc�6x�w�����Rlt��nBc�I��r�V=i��κ[H9y�= sӝ<�3j���ڡ���ێ�]9S:���=�\�G[��b�Gq�N9��e�oN�.���N�Rv��v���㮃'u�ܹ	�C��%z���\�\�33E��"8����n;9�t��M�t�bMo�J���W�/~D�α6��^d{�p&ی��W~̌��v� ��ZA�'��Q���fk#/29���r�Ҭl$���{�Y�Uͻ�7z��n�N%"14�o�j�ws83<��r��R4�	nI$�|��Z,J��]��{�][�ٳ0�w3v�����DO�W�������p��*�r�m�sne���=��A^�߱�|8�~�=�� 鴼�ƣE��N�����+���`]�Xx�����I80琳�̃0k�s�%rţ��܄��j����u��doUn�L1�I%F��� ���ػy��λ\L�,�2ml�d�e�f�3�pY�\ ��Dw�Xz	j#)07��Y�Uͻ���`�Ө8���RM�a�U̻��H7�*���!�r/0&{Ҭ���%Ș���(Q�n���x�ܸ,ߕs����k*8�*pfk���pު�v̮��-�?�$������o>m�ɗn5�,�`/<��s�;��Ę�3I�z7���X��]i˱��("f"�NC��U^f�����\�h�1�!1����x��  ��sʽxN5��#����9��e�Af����0����>zVYZ���$�����]��;z�Գ5礷$�3h��rc�v���A��Z.:�Y�VW���a�sp�wʻ�܃���`��m,L$\fHX�������o2��\��m�Z�R�|���̃��=��p�Z�X�EȘ����M�$s�pv���v1�0D�MF#�wz�]���0=ypm�T�6ؐ����H�`lSWk0     UX8��X[7<��u�7g�+,�;F���y̘��ݓ$�C��{k�,.�g�\W\��ڶV	��i#�&Si�*➻t%���/=�җ�^ݻWm��ôI�ђ7𹘰�n2�l����s.n���������㟀�����tx�������;h��YC�͉�=�M*¶e��iZږO~�ރ����:ꭼ'�Z��Q�^k�5[��p�s���J��E���$���t�*�v�oX��Pq)M$���Z�.w/�����:v���N3$,�v�&��`K˃����WOm�}� J�f����c�.�CN���$0�@h��{�6�@�*B�S��X����Z| v��t�^a-qԍ����uC R-F@�H`@X�5�X��E�H FX��łH %B4�P�20��FQ��*��'C���nNް2�c:`����G8/��������W:-6�&G#5��o۸;kMm�8�"ӌ-�^k;wmi���A"�"RI$�&�k�y�#k�u\��]Z�ܐ�GD���z��{:5���̂�Y����`s��q)M$��Z|F�d�tO�w0��%���qHP1���J��B����
�C�y�gU��=���Ie)-N^z;wmi���6V��8�.�lY� �m᭼�;x��v��h��C#$5j2Kt�`��;��f�a�/��$�I�`����G8/������=T(�^d���|m�L���=��z����gqV�1����B�^�3�pY�U���vU��Y��Li� (�݃�v�	�8 
��t"3{�S0�m%�#wgn��{w�2n?uUW3��s[�3s�v��uv�0����odZ�ӉD�M	�ڭ��/�����gq"9���@���,�835���j�v���^a,q"�F��̂�b�m��`]�[:`��mD#� 
��*�܂��[UB�n���|i��5]� ��s.:1T�:��o$�I)�m�����     +�[�FJ���/fzb,���y`;s�i��3Wmu9s+��d6�Ļ��h�{73vn�gFv68�����ݭ�;g�v�䜾1��lj��z�)����DB�Nt�����M8)�xqi4�ݸׇ�,��']suc/��{�{����u�UT-98�y��m���s���N|��mZBcF�fO�3X�pY�U��ʻ*��L���&���*�C7X�~���1�;��S���F�|���s;sN_��[�t����MHd*&�� �lz��]�0��w��h����+/]{6�=��א]`�0��M�$�ʝ�ܛ=�Ȩ������e��R�+���3b����W�^��_V�E݋miB6#.d�wuʫ��e� ����d���a���ƤQ�Q����:��	��[vN4p4�0!�e�so%gq�}	m�\�����
�n�o%^c��ܫ��P
�l��$�A,���:{su�Ův��ҩ�5#��T�✝ش$��W�~�ם��-k$^����K5!���u�y*���ܫ�~U@�ﵶ�:b&B�*l����o���k�si#�/<(�OVo{�ͭ֔�P5c�����dӶd�)��;��M乳�Ù��4`6�D��B^-m�ћ�SB\��&h�t�7���q	L��o	q܆�ڭ�C@RJ�fT�$&B���Yr�4�;(�1C!U���[#
�t��\��.l�i��ۘC:�q&`B��H1!�c�xp��JŅ��L2RI���0��a�1)mII�tK�p�N��� H���}���a�i �+
��.���=��﫼=:������s�LͭB���	XE�*=�� �\�^�נ�u��ת�C����Z<�i�T�Uz�[0�����zJ�c�
��Ɲ���u~����:����#b2���9��y���y����}�͢�Ԗl��I$��IQڅl��xC=��p�])��R��Z.���Eo�gZ�|��񎄒G.ٮnW3��0�LMK�
������y+=��ݸ�f���0("�V��_ٺц{�>���w�bpt�6�0�^���J��7�EU 8�R$ 7��� P����i�KS5���u���6���f��B�õ�,�G�e��gò�<]��@;j��n�A2�	�
������[�m�Lh�V�{ߟ�7�g��ꪭ�V�͖a���^r6()Do���?yV����698Ffg� ��˅�+}�\���2��=y��|$p��qE��f���\�[Pi�kD{,�h�h8�D�i�[��Amo:��7+�(��2�
��g��v۹$�)�6�F�rZ��&��      U�ɬݳ���j���թC�^��e��b`��;�S;-�ɹ�.<c�ט�iغ�m�b��R��ړiׄ�s��x֞} v�3�٘�⣔8��m\qo�_G�0�2��0q]i�Y8�3�^�-me	ԛ2f��0�<��������Ks� �Um�;Y3IX�Θv�x.wV8z�4�R�>���P("�_f}4��u���V�g��.8XN$�o�����!�͜�7~u�U�f���KSE���u�͕}�6�=ܿ�����6�K�A5֛�f�%f/j�g���GE�B�$#�ټf�$5;�-s:����"hc.s9���(iwL�7h�Z����/c<�AP��oD�q��7|�#b2�FN�>��Y�������<I�kꉒ(� �g�ٝ����H����M&���˴�̔�}�Շ� �>�'Z+INCb)ρߝf�A,5~��vU����Am��87�[���x�m|Qw�rU��=5RI2$�|�?���V�ξ�ۃ�M}�KuT���[�8����puv񸸮պ.͉�s7j{J�F1F}�ܟ���g����M*���M--D����[���(Q��}�?ϯ ��_0V8Q2ɍ�z�Ň��Tw$�U�0$��������\��u���lF\(��� 5��Y�3A��MKq��yf�d�>䍩!p���*���Vz�<�� P�����UUF���/X@�:2���]�9�msR��O�XF�br�D�[�f�%w���w�3
�}I���}�j�W�����(��>	��H�m�w�?�#6�V_ίݸ=iZX�1�J���p����אp`�(5�OH�_�i���`���[�cNm�妯ݹWv�h��U����7na�6`V���"TKg<�&�Mq��ؤA%�o����_���@��]p��^32��J���Iu�ZuVnl�W��f�OP"�j?B��6���[�l��1�
�z������ak-� B'���rM�o:�<�3hJ/9�k�������e�:*I���gUg͈��mo��,_s�j�uOo��~ՠ+���U��4�v�#      =aι]]��R㦝�9�(�;Z:-S�7�����{x�5����\��$���w�������=Q���g��d���O��۱�D�Wf�{��l�:��"��ѯX��.M����sgs�OWS�4�m��0��@�1���U ��K�%�$��������m��t��h����kVnz�f�^����,q"M��9�Y���ߞ�P�A�^pY�%��QĚ����o9@D]���f;�T ��
b��[i�<�0E!��~c[��`��A[ܭs:�;f0�q��fC1��*��ٲ�u� � �F�γ0c>0F�i��n����s<���mJ��X�o�I	�J!C^^��-/Kf��9b]�t�ۑ�ﾫ��Q2H��?��o�����}y�C��n���:��Sr�O��nwZ84�� cBի�Ii ��</�]��^���X�E�0Fo�o�en�TsאY7�0�g��M�XR$�}�>��f�g*��_y�̓�/&��R6ސwټ�7z�=y+ٌ9̿ѓw�ꪩػp�4^�ͻH�WZ9�%�R)g�������M*�TW%��^��f�'���&�߾����+��zD����u]�%7��%o������(5��Ӣ�i�M8uV\�'Lα��$��'{�R �X+���ku�\�&ʊuUP��%�(޹����r���� �kR�xu=I2���"|�3<��(UUUV�7����:ϯ&���=�I$�C%(�ʴlZ��'U<w=z�/B�(0H�( ? ��L��(��0�| ����V�}��W�8N{N�ˉ�"M��#��0
ͼ�Y�����
�@,?j^Lʎ%#m׾�J�q��@��f����f�56�ZZ&�����ι+[γe�jN��llI"�@�! �������@��dJH!=���_��Y����	�7Vo�e��@ ��!߳e]�������񢛒I!;.e8�X�s��X�F� N�2:*	#�h���Y�F7N5�X���#6�U�� ���*��*DԈ��>���(|j�9��k��.g3Ҷ��IP�����.&j�O��~^v�Љ���l���LӨu$��:HAƔ��-�re�ͬu	$��%;�{ ��.*�&fl�������ur�9���f�$�3��gn�ªtO1<9��dQd�A6�B��i,����F�v B永��搦%+6���L�; Sw{�y��[ë��xq��{�#0H\U���4`P�B�č^���4��b� ������޺�)�J���fso8�Dd��s��IVH�qaQ��tH�HT����4(B
n㆙�λ���9sni�ۄ�l��w H@E[�I)��@$I�dB0`�[�`@XfT1�]�4 Ǯ��/c��Va��Ęr����Nr��/FF��}��%���4`(��*@ � UAs����}�y|�s�w9�\�#.V2�xjd+
F����ԉ 1�#�*@`�&�2i�/{P�12�!ʡ��@�;�cN1�=o�q ���B�:�|�`�
��U�$YG�|5N9a�%1 �e*4*1��1b�M0i�|�-W'�Xچ�L�C[��]|�o�p $   ��@ ���H   �  -�m	    &�Lݶ���%UU\ $                                 .�����x����{9Ūq�ۧ�r<k�V�ۋ�yLj��{H�����%���Y��N�>{p�9,��nV���X�X�G:�E��6���e6|��P��%����Rb d0��X�p&!�m�tqP�a����=a#^!���ٽz�[�kv�n��M���耋c������gdL�U��l<���<�7X�E�������k*s��y�n�5p?;f�ϰ���o8��:��fx��	���n3M7����'R��k�����[�cd7�ϴĚ� �2�yQ��`��}��V�@��h��լ��s ��ƻ$H���j�6�N5��jsn{;v��v�mF9Nx\���۱�F�4 gn�U��������<��\�y���Yv�j$�5��ճOd�@N�P��}\q%� j��d�Cۄ�S�6����m;p)�۱n����v�wbeI�sa8]�I��!�c�2��YC�*��`����v�ڨ�d�pЇ]�H���9��|m�c�j���9S94���GH���ۮzq�t��+�<��Jͬ�$tJ��T�[g�s��c/i���fr�3̛�>mQ���\�kL�n�.@|���
쉍�g.����,7fY"�l�f�m�6��y�玢`qT�L�X�z1��3پ���[ �H�Gz{E:�P�CC�N� m^��I�
zޅ\�G�a�T�����*�fN��3Mݛ-2	lr�ڻU�      �ƻG*B��\�gC]����c������;����nX^:8��^�s���m<Z5s�����+�7W%�Hx�w�goW�Gn߽�m�]8���q������P�o�}��|;�iplM�Z�(gu��K[��$���zƄ��vW�ׂ�pr� K�h�$�I q��'7����6��y��R_O�/(���U���w��>�,͙~u�Xƥg;�h��G+sv�3���J^%�M������+o ���3ٳh5`��^��a�}�>��[_U��W~cN�V�g��-8x(5�N��I(��+W�i^��I!;�b��6TS�ƣE�4���t���6��z�W�{�;��?T5UApU��%�=���q6ș��=3ѵxP��&J�M�J>���:ͼ��Ǡ�לx��#m��^C��c�`	S$%j`2c��F�!lq9	���ׁ4x���p^�$]N$�ؤI-V���T�}�h���6�L҅8�m���[�y�P��_�^A��K8�q'lh��4Ad޼#=y ��^���&�Kİ`���Y��՛ܺ�ۯ�j�J���&�FF��/E� gcNʝnֻqc�φ������V>v>�j�Ln�ٲ�1����
� k3��7tF~q��%8Y�����ꪯ����[�����p��>1�F���ٳH��=ꡔ|n�*����W� ���Ċ(H�H�;��ٵ���L>f^�[�3T�c�������6Wٌwh
�ټ�-�)�E��u��6���a����.��4nɺ��*ini��]�Έ�n��Bm֐���-�d��x�lȓ�6�k��7�%w�_�UQg�89kؖ�iGq��}�6�
]���f?�� PC��&S^%�M�Α�����6���u�f�uTzW��&�Ku2l�#�āO:�
�`�9+_�=ܙ�@o�yEN ��H�>e�+��K�C��n&�5[��w��o��:`������ֹ4��Y��}_53�۪�UU� �����]=�)��c��7=��|���Ԏ�8�hq�Po����廛\ �M��ɦ�Z��K���j���]�o�k�	�LO���~��w��7�UW�M��[�Bc���۰;�P35.�� �]��F{L��DS�(��?��P� ����Ny鄟+��	�UP���q$�{���(�N6�z��=0���
�_	>܂ {1�-��U��𵻒T�!:oH�Ũ�봱�     �yۍ��c[(:�ΜmW#��hҶ��c;[;����
�r8�v�N��n%������� '�(\kv�uۮ����m�����#-���q�{�6��8c�Vq<\�{Tlm��OA�r���{q�w7�����?��=���n�[-Us>Y��km�vM�/�+��}
1=���F��o���6+D���������$n�$��U�į�$��Ey����0��w%K�}U���n�3�H��I����JD'
rU�{�sR;�˧؀�@v�4�U=k������*I:;<?�����w,��{mAW�)d�m��y��|��lY�-�bA H�s?}�u�%����޲[��:�� ��������W���8k��m�?����ꪪ�����8�2��*j��8t-ni��ٞ�#�B"�H����ܹ��f36Ŧ9�)��}M6���� \���x�NTR(�I6��?�c��"%������fp���6��Q]$lI����q�LEMDML�ٷ���V��1�����3��E6�7���k�X�ذ�n2�i,����P1/n��W�.za �4%�-�#݁�ͺ�?~������� �'��f~sm���;s��UU�8bg�qD��\�LӰ�SW6��J*T߭ʶ+�I�'
�W${�p��	'���@WKװs���<<$�@�Q��|$�3�UB�UT�9�p��zT�3f��!r�r��|@g;�m���+y����Z�m�oL$��W��N8�a����*�` ��� =�8�} s[}��b=����F�MՀ{u��/���l��;�8������frI##���HP�݃ۮh�v��d�v: ��S�{ꯅv��Di)�m��� 9�{V���Pۮ�LlX�TLԻ6�1��$Sz�[��Y����?%ߞ�
��USg<�KR^��"h����* fc���� �|����bR!8T��?}�U,��ׄ ���>?}#�F@"HHA�`I<���MT�(��.��N��Ԓ�Jq��QX����p�J�qn(����I$�DFEQ��q����у�юu�\Ըdy5��wy~ў>�kk�ߍ����3�*��^���A�< ��y	�Ct�w�ݕ��U�W�����:m�c�[BA� L�sn�4��Q)$�X�~P��qm4w?8{=*�{�D�L��	��\GE
���L$��ps%@߾���<�T��cb�tJ��� �y�%���ܮ��j�_�ٲ{{<��T�#*!Kb�w�����~����(
y^�&���v�k,      	2u��kW-�ۮ�˘�����ږ��)�X�#�9��{�G.;T�vG�+�rZ%��۝1��nv�?��p}n-�X�ΝJ��{o6��@=����'I�8IV�Ĳ���1t��ĞH��A%OZ�hG��ꗝ�w��T�75��U��v3s�W0�m�"L�.6�k���{����O
*7�3J�qf(�} �^Z�0=���E���p���O��� �~za$���'��@ ���������j+�z@�8o�{�*��P��È��rL��T)���=�tS�s1M�@lBS�[N�x˘��q�7M�`~�ʀ?f^��;� ���=_}����FF�J�IG#��N�˵&���s�1j��W�_��{���ͻ��/~0b�����?Zwe@:��Ъ]��ˆ�^I:�<�y)����T_``�ۄ�Ĥ�8�ι�<Pv/��'<�6I�~脞�b�СM��2��E��I��I'�|�v�~����.u#�?I��/�Z#	Ȝi7�~��T �~脘����} {ﾪ��g� �u����n*�U���J ������� �y�=ݕ �.$���BF��O��>�f7K]v7�<�ʶzL�枼����ߏ�������[����3V����P��ې%D� �y���U|����.�_�I�_����$ۨ��۰;��T�g1O�%m�X�(�:�:��F�w�u�#�g��W7ty��GA�i"��G30k���2�I
`�˙��
)C&i���$�+�����Y|�%��e�xƱU�v�FU0fY���tx��f���$��L%ax��R�	I��H<���B�`{p�	�Iq$1��4P%C���fE� �#
����(B�/:���ōM8�xkx�1�k{��[B��#�@�3Q]�����U�=@�W<�T�Q��S���
���_-��$M�I��5�T�)�ua�������?~p�M,���v��!��$��kE�JB�m�s��c�ms%@�p��+^����l1�N�����%u��s<�K<\rO����)An�Jj�n3�Z������ �n���:ɿ��IՅ/�^��M��vT�A���< 9�6����U\�뭧�1R������k�^��`�� �2TW��r:���|:��P���w����N��8b]�A	�R�(L �p��,R#d�1 Q��/@�A�5�V�LC��N@��Z��%�������p�����+�Y�V�M�* �$����U�٭��z�Av���[v������w��k�I&�n�o ���@�p���<��\@n��74��D�MՀ{u��U|��{��3<��J�qw�Є�F�e���'��W	&�\>�)+�� =���,���Dܑo�-��q#3ҠZ_�Z���ￏ����yp/	~I~����Q�Č͕${�pk���$￳�Y'�A�"����$Z��;�{���m݆�[I�F�b��X��     ާ+&Z�n��N�8��jz�y�Mn�q��3hG��^�k��Z[K['&��n����!v�ޕ歂�rΞ]Q��@Z��o2����n6Z7���b:l�ݺ���}�#��ә+&0���x��.��C�#>���t�fL-U2��P��^��(m�u��3p<�ש��$�� ����2����u.%�����V����>��� �����#k��u)��8��~�W�}�$�pcTSm�9���v4U<��9��D�MKuQH���ps%@�� �y���n�Sq4[��P3��wu�/�1Xm%��1#v\��$PI7V��� e��_}\��\ �y�7�۫�������g��UU��h^h:����7L���E�*6p�lN4*��M�m�h;��+ �u�܃�@
Iy���'��mk�p�ݼ�w�ټ��� �*Ȳ,B�f�)TYy��|�O/~ݒs�1gtU
��^���mF�I�����U��}UIw����f~p̕�yJˌI�GG��U
�}ߋ$�_��I=�=H�� �"R�p|�@Xp'��s�ś|@HD�\����M�Fs�V+�H6FƤ�I"QP����[3����z-���-��l�+#��tQ��~�_���d��[�����<�U�l=��M�m���?$j�J �纬�󟾪�H��k�8��	&�����]ٺ�Z�P��:V��ԭ���y�
�tGj6�������+ �y�9̕���u@8�-�]��DܑX{�(UW{�V��_�b��ҿ[��v��+�5��q�㱮ȝn��V�sg��S:���\�ڍ��J�H��mZy���Ng�$�e!#*1$!�~�9�uXN�@9̕�M����r:�:r����=�ך��^f]X[�bG=�4�&�8�TR+U-ɫτ��{���[�9�8�Jê P~�����kڒm�l6߸�3Ҡ_V��`s�uX{� �~��������,�gy,�v��@=�k��QI�m�dh��P�$LI7V�� �y��;�~��ʻA՞օR:#��V|���H3<��ʀyf)��#����%$ܑXg���P,����VD�`���ۍ�{���� �<�`��F묭��T�QԒ�8����l�\ �y�7�۫	�  /q6�$H�JG�����%����     V$idĖ��<4�+���r��3�Ga�y�^����h���θ���:Zt�_5q5�^u����gc�m���/>��9x'nQ��V����)ɳk��r�gp�v�ƈqaHٱ+0�����Y��6��{B�
Kjco�p�
�`#v ��s��l��c���0t�z�s)8�����;�p?.�K��}�����|5q�J�Ez�f~p�ee���Py�ߪ���ѯy$�n n�n��Y���j�P�o���fz�h1�1�$��&��/ʪ�������o�
H�|�?PK���[��(HҎ'mp�=��6�UB�o<����,�s�}��nI$�͍�#���vM�3��~���b��̌\�l���r�,���6߿���/�۫��Y_}��V��y��%�����L˹����w��oK "�Hq� Uu@�T�qs�o��p�M޿q��kdcT�J:�U���(��+?�� 6.� TF��ٷ�r�m���$�:�*r���@�����3<�̕�������s٣WLq���VjFg�]ͺ���)� ��`g���u���ͻF��E�nk���'�Fԉչ�s��������|-Y�6I�6�C�7��Z�T�>���>��k��I"bI��<�T����US��X��5#��P?cB��6�(ڰ9皬�Fg�=w����,���BB�+�"š(��j�� o3ϴ�:�T ��>x1�����%�-%̕%庠��V.�y`�mF�F�WvT�_W��U��<Z���U�0��RI$�m�ʑ>n�B��NȨ�A@�T�B1�q�I*Ȗ�� �<Ŝ@fk�}�U��zTWQ��ڄ�S��V<�U�_�785o��带UURIs�h�#i��J��`�p�J�yf(��/qh���l��q$�͛�`B��r����Sn��=��r���s}� � a���l����!�e$��'�uBO��UP�s|����/�*ϙ��ܒH��A���n�6vŽ��NKN�j��|͊Lu2�A)�ך��� �d��� ,՟<�$"n8�O�Y�s�@${{$�n����ׂM-��4�r;��T��g1O�1Ug��"ͷ��4��1��j�b#�%X~_��Pk�Vu!w��ox!'�����q�{皸I� )n����>�'庡&�tP4Y���8�Ǭ< bF�# �5#1$*`�Sb�T�
$UP��&oԐ	�$0	I  0�@@o\Ρ����ȪA*�;0w��%��p8m  m�  lm��  �  -�m	    �m\��e�Mmi&�Z 8 p[@                                mݜ�\˧��̖�au�TlƍW����vy��]sY���6�N�7HM'@��sUݶͷ&œ���@�〚���֞wLldu����a��6�5��qnMvN.�Kk��Z�ۣ��2�+9�1Mwk�6�����v9^�wk�9�ku1�����Rf��3�N���MZ��s·eB�7Eg]U��E��#���*��5���ѻ\�2��ͷN��-��=	�R=\�K!nRg�&�����ugH�Xۓy{D��u�s�����r�l�FDHj0�b�����d�vnQn�j��Y狜q���5+�G�j�[J�h뱱u\�\��FC�уB�=�m�� �{x��]*�k]�4����M��-r/7H�<�Аs�5��ոY��[<v��Z.��Ŭgy��݋/0�;qہ������EY���i%�q� n�u���nt.㎚�`��a��:m�dY^ޅYl���ۍ@�tc�A[�j����8����ze�^h
����/Y���T]�i�] gΡ<�$�x;"ri�V�ɇs����+6�g&E�j�y��<��m�v��yf�uV!C��Eݫ���gg�i�y�Іl�&(�zm���&���\�/�M�����ȇ8���Gl�!q�������J��#�*��� ^��ޠ�5�A�����f*N�5 �@���{����f{����n�m�ֱj1��X�     
Ji7^�;n�E[�����5������,M��-�r#���p���-�ZYYwb��0������n6�^����Q[��s�m�/�a;M��VرY��ߋ�|s��A�V%��;�.���1���ѩ���e;^v�ko�y着�:<Lp4vwcl�����-�cl]T��(5#i��J�ŀ���%@�b�}_}��5X�^<��%!:m�6���|�;��'�y������ꪠ>���������)�bI����� �}�Z���̕ ;�hU����Q�6o�	B'<��m�k�M�_4Sm�9p�Y�)*����\����8��
�;���Z�?�I.0Wc7V^�Z���+����=;e�2^����|��B7#���H�fc�s��V���+��#-Q�9��I���U�ZPa$
�I+Am��HI ��bv�ߞ�����>�w�qX}� �b� ��;YM�J8���j��\=�|�{���\��I�JS#h���;�89���8��_���֞Cd�	�m��ʀz��[��y� �|�\ݔ�4�IH���������o�i�՞�fE �7#lI7\ ��^<�`�U}V���P=�
����nή��m_��}T��g�w�u`�p�,��D�DܑX{��d��HN�O�3�rA0H$�X R �"BB(\W��VHb V���w��z)P*�C+,��$���O��)5�$$�Ga�_U|�=uR[�/�1p?UR[��v�j1�q��H��ۮ�w���w��{�BO�T �v�'�U���d��A�T^��웶X�{Y
�e�L��D�S�q�����;�ps%~����p{4jҔ��%E"����d���z�����Sf�k���D'M�`n�� 31���b�w\Y�.��bI���}�U�y�9�u;��1���F9��#�r�n��Âv�n'm�����\��Ps$�@
��b-�d�I#%B
qc3�e8�3^���x��g�#����|^~ܖ����n�ps%@َz������I�q* H�v{���꤃w\�{��;�8Ur���8�n�u`���1Xw���J�j�;YM�J8����}=�`�ps%@<���5iF@m��X{��d�$����'=�<��Q��YD�O!�{�T�@S��*�M�T^��Č      ��H��7R�k1Ӥ9��wO2b���GFX�N�� ��u��9�z�p�]v�5z��lO&h;&�v��Z��LuA�\=f;����wi�Y�o[s�n��e�j�	�;by�g�d�'3�fݬ���;�.�2ne��UM9�`+�� EU
�,ZC��)$�Hc$�#��A�f�U�G]u �f��ݺ�%��t뇕{���*k1B%�b�������8�ǭ�j1$�Y��E=_}Iך�3�\�J��g��S֣q8�mX��V��r�K�遫1@5w�hb ~�UT�g� ��J�~Y�����\�3U��:�&��T@��ݠ�vU��}�k��y� �|�YՃ�����+�5�ԻT;i!�u����ܵ��n�n���Ԏ�[����@w��܂uuP�Pp'	=ך�� 
ֶ�����rݫsM��TSļ�T�����6�2���/�)����/-� ��;�^6�dd��촹ݕ%Ř�ך݀w��ޓJ��$��V�z���5t�s<�'��!'�(t<8�a}$��ݦ+v-��]���e��z|ya�r3=�1̒ÉF� ��XPw��̔�Y��}:�<iSp������5OU
��6w=+��K�P����%��j܍�����I����1C���4IP�@ ȑ`HBH@�e�bT��J��+�y�U��}��]$��p�hX����FČp��~~��A�{j�;�8���\��@<�����*Rd�E`s�5X��g����D��^ȕm3cRI$�PuX8�S���턑����k�=+`�AY .���e`��� �2W�Z-� �j�;���):m��م�W�W�6�p�{�`�� �a��P���$�Xy/{���Z�ڶ��8se@��
�5��n���aԩw\&6W;0��jz"Ex������|�6I<�YMb�mGus<�$������5{[�_��V�>´�\&�Jq6k/P�NC�D�t{j�T�.���3\�`Їkjd|��P�����^�����8!�4F�D�A�I�� W�6o�|�<����9ݕ ��v��P�I�$v5�ă3\��P�� ��<IAl�����$��{{�֟�?.���`n�i�C�)Jm����ؗkvۻo�n,�y�&�x ����-2	l��Wk0    UV����IKi�9�n8lx�K�(�L����T����j���á.�r�[-��Il�ڲ���t79�g-���&��6�]ZqoA�:�^;vum��3�o,@�;q\Ws��')o�v�:m�N�7X�����w��������g���4��I�%��G<��{�V�23[qN{Y��K�^���P�&E`Q��]s%@:��E�F�q��'��W>�����}�8I���W�P��)�j����%A�x�T�}�`mc�#SJ��F�w�W˹�-� ���\$�ߜ$�/m �J1���[�D͙����̕ �do���UV,,��\nl��ɕ5�Ùc\���u�������w��I�%@��ߕ�gu�/�*ո����IJ�l���3��eUWP�� @@f�$�{T�y�.w�}U!<5_�P��JQ��-,�Ҡ������}� �a��P�Q���Y�����U}?K����+)/�* ^��1d#�DFՁ�y����P� [�ϑ��rI%8�N�i�bv�w[��������:����3]�-��8��ʣ��yo� �d�W�U �}�`mc�#SJ��AȬwe@:��������瀞5V���t�II*��s�M�fq����s�C����jxVQ��� �7Z�� �#a-K,"���Q��H���"�i� J@$a0�q�\U3�tqT�C���B\��t����R���ьa ��,��9�P;�	�	��F�#�i�/1��# �������h����!�K�����%3%%�4-eԅ1��1 m�鄸��0�JK�b�A��ˇ�v���ы7f�w5%"1����
"�E�: ^��Q:��� 2.��E:A; Cj'�({�u 9w��{�1@/�*��v���I�%��<�}HŚ��ʁꥏu@��f�q%*�TN+Vy@/�*��P��>�_��������O;��[R��������u�!n�ʦIL�T�48�J1��(����qgT����j�(�M�R��ccI��1{T��}T��y������4���	�!r"6���V.�_2T�q@5c)c�A�V+�	<�A	Ս�Ұ+�
�\�^ڰ=^~���%(��X�ʀuf(��+���0��RI$�	U.���z��1(%��.
�m�-����(z�MI*��z@/q]�b��h;�*��em1�R�$,y��`b��ׄ��5i)Pm��qZH��P
�d�{�K<�s�5X�*�Ԥ�%(�Շ��w=u �ɥ��<�`j�(s��r�⍍&��,٤¨C3x�t��g�$�$�)�3B�J	�
H�K�g��n��a�m"�d�G]��      h��݋N���0���ю�i����k��Q�l<=M���x��r=vL��{6�W�&��\&�;Y�����m�A���zt8L��8�֨۸��<�!���q��:�K�y����i�6ܙ��;j��ct.��ٺ������Eʆ��KrI#1�8�A��H��vn�I��Ѥ���t��i9m	��G$�Q�����h9ݕ����A������R�D�j8�]��̕ � ����G�^��Ҥ�r+��P���za`b�ew*6�II*��z@9̘X���nʀZ�;YLqT���٥�����*�x@k�W��'N�I$���|���nv6�=��`x���Ӫ�1&��JD��6�Q8���_2T�x{ꯪ�s�7 �үz�&J�ܙ��RN��6Ώ�#��@�h�����e��w��.%���Σ-��64��5� �y��cz����P��hLYR9$B���=�`qwT��P�� Y�KD�RE`b�j_�����Ձ�z@/�1X�1!�����I%�jP�9�ש�m@v�d�*LeN�m��.̓BG4~v߽zD$�<2�=���ug�$�3j6�H�qԒ�-�<��{��ŞS�#��P˨��c��&J$V<�U���P���뵞�P.�_;�ݤ�A�J�E`uw��d��� �y���4�v�7R�(�Ձ��,� �y������VVh7$�:\��p�G�c�*,��,cm�i�՞�f�57a�cI�������+��J �2T ��Bbʑ�"Q�`s^�HŚ��ʀb�PVj�b1�D��$VWu@s@5f(��Vּ5�BR����}�,�]@5n(�����K�A	�D$R�6|���翼��v��(�RAGRJv���P�ٺ�/j�_2TԺ�Zy$�q�n�^�:���8��wi�	��X��=s�huڏ���`un(9��UUV���s٣V���*)���Ps%@"���湊�_$nlI��N�"��ަ{ꯩ+�L,?,�(n�m��64����� �Ʌ���Ps%@�Z5�n9"M�ݚXN�<��6I=���$�+"�##	0'@,K$��� ���{۸���ߝ���U@S��ְک8�Y`      I�+,ֹ�(��/0灜5ˡ��^�1�m����*<�������y�N�g�'x��f\���$Xm&�NŒ"L�w]D��<c�ܺ��k�;T��;pÎ�G�Fc�T���Nj���*��e���Y.��u�<�
�v���s���Y�4 r[���f<<�탘��C�����Vp�<�PӴj܆�|��* {1���ܺ�6�����JTP��R��[h�p��u`s�Hq�+2�b� ���`�ps2��~���Z�wޕ ��v�����#����կwӕ`j�(�˫ �c�_{��J2�2IVWu@/2T �� �7.�UԫĤ��KK��J�L�,�'U����gZ��S����G98�V7eB��� �7.���s���
�lbn�w\���}�y�k꯳��u`qf��J���И�D�F۰9�۫����.nʀ�p�u��a"i�*�2g���;� �� �=�����D�*i%**r+��J�5����{-�WuM��{����Ʌ��6.��]�F����.�L++/r�$�7N��9J:�U�n�w��Vy,Y� �����c!ԢE`g}�VWu@3�*�1O��W��y6�H�dd��Y� �d�d�tV
���Rb@���E�'��!1���
��~J�!�?t�U��_ߔ�~˫ٱ-��8�V��u ���E�nr�ĺ�j�;���(n���X�T��;����̕m���&������'q�k�w�c�����8��vX�	�*�qH�mX�۫���̕ ՘����c�M�Vj�O� 6v�I]�	7�gG���H�����;se@1f(y,���Ky@���R�U��9VB�P�2�������ܯ�+g���@8�#Ք�B d�E`g}�u`uwT9��E�M�`~ؕz��ԒI$��j��m7�K�N��ΰr�'v���\4-
�]$��ZX��_2T�1x�3�۫�藠���Ձ��뫴�[����X]򟱳�m��li7Wi^�g{�VW|�H�d�{օCx��6Շ��{ݫV�@3�*�1@7c�M�VWu@3�*z���ݺ��ª�U}W~����!$c�\fi*Hϵp��xH��	!75�D	r�|�,F$D� ��4f�%��%i@]�!
K5���8Č�#;b�� F�;IG���,�&���G	It�%I�u��p���D��$�X����GTXB�%�5�#wxN�d�e-�ČaI�T@4 ����Yf�x���i)$���h  l�  �      [@�    �\���[���ٗ��  h                                 $ݲ�s' ��9i3fk1�<!�]poeۈ*�k��	�#�0�m��FP�|W��^{n�Z�����%��a�����"ʔ�[;vs�n�������i�%��7[1	VM����.�^�>��cv#[=���3��n�n[������M=m�I�	�v�^�yî�^��N�DnŜ���f����M�ju��!�2âm���v{l)�fn!��#l]�5h���\4��g��&��F<�{���5 ��I2��3�a��x�3�p����_1,���i�I�q2zkΖn�/h$�%�8]h�u�N�Z�Ň��U�����v���H��v��+����]8\��]�����rt;�ݞ�s��q�.y����Utm�s�ean-�WY���� ՙ�\Dh�j^��n�#��U��/qf���:���u��G.[�ØM�nz�9��K���U�&{[+���ós<[[�H�ݸ�N�J�mS�}�� �Z�Izk��	Jۥ��:�x �4�]*��gΌAag�۱ӣ��n�	"��[C�u�B
 �s��UUO.�K';Hm�vxMg�w<����u��تu��Uj(N6�k�fZ�kN�z���q<ٷ�Cu�<Gv�.]��;��l7"Ħ�����y�y�[y��υ삽���q=TL���N����ҝy�S�����y�����iV�X%�m��#��k0     �9zc�t�&��F�vL�@��;����l�g6�D��9� wk4�A�����w,�;[���<��;h���..w;b��r�b���r��{gV�pڧvP�s��u��6�Q��:��sa�&a�r���$��ܛ�e�r��S�{z�o�~SU]NM��o82[	�ܞڱ�.���#6��"*��"����PY��{.��� ŞS�˦�&�**nU�庠�eՁ:�����T��H9�+i��FE(�Yin{�V,� �d��� �wS�q6�#$��+����ʀj�P�r���ؖ�%%TBj���,� �7.���{�YS��UUtY�jŲ�Í�l�ݙ1���uN��3�P�#cI��E��(_39V|��փ��� ��Шoȑ8$�Vw��9=�o(�B�J����o�}UD:��(^zTb�H8<lU��$M6�X]��,�%�"�w��VwiF$j��**r+(9�*�1BO{���~�KyBO�

��eAʉ�W ��� �3.���@/2Ty�`S�)$�H(�j7#J�T������a�77>&�J�m��>(\J�H�{�~��b�)9�*��P�|���p���J�$u=P�@5f)9�˫w"[D�(�Q	��v��ŝP���G����A�<�{ι�m�7Ȧ���r�p��MՇꪪ^~�w��VUw���\ݺ��hT7��H�n,��7�x��*��ᆈh��h�7b�h�%�b~�}�{�dK��������W3��4�����K��$Cf�/E+k�͝K)�m��.fi�wı,O�ﮧ"X�%�׾���Kı?g���Q2%�by�=��uı,N�>�K~��M6��/��%�bw��59��r&D�>Ͼ���bX�'�~����Kı<�?]ND�,K�w=�����6��8�D�,K���Ȗ%�bw߾�q:�c� HdL��{��r%�bX���L��bX���x~�"C��TYh��}�%�޺�8�4X�%��}��r%�bX���ND�,�!�t v/�%���K�>R�h#A���ě�F`���D�,K�����Kİ�*r�y�f�q,K���yu9ı,N�{�<��A�F��$�lzI$�B�I��dc��0���{&��s��K�r�ήl�F��k�\�N�X�%��p��Kı=�}���bX�'_{�g��&D�*dL��J4��ho�uƓ�FYM�P�%�bX��ﮧ"X�%�׾����w"X�&g�]ND�,K��xjr%�bX�ϼ�)3=�v�ۙ���Kı;��}8�D�,K���Ȗ%�bw߼59ı,O��n�"X��F���6P��2&Z��Mh"x�"y�}u9��*dO}���"X�%��{���K���L��Ϻ�q:�bX�'����%��.M�n�'Q,K���xjr%�bX~����]O"Y�2&D�ߟtq:�bX�'������bX�'>���ƽ瓹}��wM݉i�H�ƺ)�v�     .�(%k *3X��\�a����v�#l�O�g�7=u��];Zݷ`�V�g��P���{]�P+/;;+���lq�^v��=���m�;T�����8)�ì���Z+M�����a�׺�m��۞K��9��j��/���w�U :�ԙ!�$�H�6�(=8>:�R�Zs���@��Y6���<��\Y����~7���x�;�~���bX�'���G��%�by�~�9"X�'}��S�,K��e;<>�.�ܓt����Kı>��}8�Cc�2%��y���Kı:����bX�'��S�?���0�F�����I8�fB�<��A�E=�]ND�,K���Ȗ%�b~�}���bX�'���g��%�b}�<^&0\M@�%7�4��hfo6A�Kı=�}���bX�'���r�:�bX�؞�߮�"X�%�����Y�nl��%�8�D�,K���Ȗ%�ٔ�¾��vq;�bX�'���S�,K��8jr%�bX��&�����j��dc' v�v�Kcv�e	����+��cE�Q�"M��"���h{=�Q�Kı<�>���bX�'}��S�,K��>�yu9ı7*gS�3%=3nݙ2��'Q,K��<��r�C��L ©.F��C6�-p��	T�U��P�l�X`���<�q#D�R��M�� "��O"X��y�S�,K��;��r%�bX���=�N��eL�by�?s%��&M�n�'Q,K��߸jr%�bX���ND��
ș����q:�bX�'���Ȗ%�bW�g���˳4ۓ4�uı,O���S�,K���y��u��*dL�>���bX�'}��S�,KĽ�I��.�ۤݼN�X�%���s�����ı=�~���bX�'�{�S�,K��=��r%�bX��y9�{�UU���Ӭ��s��l��x�uS��V6p�E8�f@[��t�֨3AȖ%�bwߜ59ĳ����z��,K��s���%�bX���9~�p��i�\�N�X�%�����Kı=�}���bX�'���g����,O��f�"~ʙ���l��ܹ�n��\É�Kı?g�]ND�,K��糉�K��Š@�E�b�
��è�D���59ı,O<���DȖ%�{�ܲ�=ݹ�r�̼N�X�~U`dO�~����%�b~�~���bX�'}��S��dK������Kı;s��fJzfݻ2e��uı,O��f�"X�%��~p��Kı>�<���bYA���Mh#A7R-�d����ػ9����*[f1�O+,��C��ec���;=��fl�;�bX�'���S�,K��<��r%�bX���޸�T��Ȗ%����jr%�bX�����.dٺmɚq:�bX�'��۩�@?(W �Ѽ�t�1���n�6��/|J)��*�F�уGĵ���r�Mi"X����\N�X�%������Kı;����bX�'_o�S�,K���%��˛���K���%�bX�y��Ȗ%�bwߜ59ı,N��&�"X�����C'-f�P頍h#C٧�����Y8�D�,K�=�Ȗ%�a����[5:�bX�'�>�Ӊ�Kı?y�2�h#A���}�I$`��x��s�±����۫��ٚ:]/W�_���|ȰNp�i�Kı=���ND�,K��糉�Kı?y�MylL�bX�{�]��A�F��֊%�m�	��D�,K�>�Ӊ�K�ّ>�MND�,K���@�&D�,N�|���h#AY��Bf�e�(t��bX���MND�,K���Ȗ?�dL����jr%�bX����N'Q,K����2[>��]2ٛ8�D�,�@Ȟ��F�"X�%������Kı?w�=�N�X�%�'�7�Ȗ%�bW�a�.dٺmɚq:�bX�'o�S�,K���y��uı,O�ߦ�"X�%��~p��K�7��_������W�SAi�]��    ���
��m��'g��'Jr���9h(�v����o`�A�nt���v�n�s�^��vg�c[q����v��{c�tau�3ֺ���g�*l�2\��b�����_{�Y#8�V�ge������%��k�'�]h9����}��{w��	����N�y5g[��jxǘ]�.�N��v�$իI��6t�ı,Lʟ�{����%�bX�y�MND�,K���Ȗ%�b;�P᠍h#C��.y䑘�nN'Q,K����jr%�bX���ND�,K���u9�ı>��{8�D���b}ﳗ�7	�f��rq:�bX�'�zp��Kı:�|���c�dL��~����%�bX�{��ND�,K�w̞�n\ɷl%É�Kı;�}���bX�'���g��dK����jr%�bX�y�NA�,K���m��wn��K�8�D�,K�>�Ӊ�Kİ~�~���bX�'}��S�,K����jr%�bX�����ٓw��UW%��3aݰs]@�$�Ω\cD�f&҅�b���=�f�4������Kı;����bX�'_o�C��L�bX�߼�q:�bX�'�s%��L&�l͜N�X�%�����1���ȁ5�*	, 0.q@�OEPǸ��b{����Kı<��{8�D�,K�7�ȟ�L*dK��>���s&��s3N'Q,K����59ı,O{���'Q,K����59ϠdL�����Jh#A�J8�eF\<��A�0��k��E�v�h��h�+��f��bX�w�ND�,K�����K�hw0�����Fd�yC��4-�ș��59���L��H��]�D�,K�����Kı?w�=�N�kT��P���?�RI$��Ev���k�[���Ү�bs�u��Eh�-�.�'����bX�'~��S�,K����jr%�bX�������ı;�~���bX�'������nܥ�q:�bX�'�o�S��9"X�y�>���%�bX�g��ND�,K�<�ȟ�ʙľ���[�����K�8�D�,K����q:�bX�'y��g���!���{�"tʭa_c�D"  ��h��.0�	͹�,c(D��f.4�3@�B1@��XV�Iy��dH���#	�H�H�`�`A�C	�!Q�p������Na@@��ȟ2p_oxe�i���z����<N 9�h '�'�(w؊oi��:j�
����բ��x��'j�)E`�Qλ�ϻC�B��؞f�MND�,K���Ȗ%�b^��̶�mٷfL����K�yCbo�����bX�'���S�,K����jr%�`~�.Ǩo�w��wı,O��[��l��s&�q:�bX�'�{�S�,K����jr%�bX�w�=��DȖ%��|��F�4.�b���M�$�&���6��l������͉����kUQ��؉�sN'Q,K9"y�>���bX�'�y�g��%�b^��59ı,N��"X�%�z;<>�73nY��6q:�bX�'�}ϧ��%�b^��59ı,N��"X�%������B"��������F`������b^��59ı,O;�"X���<�y59ı,O����'Q,K���g/�]�v�4�3��Kʙ"y�59ı,O=�&�"X�%��5m;"��R�,7z��+%R�+[��9ı,N��l��[�Mٔ�'Q,K��>��r%�bX~P��}�Ӊ�K!�2%�f�"X�%��~p�p�F�4����%���I$0�R'7��9��n�����;���"�>�~7��Dȟy�>�N�X�%�}����Kı;��9"X�'��S�,KĽϯ�m=�fܙ2��'Q,Kľy�jr�9 {2'��ND�,K�}���Kı?w�=�N�X�%�����I�e.��7s��Kı<����bX�'�{���Kı>��{8�D�,K��٩Ȗ%�bS�߳�.d�7M��8�D�,K���Ȗ%�b{߼�q:�bX�%�ϳS�,K��8jr%�bX����q0�E�4��h{=�'Q,Kľy�jr%�bX���ND�,K��۩Ȗ%�by�/0D^�"5XR��!*԰PB�!Cw�7�6�IH���ؑ���`��v��      �޳\��������m��Yy�Nrӫ��,���B�lC��Yc���v�wY�17.K�7>^�Ƌ;$Ml��c8��^]���Z㝀��[]�wG$cu�mɽѯDuuF��K�k����I��%�z���1�3r�6̟x�</\;��!��*��X]����K�¼e�tdܚk�ݬ�N�I����p��;O�X�%�|��59ı,N��"X�%��{���KĻS������%�bX�y���Ji�n�[���%�bX�y�NBFı,Os�n�"X�%��~����%�bX��>�ND�,K����{na7fR�8�D�,K�}���bX�'���g��%�b_'�]ND�,K�9�p�F�4���AjqĚI���D�,�=�Ӊ�Kı/�}���bX�'}��S�,K��=��r%�bX����-��vmɓ.��uı,K�f�"X�%��~p��Kİ�3=��r%�bXr?w�^�'q�F�46��>�&�A#-�.]�B )ҝ���DNâ��+6y �)�e����oq��K�=�Ȗ%�b{��u9ı,O�����D�L�bX��f�"^Tș��>�is%ٺnfi��%�bX��Ϯ�!���� @� �D#�9ߋ�)���T�{���'��%�b_<�59ı,N��D����;"_=?I��7	�f��uı,O�~����%�bX��>�ND�,K���Ȗ%�b}��v�h#D�h.��rH̀�(v%�g�X�=��jr%�bX}}��S��%�b~Ͼ���bX�D�Ͼ��uı,O?}�uM)�ͺin���%�z���juı,N��n�"X�%��~����%�bX��>�N�F�44h�Kd�I �S���\�=b��m^be<��a���9�����'�{��bX�'���S�,K���}��uı,K�f��	�N��D�<�xjr%�bX����i~�we�nf^'Q,K����tq:���L�b_}����bX�'�{�S�,K����u9�r�D�/s��-��lۓ&\Ӊ�Kı�g���N�X�%��~p��Kz��B�}uq4.��yș�~���bX�'�{�G��%�bw����}�R��ɹ�N�Y�2~U�~���Kı>Ͻ���ca"X���ގ'Q,K��?o�]ND�,K��>�is%ٺnfi��%�bX���n�"X6%��~����%�bX�g��ND�,K���Ȗ%���{��?��ߓ��UU��vƔ�k�b}����$(���ָ�9뭙t�\���~w���%�!��߻8�ı,K���Ȗ%��ȗ�8h~@�L�bX���n�h#A
�J_r3.A�	�b_*dO۾�NC�r&D�<����bX�'��۩Ȗ%�b~��z8�{S�,Oߺ����6��7fe�uı,O}���"X�%��y���Kı?w�N�X�%�|����Kı=��g��ve-É�Kı>�~���bX�'���G��%�g�2��jr%�`th$$��A���z���ѩȖ%�b_g~�K=36L�m̜N�X�%���}���%�bX��ϳS�,K��8jr%�c�2'�s�Ȗ%�v���z���l�U��yKRɋ��o�o��t|o���r�26����e�ݙ72d˚v�ı,K���59ı,N��"X�%���}���L�bX����'Q,K������~̲nm̛���%�bX�y�ND�,K�w٩Ȗ%�b}߾�q:�bX�%�ϳS�,KħS�}�L�vn���q:�bX�'�o�S�,K���}��gU2%�b_<�59ı,N�pJ4��h.�<K���PH���%�b}��tq:�bX�%�ϳS�,K��8jr%�`~BdG�猡�A�F��җ������uı,K石S�,K���糣S��%�g�;��59ı,O��z9C��4���<�r!�&�6���Č      ����7�f0�u:7�8�j笹��N*𔜝r3���	����׬xw[^3����(�E�2ڭϤd0㚺�:q�d���+�u61��9��u틡��[ݘ%^8�u��\=��[���6�t�۹qܹ�TO8�u7߀y着�����C��r�ƶ8����s��C�9l�6ilˤ�M�t��ΓȖ%�b{��59ı,O}�f�"X�%���}��uc�2%�}����Kı/K�[�Mٔ�'Q,K����jr%�b]��~����%�bX��>�ND�,K���Ȗ%�by�ym,��3L�n���uı,O���'Q,Or�D�����K��2'{�ND�,K�v�u9ı,O3���-����2e�8�D�,�D�����Kı;���S�,r"}��59ı,O��ގ'Q,K�����I�e76�M��uı,O<���"X�%�����Kı>��z8�D�,K��r�h#Agq&H{
�I$�K����U!e+�݆�h`n��v�l읲��qj���8�D�,K���٩�KĭֵrȻD4CD4Fs���	�4S��=�Ȗ%�b^�O�f�m�sMܜN�X�%���~��u%: }7��E0��DȖ'���ND�,K�>�Ȗ%�b{��59�TȖ%��e���wv��.���%�bX����<�bX�'���S�,~D�Dȟ�ߦ�NDȖ%ʟ����'q,K���ӗ�i�r��q:�bY����jr%�bX�g��ND�,K�|����Kı<��jr%�bX��v_s�s	�2����%�bX�g�]ND�,K�|���N�X�%��sS�,K��8jr%�bX��a$�߿��UN�<6�ɏm{td���(Wk��!��� n�e�2�s2��ı,K�>����Kı<��jr%�bX���	�Eh-�B@�C��$q��ON	#�[�>�؟D�,O����"X�%��{���Kı<��z8�D�,K���-'ٔ�ۆ��uı,O����"X6%��{���K9���  F0b�"F�`H!	! � ���G��ȞD�:���;��,Ko��q�f�4���l�d����%�b}�}u9ı,O;�ގ'Q,Kľy�jr%�`~A&D{=�(p�F�4��`��.7��N�X�%���uı,K�f�"X�%��~���Kı>�}���F�4>�O5&��I!���@���g���\=ly��O��U"˖�,i�\�����,K�����Kı<����bX�'��۩Ȗ%�by��59ı,O��r�M�6��Kw8�D�,K�>��~�DȖ'���S�,K����59Ľ�ș���ND�,K����~�0��)nN�X�%��}���Kı<�}����石d�v~� ��Ԓ(�r�I6Ձ�z@s�;��6L�A{�$RC�U�����V�֡'���cIh�c6W(y������~Y�CGJ��]����n!-�ۧ����ҝ����F���6�8�8� ���,� �.j�@R;�R�7P��nU��u@;�5@;͕ .�]���r�F�[���P�eMHK1@�D���Rm����?TO(�@����꯺�~�~�z��&�D(��ʀ<y���ި5@7��晴�>�{���Y@�����`,XD��$���a83@��HXc)0��ˡ�i��R D�ŀ@�) BM3BV�sH����`B1�c!Ir%�B$! D\c6jD"B0�� �xdb�B�0g+	!Bk�\!$�8�K��
K���$I�Ϙ���"B$��aYx�8l\ч]S.k)CL2\�Ws$����0B2!"*͝u�:���BPUP���QܥJ�I$�T�I"�  �:  �lm��  @  [@�$   �ܒ�����d�'Z 8 p[@                                l�]ض�]#��.��LrTc˺�5���չ�lVЃ/<1�G;v�f\M����ͩ���ݧ�:}9��G\p��nonPƣ)"�=FM�q��wm�c+
�N9;�
�n�+24q��}�v}X�ln
��.%7nO1��h��tCI�Q�;��r��Ǭc�`�8�Ai0nLm��Rdy++U���h��ֳ�p�5�#�J����I�7m{<�s^�l�0j(1�ݙs��5m��F.�m4=>����)�"��[�h�S�ۮ�Y�û}�e�g�qh8w�F��T،[C�ӓ7Ynݝ���UV1�U�1�Z�'"m�V���u��.��wm�m7c�O+��nv��d
�,X�v㠮6��zSg�-�y9���;��\�cc�����=�F�Nn�r$tE�t���D��r�>:��wf���<�z��W�s��}ͮ8�ζHq�n�'0�܈X.�e��vmZ��.zI(v;vr������EvY�g�V��+�Iġ�di;=�j�e�.۞�G2�k��'Vt����n(�Yy4=��]�ۚ[�Me\��o5U*Ơ�zq��++<�e��j��M��36��oY�<vBr��V��ˣ��*1.�K۝�۞�m�N�c��u�����w������b�t�S�M�8��ﺯڔ���`/@���D��
�N�z�OLG�_*�������$�,�y��$H�JFd�dq�Jtu�X�     �Cڢ�$�d�g�������Lv�f�:�Z'�?O�}�C���o �Z��un�T&9Ϋv�m�4��giNUuŵ���;k���^���b��[������9������a·-����m��Unݼ��ѭc,2nSM7f�8��~ ����
�����*�q�m �(�m�	 ��i�Ժ;T�2�(�'%%�'Z(Vf;���;�P��I����j�[���P�j���?�H���ZM���&�Y� �2T�1@:���1*1�Q��Ƭ�ʀb3kqBA���GK�Q����pp��� ��P.j�w�*��tx�-UfMٶK���8@�y�֖2;��f�箲I���V-� ��(y��U����S��N@M����)*~��P����Ř�&ױO���	�LCI�"�TB�����փV�b�� s�p.!v��n��'Vn�T�-BI�u�~����$��$���$$�VD�{T �q�;͕ ՘������7~�UUr[����4w<�����e�^��r	C"�$�jH:���w<�igvT�:�^� ���J�mTq6F�^�	8�$��P�{�s�RG�);�(�MB؍�:Iߟ�BM���JX6"eR 0�	T�
@�����U������ uDUUNa������N�b���\L��t�V-� 9�p�e@T��(}����QX{���}�۫�u@:���\J��%$�I+`��ļ�Og���\�E�ӟImm�����J�M�%�fʀb�c���z@� ��Rn���'V�� ��� �6T(;Kz�Eb�$$�Vk� s���ʀj�P����mIB�`�y�����꯾���s�������O>;ܖ���Q�ؠ��@1f(w%@s\6�߾���Ʌ���-��ϱ�W���q��1���n�*⎓j	�mʰ�p�J�O{��u���!$���L�ĄFd|=��9��l�����l�� '&�*�3?8y���UUI�p�ʀ{�E��T���3�� 31����P�� /��ԛ��"��X��v��;�8y�P�������/��jy^�&����X      �k��j��u��uI#XJln�גy�� o)�M�Ol8;�k��:�;6�Q�:�^�\6�e6�M��6[�n@N�%��G����Z��$60jv�	�,�[��R��ɤ�ζ�]v��iFݒ����O�.5'��� 
�t��I$�pRx�l�l��\Ȏ�W��L�v�#"�kWM��R+�$��$�~��T*��>In�.�Z�N6���J���s��J���̕ ��ͥ�Q���3�* fc�wrT �5�
���&��ەaķu�3vT �1�𪠻�����<d�r3#�&���qz��o��g�@f8���3P�m�,���&y5�ٺ�3�Zn�����ۤ��%X{�}�Ps�k=$�4�4FbQ�Q�y�&��
�6$$,��Y�s}�6�nśo���<I�JB$'W�$��s�*����;�8sҠ^�#NJ�m�j���ʰ�8q%�Ҡj_�\������� �)V���?}U��o�p�\���s��ԭ$ܒIR1�wMq��S����m�q1;��Y��������m�͕ 31�9]�P�� �:�R�mA:��\ ��s�* s���ʀ��i%7c��;w6��;�r�uDH)AHB�_�pP��[�'%f��$�R�DN2SqJ�w���P���ʀop�`�ģ���&�`���P��o=* s�n#��z��үI$�J��Gqp�n{il�����㇥�S��)b`,h0� ;�p9��p���W��;a���/h#"�؛m��J��8;���8�%�$�jH�R�$;��d�����zT���J���H�#v�ﾥ��� n�q|𖔜��B�  hfgϼD�!�~Q�\I���V��DǄ �k����T�{������߃��UU��x�BN�FW�;dx�;HZ���Д�D�T$�"Q�FH��~ 9��zW���\ �pK�Q�	���;�8y���8u� ��eFD��)(��ʀ��ׄ �5��4��Z��HN���w���Y�]@1{)���|妯��/���̌�򪀧b��ζ�X�I�m�Z�iKk�Z0     �9fgV���hiY7=��Y]9Ȧ핥�N9�tK"rj��Gl��P�7�U����)��^��q��y�rf��C�3�J�����63�5t�Ù;l�k��R'B޵%��:vM;q6e������3��rj��yK+���"h�]�3�37wwL�s&e�5�.y�n��nۣ}�֎��b�8FS�Q"Q�'�˴+e����Yz��̂�a���XȒ&�|z��!����ڪ��O�
6F%*$�n{�8,�!�.�_�΋0@�1�#2p,^�W���`^�J�l���M&�QV]�����݁����t�Ԙcd���ig�m�a��pqs��]λ\L�V��=��t�B�S�qۻ��mU��*�Ie)&�.?O~��$��`��'�׾w����E�1�$e��l�;����/���̃�m,l��m������A���dwM���D�6c�z��fAgqU��*��-�$�H�&�1z�nd�ά�`���3�)��Ģb�:��U����W���~`gl`�'e�̜}����7-0/o%s�R�A�"S�EY���eQ�N��n�z� bb�Lr�2�
�ː���J�A������BRcFN$�
a`�$.(F�
c.)��,b%W`�.H�H2�*���n�01b��H���!@�!�1aG
K�0�	q��\%0P&9pJ1��L����*@�B�(J�)$�
0�(��E`�22ʖ�0���F�"A�Ff�q:�$0&�n��3#\.�:3H������p`p�,S�\&a%�A�:`F����B�+���Ȥ�p�#��F4JIJc�d���L2t@!�g���u��9Ĝ�ˁ�+h�@j���l%��bd�A�nz�;s���I��È��'B�!�� N)�{抁����*��H +j��.w�t�ol��c0�!`�82��yy��W�쫲�=��1"�iջ��W���`r�$���-U:D ��9�7[v�jZ��B���
�y�a��"H�e6���܂����:v���N7���^fo^���̂�ګ�m��D�6c����dw�˿A���c�Dʉ1r���ރ�uR�����Fb�����:�m����ّ@\1�#2pg���]�Y����������a7�j�E���m=���MۢvF��l���uR4�j4"0c���M�[��3���g�Wyi�^ZLf�(%9Ӌ���/V��g��`�%���$S}�@oE�� ��0�$e��o�5i��r��yN�X�I������`^�Az���Ί�"��}M�"Zd,1�Jz�j�� t>   \���������B�1Ǫk��R	dq�����c	�Uq�6���\�P��:�a��*��L����d��-�<v��r��E�X1�fԖ�m�sI�1`Z���ܶ�x�Wۅ�:۸�ۢ��F��\�7#~,1UC�K��GY��I'#%@Qw2���bqo�w���˰-��pܩ�'uB��w���0// ��a������L8B8��)�b&�Y�l��a�;�s��ӝ���@d�#2pf�5}�Nǰi��]��� �	)�ᬻ�/���̂�a��Xbj�%8?��f��yi��n �������t�<Eʼ��Q�([�m�܄���]����1!-%!���݂�a��w�~`^{	X�2�M����H�:�IS�B"J��浝�k�C�h������j")�Yw�_q��UTs۰g���{m�M��&_�i����Xj�ݕ�fޥ1��M�3w`�Xj�݂�u��Յ�E7$�!�������S��t��|J��9$lA"��#.Fd��/�� ���{�+���
���.˽��]�7�o57�qCqF�A)�����͝xFI �a A�� ���"�0���}�F���%�[��We�Ĕ���y��{<�k.�a�B�^��xH�đ��m���^˽��y�~̃�V�Dy�$�NŸ�k{\۸�.�uD�n{��U�"�jx[1Ƌr˽�����;��g}���zȎ&�|�~#�@�����x�]�<E�8�J&cE���o��1a��}�]�E�� ����f�5|�A}�Z:o@�I�Ab7��� ���[[�h�JBKp�k.��d^�A�XzFആȔ�I$*Q)H�h)at�u��Ŝ�ܖ��g�&(�1Cq(\%82��y������vU�����B�`f��x�����X��F$��Sm�^k�܃���Ɇ��Z�M�だc#�B��w`���2Wmx��q��/�ُ��X���^5}����
�����"��m"��C���      2���r8�x�5�
�j{N�6�fn�Β��pl�C���뗇 �K�;�nrM�tgfz	��kh�r�z\����I�!ڸ�h6��X�vn ���oh6y��;M��>]bx��𱑱�r�.�=�����@���\B̧����q{}��GY����*m:ɫ�Izq���&�`�zl�����n$cQ�َ8�~Pv���}�y�v�E�F\���x�j�ܐ���k��0~sx5�EHI���ng�v��}��x�kݲsE���‪�@3w`���һҬl%�������v���goX/	al�I$B�Rx�������oNSƥ���=�dL[Y�F\*�׋M_{�ް&�YN�X�M��R�w1�U(@Tcހ!�N�$sv���ߵ��/Y�ُ�7���f���vW:��F5-���(��/����v���tXؠ2��8,�� ]����=ԕ�2B��Ub�j��!]݊�p�b�g��ݧ�$�n���bY�F�U�/vp^ks2��[�'24�Q�Jp^kF,�:oU_{��Ҭl%��7e��}�N�~S��UR ��<�I$@�Z/�-��_��Q#M��g<���o]}B�={�bZ�M��r@�_b�z�=5����v�E��$ܒH$d�Ԇ8	��n����:���tݍ2��F�@��%��*p^y֝��,�#��+���F5-��nnA�x��ۃ���E��P9���j�w.ް6��s���Tn2dn5]��;x�����������sD��З��5�&
b�j`�1$$�Lˉ�Ԅ��Q`FR�@ݸ2ˢX�7����{����z�qF�AG���/.��\��w�������-�a_f牻N��vE'y���Z�ӹ�-�TZ��QL��:o�w�f�;y�q)����Ú����M��3<��eͪ��-L&�.D������`L˂���q��/��R�ЀַA��4a�pi ��i_��C�F�fI!ٹ�T��α���}ǻ�������z���m�6�@5 ��J�� ������("3� ��% �o$~�˩Uu
>��*i'����I�g]t�!ZY�̰��[a!&�`��HB܎�2% Q�)r"AE D r ��#H	�TX�QBA:�"�H��P�2"2"�H!E�	`�"�H(H## ��!"�������*�QldT$A$U$di,I ��QID�I	D$ Be,ABD�	 VE$$@RD�ARA�DP$d YB@EY� 2
�
����&�OIi(
; @EdQ�P��Ob U:��	"uj�"HȢH�DKd $@���!����	�٠&�ATDP@  l@@ S �T65T���D]������������4d�$���l)$#B;<�z��*��@�O����H��y@�_���?�(
�"��Ȉ��B!"}$�3����[�~��~��%҉g�V��O?�f��8�kYs��{<���^P��n�{`��h_�׷�/R���z �[AD���0W�2���c��t{9��
��$��-�?�E�~����������щh�x�H_�� I!�B I�aa1�m(�Q�w���(��ڏ��=G��/��(�%
������@�z�o�� ���7����]�B��?�BI	~=_�4��$����?Y�����?��41I��OE��c�iI>$Q�R%�i���W髠,�L";ɒ&�K��
�����Hj���j�kn���d �g���>Q�����p��>��Z�hl��_�4���c�������P���@�$�H(�)""�*�)"��H�,"�0��2�
2*���b�HF0��"H�F "��� ��	* �2�4�"�$�Z������� ! �H+ �"�H*H�Ȁ���H'�*Y"��B* F ��!	"���$"H�"�
� �H����"� ! ���"*)! �Ȉ3��  Ȣ1���F `��"� ��(	���,"��H�H H$"�� B)"��"	 0��B
�0����� � #"�"� 
�",��1,T	IFBH"( Ȩ{��/0��T�A��U>S�<��z���WTpϧ����B� ��_P�Gi K [#dTd�D#3���t� �>^�Ҽ����#�ak�IHz�ˋ�׶��Itx�w�7�gpw������H?O��f��S?����폪�r���� ���7@�HH�#�� �c���B���~h���5c�8���ɒ����c��@�.�{�E�#������i[B>���WvO5�2-���������3�L=����������z�z�z�K�|��瘐H�z;h`!�z��������O��χ��aveɸ;=�j�i3��d��`	 !4z�$��/�j�L��(�Q�����%��lI ��I�㲌!A���߄����+�`=�<]�i��Kl��{�7�	;^B�&Z��.2��e�3V1�"7� ���dE"��C�d#,
D?���J�KZJZ���dP����%/��h5�R�Ő�� �
J����_��+�k�Б(]���	$$؅��;���;�����W��c���M�!(��=���~��_��z:����=��M6���q���{�O�tx��^��&���]���O�H�V�g����4�j�hWE/�hHHw��W��=����� l_䔙	�Ϧ �a�	$$
~�`� G��'������]�#���;����h=]�0Q�����]����@`�{�_�؛�e%.ىI�	����z�D%~q�χ�{��#=�0/�e�PN��.��R��י�eI	Ҽ!~�W����D6�S��	�]���拇���b�O�ǧ���	�m4t�I �r�����O��B�xJ5��};�='��<<O��{��BH@���z�9G����.B������S��yZ^]� !�bHBB���-5ߐ�I �=��JG��"\{��a�k�Հ�0z��|=2C/�����e���2Q�w�H�?�.�p� � c<