BZh91AY&SY�1� �_�px���������`�}n ���-���  -�ޏY�p�tZ�hH���S�T�T�Q� =A�S@=@4II%P�     �A�ɓ&F�L�LS�)�L��j44i�  FA�A�S&Q�j�MA����4��$�BjbSm4���ML���� 4�NK����*�`D$Eu"H3��Q���	$h"0)i��jI%�`���q���QD@1��SZZZ�Ǣ�&�t�����d���&Iɒ(�Y$�B(�D$��E�	:(�B):!$�'EB(�d��D"IB��8��8���Ȳ(��I%ݼG<Y��x5�#����8����P#��__o��T'NfEN��Ww5��Cn-�od���0M�}��R�c4I�u�h�Aq"��|E�r ��G(��0f*T`��a"�j�:4��w5@5�t�اw�SR�	�����N/w �(dx$�3��Ʉl�	�efI�a&2d�d��[-��$�d�UݎG���@?��X���NN@e�_]xM:�t���
	�'e���6;r��F���y0V�YF[���s�E�2��"�q���2�IM�}?K��bi���w�_��AG^�hm�P2_j{S���XF~�߅����$�In����I$�I$�I$�I$�I$�I$�In����I$�I�I$�;�Bׁ�a���B{�8�!<��;�{hқjw�7{7��5d@�Hk�	��mME��{��[����R'��/����0� X�n�.��-`���w���4f�Ͱ�T�Sz�B�b ��13 ��$�����9Uc��y�}e|�����?ɋDk��O@��t弉rс��.UŌ��N�j�f��MM�٪���0*2e���R<+0��#h;�ễ��	��f6� X�T����Ly9O�x��p<Z�5�.�]���<�_e������nC�wn "7z�`KCi�W��4@��g�'"b`�B�fg��s����O�G%��x�8�S�G�4�8f��.��p�IP�Z�/y�Kic�f ˍ#ۜ�Ő��`��j>;*Ȳ�o0,�]�X	Ѧ����:�վ�J�I%ad$0r�L�$�a3ow��UP0�"^�ԩܿ_8�d0���Fmz��'L�l��T,�K Y�{"G�6<�{wf�V�㥄$%��b�lɒ��M��7�t��D;�wC�iv�M`��,���;0:C۹klЀ�Q'��|�|����P��߰�/�Z�ꌘ�sf���@�/'�>���t^hj+�e�����.s�:�wd��� t�\8��݁߳����ﵣ���~d+ߦ����AD"�{ɘQ��r�f�^kU�C6����B���50� fz4e�!ޠ�K��iU�l>��7��ǘ.ꋶW��6���#V�����t\��ȓk���]f���R�Jt�h�3�B��ay����`1�8{<Ng�»�v�Ï�U#H�ڣ�e��9��͎�9J�/5�n�C����%�|��˘�z��v��k�2���؉����YOQ����¸ǚv���8���#��� �W^����8���58s-�7�b�	1��u��;�B0)P��Ŏk��ou���l\?���!ޖ�g:��P.=�xQ�$�p���8���Y�8[�A�j(�WE^�wC�0�+|۟N�[������Q���e�:�`d�ϱj�$Y˷�s7�30� N4�+�Bz$g�m��tkƍ�8�o7ׇ�VٽR �������&�W;�_k����=[M��[ �w���+c;x<>�b���=��rj���jԺ�dN�6���6;��z�e��,���F@:ҋ��O����y���2kq��m�� �|�c�F�c�}\^�-�F��t�h�ou�WD�}0,�^o3����|�|5�U	v/�"	.���LH�F�Z�{g�4?�A��{/�Q�]���E�A�
��{7��%�<�|�^���q�i��H4A���*fW��d�=�~��G���2�?$&a���v\Z���;60��f
�(ߑ1�'ǫ+4>�m��Wo���4Ջ�M�/�8b�k��9ģ1g8A[o{e�(TƊthk�8]�e<A,�"��"vf>�����gy3�z�\\x�����̻�����C�KH�Kڪ��,F�:���2X���|;|��v/s"�[K{�h�)��X|�p�4ak��4�J�TH��������#
R"�����K���%EV�UUDITH��-��EF�P�MX�.PB��h`�$",b�b��e�TA�m�R@)�ԵD��Yb�$� �6��4�K����E(�%��������o��|h*q���DDdCTҍv���׫<|L򶾜�dLr�	�__�i���L�Qj8Tn��Q�\+g�X���Ẏ��ܪ���K��N���Й���}\i�؎�������E��BA�����u���iDv�9�	S�5���3I#�8�נ!
�@xn=�n���lC��#4KR����&_$�&��)�B�
N�Y�ssH�W�ǝa|[�(/p��7��k�bk���~I��&ɪH[@��)A�B4

���R�*��
�"�cZ�PTZZiUAJ��)���B�J��0��tf鸆d3���578H*��>�����D����j	QHEI�I���feӿ����s��k�0C�����L�,9 /�"����R�#��ds�`DDi�)3�����2v��_�s�lM�����ہ�Jm���bR��3	���6����X�%�}� Dt�<�h(k���>�e���2�O� ́�u �@�#�t�p`�a��C�wQq�;C�p���Ĉ�GdD[
f#Md�L���d�Z��7��s
�qa��j� "�-7 �%�a�CE���	�����P�MB��r&n�/^�	��w#�l,�?��e��������π�R�$yt��[ˡ�r��O�(��w���u\��U�F��0.1�#�v]Anz����ώ����lJC�;˦�QŐ!p!׹��QAK2��m8��LN�ukL�zǍ��v&N���զ ���M7�Jj<��`k P� s7'ǳQ�`��ؠ���ᕌ(1�+��q͐]����DE�a�*l�LDGJ��]���7=Q� �V�`.YktZ�"mTTʤM;1lޡ∶ ��̸���H�
�#0�