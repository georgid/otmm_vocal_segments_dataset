BZh91AY&SY��� e߀Py���������`����4���uT
U %PP� �
"(��+^�-�:w$.m]SUB*F� "����&�6���@PL5�OԀ244   ���b�LFCC �#QI2�!��4�F�  OP%�	�Ѥh���~���h�P��6���	D����2&���� 2����}��5�Ds y�D��~���+T��
�&A��q����< ����Na�Xhlqz'�������{�>�����l�}�Cl�"�9�q�g��N%P'���	)�8���N'��%,�I$�����`��]��N'�R���JD���N'�N%P�Ĕ�)��J�q8�R�$�I.�N�:�~���P�:q:JD�Bt�ӥP�(I.	҄�:u��5���6�5��}�5�#4�>h��{��|~%̢�Ƿ��=K(���n�e�YfO��b�c�ZΙd4`��Q�&b��$rK"� �psh�\6���S�$�NI��I�r��n�w(�OU[y&��f�ɪ|tq�&��[V�N�a��ZN�M��_#F`6Q�a�̼�s1���'�^]D�,ݯr�a��B��t��u�"���$�vs�����qs����ū`�UY�Id0YE�Qc �0��e���1B�d,(����1�e�L��X�B1���]Pꮬc�ݻ�jֈ����ϛ�}'�����X�p�g}��Kjz�9{���%���c����X���X�<���
n4�� ӈӄ����eZ��2����TE]�2�XP[!P�gؽ�u��_� 44RqbG��M~0��DT��n����6��d��ڴ$S�jlN��
��K�KJ����!B�!B�!q�!B�!B�!B�!B�!Q�I$�I$�I$�@�"ᥒ�c�D6P�h��,��H8i9�ք��n�$����q��`ia@�>C`Ch�9%%E�p�5�zr��Go�z�P�R$�XH��;kF�vt��o���h ���h �)
ZhB�G��ge�ԕ$�{|>7nos<�!�dac�l��FR��a��Ʋ2�%8h��������,�$NF��q�rtm��6����c oe}����7TN��2o�l5�G.��fߺ �����s�?��&���$��s�]�o�{L��UW:���t�o3�#9+�2�f޹���~�XD�t��J�ih}1:rkH���� X;cn�v��,�<�F�4���ċ�+|O!�#.�7\o�v""�4�ӧ�{uIN��(8c@�;3�R�!R}�u���a��C;��8Ps&���Mv"C�C'Ñ�l}KFތ�jƅ��F �i�46dcγ��Yh�2΋+��X�<ؗ��a�ё�׿+f�d��A�F����,h<gpYȇ� 1������ ?F�Mc�8�R-DU�H#� �P�e��2Q���]���P��q��[XæH�5��fݐiV�fN�
K: �XAi�F��k�}f>�,�x?����>�����9��?:aChe�2cŦ͕�9�
:�6�$q�m�$�g<h�p�a<<���ɍ-�[����-��^��<�Xx5��6j%. +< �V3�Fa�Cֆ)qfh����q���Ip��lG���#,3۫.$C8m%Ӧ�
2!�04�3�B�xyAM��b7�K�j��@�l�f�44q��?;�A��u��z{[ɿ#t:�AXW��ġ����/>�0ؘ� ��&¬(r����|�tək��͐U��ܼiܫ��A��[x���x)�GmsJ!��q��.L�'���
�O�Hf�,h�S0>�e�*�1h�P��>��=�5�-�Y�3�_.��Cy��f�Eó}�d�MX�X�Gl~A,ɖT��p�S�9�:�j�4�gDQ�C���;\�"�i�(�<_���@�~<O(�(q��r��޷��w*��tTn�v ]6J��ُ3��`�8�H_}^����k*̈҃��h ��0��(�8L(29'	8Px�gL4�dxӥ�83��?c�<(4z�DZ�J�������?rc��#�᪉ /�V�g9���q�����$�=�$fq�@d<e����;�*��E4�3�LE4��̴Uې�u��(K�8;���6t�N�̮��d~x�v�]HQ���2q�.9��]J���$���Β"��⹉�|گg�dt���A�(�N9Cx��U�[�K�T�d�ųaFԕ�>NM�G�;	Á<+�%�k����)���7+�6Q�W�8ږ$u�(����u��t��4X�>h��{\���(��932�8m�*��byuq��>~����_h�C�vw�rj���Ȏ|�hh�!C)Q5!X�8Yc(gA'��:I��#E�e5�.�A8�H�$x����3C>�9��}E��������2���N_L�8E�P�i*��!��D6�G
晧~�_є���Ξ��j��J�,��a�B�:T��c[4G\O�����X����/��8bD��׼��\��>��4�,�\���ӝ(�F]�j��᎔#N��{�Q��$(y,��5`���q
iٸg�Yo"�)�g1x��p4���L�`��J�Հqя9&Yr[4Q��V��iݻ��漒L�X�/�����, ���
��h�rb�
!������7�>͡���&1h�����ï_/OY�T{nsܰp�42
��T7D(�������0��s8s���rB�}����l^I�.o1�|��*��Y�DS_b^v��'�u�����o�rI��1�-�l%!+@����sW�f܊)ۻ�Y�x�0��Xw�މ�Wpͺ����cb�A�qΟ[�3�s���-�
\��9����,�b;��TY�!ݗ���J��$�G
<.zy��)Y㙦l�,;�� �w 𫙆�kw��ӥ�<9��anOv��e/��i[1�l�%¼�̽��R��ô1$�9l�4�y���#>�ϟ�'�t5�%e�Xz�/��l/C}>��s/�B��"�=s�o����`pp� ��UU�!*�a��������@|�rKT���ۋB��(h->L�J�m�k"oA�!ᤱ�wpxVP�c"����",0�(-�bb�b"�b����	"bp� ��	"�&	���(�I����3
(���"b��H���(�'"bH�4#$�
f"(�������նJ
�)�����bj*q3"j�)�)��x���qe�N.�������6,G��u#T4�Ϫ
��E�"AX�����Ȑ�1�4Y�����a��̀`�sϟ���2 �L4���]�Q?w�S\��7�w�������?�����q�$!y[�����hP�Wt��xg?O�(����Y�g�Fl���%����l�jk�K4��FAU3��%�'Zt�70ۼC#���E��
)�e�\�� ���=��}X� �$

�5 ��W2����~$1���oO_�R�㭧���M)�Z���@��:V��7�Nq1��:;:�C�D5�9���1�*�@6��hY�,�4���RUS�|5�PI.��a��6@��@.��mOjl��ލ㇦|�1�D�&B�))�j������(���(�(�"���B &B`�(��& "X��b"���� �F!"`�
`���=1�}��Q<�9�Mq_�l_r0.�pߪ����N��c�
��I % ��	J��4��(N��SX�՝����&�K�!� �0n�`����j@U>���g�wpV\��������jX����z㗘�����C~�!EK�'C(��G3;��e+ ��(8�����v3`���$�:�U,�` 4
L��g=x�o����E&�ՉEB'`*��{��s �;̇�c��@�<C@*��&bኝ%E⺊kjS0ʕ��\3Z1]$�gI��$��mIJ Ȉo��T /�a$a�0T�ΟeB��eP��_�&E0=�(h�����ӣ�y�έk�S����f�ȣg����y�6�gq�>I��@�KU8��I��a�xN@T"�I1� �y��`UU ��#��^�
���DZ�{�yeU$z?�LF��w���`$�^�� $�<�� ���3GB-'-L^I�b�V�[.FʧB���(�x��@Ё<��8�@�����:�J0��
#3�$@�6i�`d�nʷ!`AU6�4F�Ȅ���4�w�izH���ǡ0 �@&<���'�%L3��P�������*�ݔ^|e�dJ�M�����y���q	����(�9���ܑN$8p4��