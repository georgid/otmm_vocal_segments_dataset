BZh91AY&SY��  _�px���������` =�G�{��&l h �
 � G�ĸc��v2�#FSO)�&�������h���M �R��@d��    jxSSM*hz��h !�  M$D)� @�    ��4�6�ڞ�ɡ���0�$�1L���ؓ�z��@hh2z��7f(����XA�Uj� �w�S��H"����*��A�I%����#��  5B�J  ��J5�D��kFڋ�P�s�����E�BP�t=�8��n<YB(�P8D"ȲJ����#���QC��D$�Z�QI,��f@Z��������I@I.]�Gs�tq�'�K��� �g�_��a�~/��@x���C���T��=��g�\9�{ȣuD<en�[NȁoYX+a�k�ٍ����	�z(%*�����L;��A���_MH�N�Gn�8�`�1��NT�
�bOo���dm�B�Fjʹ��/8���1��IXv)�Xw�5�DL���.�
�9��f[��E���hf(�H
�*H�d�a$��J�9=�H��$$���nC��S&3#2�:��& ��{�@���p/JQ�
"% (��2�9	.C�B�	�6�H�d%�0cQ�@�H��p�N���i#[RŤA&����	� �l?ч�pa�߂�|���}��$�I�#0a$�Z�I-�ӻ��-�S.�I$�$�n����Q	$�I$�I%33)'
	f�cn��C�z���������z�@�h��1�$�|\����D���MO~���
g�l9#�*q��	jږQ�b���V����=X�\<|��ir�͖����3v�� P�	�����
L�@�\���F۪��3f-3Z؟�X@�4b`@��+��
<H�l#>(y�k�f�D�Qd�/'�(�@O�34'v͞B����6)��=���CFF�Cظ$�͏�5�C�e�]�I -���_7�81^�E��UT�͊:�����屽���F?D�m��ѱ��*v�<G[�%��&���@rޟ>l��l7i��l���{kuMD�=p(�`峣bFt�&�τ
6G<�M���'W�t��9�^^�zt��c^�;���³�.3I;1I��xۛ�u��IU�S��w<��u�ٻu���4�M8p������1�k"̖D	�@�3A���j�s������K�I�&Ņ
��m�4�!U�K���B�W!���Af���k5t`���)C�f��7v��L�uL�.ވ�D���m��-��ݚK�(�j�'�L֐�aX���p� x�*H
oE�l�縙 M>S�',S��wma�g�`�}����ɷ���Y��#2�LH��׳$ 1�H��Y�J͗�4?^����R��8!D���=k��TU"���j*�݄z6;5�K�x}�gL>#��}��@��\� ۻ��1��͊�S�1
�=Rx�-�P��m�Ȉ�4e=��2��e9Ż��X_a4.|��ۨ} c��E=�>@�{�� �vv��l���jh��])%kaDF"a�088rL��mv-N�]Ÿ�p1bLH�a~����n�#����l���Ɣ����~����P!��"� 5p%�D�k��Qi��r�?���{���y;��E�ԛ���
�r `Oo�C�V�Ќ�n��/�3���Ù�o��7��S5^"�gñ���,�׻�Ǣ�ڨxTQ[7�W�ړB��,�藹5댌��r�fFW��e��O�O��jd�?B��;Z��&��om�s@�{�0����фnO��c��;���^�7ݣF]����,m���7:(��P�1�x�oi����I{a�n�b_6�gf9��ș}pl  �0�'@�ݹ�2|�v�M�e���Dt�Pv�ǘ��5�:��M��i7�я��P���p�A�xU1��7��c-�K3X���j�V㚛ng�WDEtƉ�����D�V�ؖ^Zu6�4�F�3lS�`7��Or�W�T=���u@!.D�
�� �z߸zdvjyU�"�b�q�!Ϧ�������C2�^��p�>&�}"�#�Őඐ�ى%�D�%�3����덲��Il�n���͂DB���V~������M͚ڳ�"?@��/&F��ƿ� 	��� �~��c�{L�����=7;� -�Fa"#Ӛ��0�3{c��>1�}�2��Y��^��K�5'�q�+oLVR/��P�/VlFiV$}$+޵ՙ���˻�V���q,�슎�����3��{���>�:%�,e�ςUT}/�ϓz7�����X� ��UUVD ����<0��� ӳ�0����2��e��M�iYevע�L�8Uԇ7Fڢh�EETEij��-DUDP���BZ(����*���j�@�wj*����TX�TUDr�m1Q��b""��QAAEGU*�����Q(01 �b��#����	�FM�y��@PR&I10�aћCd�xl ][B��lQu"b\[��P�6�݋� m"c*
��{w@� �
*����k6V�j&���:e�g�g)�����-���S(m�[L�0̘[-�lw_,�z�C��{}vt!˖�X*���f!�Uy��+��S�rx�7�ƀnaC�Ȃ��oO���-��i���=�.�
�Ӣ縂��5�|�7􊫂�9s���Iܟ��=�da�jZ��ȏ8��Ok	v2�*yKL�OW�G�fϹׂ$8���&�ꫨ�op墂p�lִ��]�^�����A)�$1�
���$P�"�EX�X����*
�1��$���$;��Q
�
HY� ��e�Vṕ{�~�5�0�Rw����M� �����+
E�� ���, ,���ϳ�+`�s��{�0Aq�H�j$��LiQ_�%�����ԙ�`!UY:	'4�ʇ��� ���M���Q}�L�R�_�M��)���yA�`ꭆ�;w��ףӁ�U]��� ACY��8�^2v�S��I�L�E��*��[��6�RpB�xp��Ģ����dDxGt@�¸��hK5�Gy��( X0��u��s���4�MK��T�  ��p�3K9CgKE����7�c�Z���&� `�����h�s����P�V�){�P	����p��ά-�' ���ȉ���� 6b�yG?a�<c�� :Q>�o �V��yUo���iU��F�z�Hb	�w�rq`'��Ħ	J����7�T�@͉ǣ���M�X9�=;�6���e�U��:Q%G���B	b3��v���]�4tb��1|�\2��.���1�� Ӑ@Ń���g�*!W��y��)@,��U�êC��[2�"X�r�j�oU�;���[�b�%�.���H�
<�� 