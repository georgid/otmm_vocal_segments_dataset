BZh91AY&SY�ʢ��+߀pp���f� ����av��*B�U
� ��P$@
P��T PH@�"�� Q.  z��E*� $�T*	B(��
T�P��(% ��A  ���U(� �) �%�p    ��U@� � ���8�H� �� ���H� 4��1}۷�S�@(�׾���@{�
\ (ހ>��bӠ.f�zq z}���C����=������� 3�>���B�>@*����@N������cŗ�}��.Z� ����A���W=��wr�W[�} �Kf�g�z���� z��yhu��U� z���R�nw]����R�Իk� �̋�n��.}�ǚ������:�����A   *�(�� �L�|�y��3�P����|_s7�G�oKϹז<ZUb2� j�#)���"�q�j�r�p��|>�\MUf��o(���<���i9�eϷR�����҂   @ � �C'���95]9:U�((����<3�quqaM��7 �ش��o� wW��ҟu }�'�*���v� 1}�93�W��p� >*  �@ �� �}A�RX���w�� c*�j�����4����_GNC��@9/sh, 41�lڻc��'}a��:14��=�x3��\�      D=@��T�H 4   h � ��T�4hɠ  z&��P<z�T��)6��ɣL�&�d0B'�T�Q%      �S$6�T� 2     �@ԥM�P��!�CCFjd���O���?����^���0���_}�����*�����DU]������*��?�EAUt�������UU��ʱ EU�?�)���"������ݢ������լ���N�f��,�O� ��MJd%�4��4jz�KI�C�d"ԫ���k�FCD��^&k�]���@�-K��l9#"�-������Fd��'վ!�&K����H��r�Dm��b��ĐD0@�Z��\��ņQh.���D8�C���ǨD��+��p'�JSz3;��4{j6�\���j�.c7iB��Uj�¬��J�!(0r��(2L��0KNL�&N.BQCE	 �K�8�uieݽ:��;�i�g��1ך6�B-�j�����:�e�zk٦����*uu��.���֪�Ӑ�U���F��BUK��BRbn�!(L� `���ν�����ĬlO`�2L�c�FǣP�%	I�{��$�2�ӫr�*2�R��@�-��~����۶��S���=�|�w��v����/{f�S�����Y�l�硫�}�������~�XuTL���ӷ�=���e�Oż�N�d��+s��΀�&O��I�1"��%��&o���w@o�J:OQ�I���_0��$���[;�=� F����y:=J���]
prF���3��k��::3��q5.:�!0�2\-�2ELzף����7�u����{���ok�!�$�'U2�#�<3��q,��_7bR��1�m��wL=��o2u�R�u;�_�7�Ǿ���[���zo��SM3�^�v,��!�\Y��.xvofF��t{�Ӈ+�u��ڽ�oŌ=%�y��=|�d�X�gj8<���ky*����5�)HTçah�ܺHq��� ���T�Icp��2������ַ��J�J3�=��(06i:CN����fi��8E#/	�_���"T@�(�e��'Ubja��0ᦁ��yt�8Ld%9m��ѝ�#�{q>5	��P�%/�o���ϼ�[��]��X[�cM}�:H쿽��%�OQi�g��a޹;���,"(h� �P����񨰃��ٙ����w�јb��=��S�fn�3���/�;̬��a&�����+}�vl��qٸ�	A��!�T+q+�۲��W	*luE'�2vE��8��#��&�I֣d�bL��#S�����%	f	t��Q�&�5!���&�*N��<�OO��{ٻ/�ԁQj�P�N�%A��:��k���']`���;��(J��MBY��S�qz�B��<�|h��4�F(�X��݉
��TT:N,+�b�[��$���X���i,��ުU�ʀ�j�U���A��0�ؾ��mq��P9C�Y�׾r�ϼ��˖��L�	�w�w{�e>�`��zCr/���N;��{��#�>�֪�U���" ��:�814';�][��E	:B�.;\�	�OCPm�7{��&�3x�uh��2i�)��-V�D�����u�݄�ѐ���F�i�Dhzz�r��J��5!�Hf@aL�JP�t�u&R,Z�r�<��^�u rƮddޗ4xY��v��6Z��0�d,Cwr���!Kc��S&��bb���ci�y����K���P��#�l��]�2���V�n�0lۡ˶,�C��Wai%B*m�b�U�|�l`4Њ�ST�:a��Y�L:���6:��n6BPe:�`hw�N�O�q��z�Ӱ"(H�"��,��Uz�=��0��i[������P�BEE)�g��nۃ_?Z�=��|b��Sf�$N�z�v��ȗ�}�yNE�&BHRM��Ue׳s^�A�WHdi]a�X������L�qww^�j�Q�{C��L{��FC����.y`i5	Ҟˆ�t����y�����QB@�@��i[����}d��+�3�T��_o*��a¢��f>�8^xGxBx�NJ��R�u��	��5Z^���^Z�%M#����̃m����&����E'�d�<G��vN$an��CTʷ�� �I��I�	�J������a����DC��z�%�����bC�6��&�n�H�{ۯw4�H���D�JһQ�[[��]��mi���U2��/���*�a�2��ٶC�8^jU�;��T�ٚ�y_y�Ͻv�T�B@,���/��m||le!*z�Rز�w�Y��x�xQ���Ĥ`;��u{�*���5N��*oq}�3m�8��Mٔn	�b2��ua+K�F
�@��t����t�����6M�J��gk��Ş^,T��R<���Ң�7�:���vt�%'pa��}�CP����N�;�	�%	E�(H�"����o�wھ��m�}�|,]~��پW����6[Z�4��諓aa���יೣ�h�u3��
���>au��`&��!T,־Tf�j�*���a��An��Fv���e��E�<4���2�"��}���>wX����|��P��DuM_w�0z��A��<��SXX������n��1�Rp��o��;�7���̖��&R�R5K��mw�f'wzVҡr0�$�d4FK&m��8�U��1�$���7׻���e/:r��w)��g�3����d�p{}��e^9Va�<$��T4������*t��a����L��]i����m��Q�[P��SU���b,5A�`G�-]gl���UŻ���׆֛�bI
y���d[�a�:)12�̉e!�oj��ώL�������2�Fa~��kx�Y2�m�:i��}x(z��y�{V��d�厙֍���QV[>{7\yųW����n$C���cPv'JZ�
!�?,��%�f���O��-����9�'j�R�h��L0v�Y���JeZHU�}�*�����w7��x��х/�)�Bĕ}���g�n�!��O1�7���כSu7ƅҊ�{�����'���P�b����Ȫ�(R�����ӽ�F��s�ɯ��1��r�����(JR��J��>��L�Ώ�.l����W�񉔶��uD��2*t�՛_��֜t��J�0�!băO����9{X�h �MD*/ȡoP�wTE�x�;��,/{��ݐ	�%	i0���7����&�b�g��I�=��21�'$�X��P�LI�Q����`�V��n�e�rf�
��BS��a/��;�������D�$""�Cp\Z�%Y��@a�%.:��%i�)��a��(pF[���K�P���N�����ք�����᭝Q�^jpܱIQŝ~���Ë2���'+Fv-U	�,.,0�?����;Q��{x��8���Y�3�P��oz+>>����Z���`^K�jf�3h�-�Ӎ7ov��P��;���B� Wvv��޹^�{*_ec���=�we��y�.�����=P�P�Mz���a�<rĸ}�}��n��aQ;�W���P��Vv{٢w�;/��Z�5%y](3�=���ھ�����|�ط��y�)u�\�ޱ������$K�J�����;=5�N�P�w0x�*��d��Df\6춵B�9�6y<�{�O���19�]�őw;Ɛ*I��2vi�%�ؕ�V��C�������?��Z�R�j�W.Ċ��- *�� ��LZ�D���÷A�"���Y<��*�<�	)�,�0��.�?�%�ɉ�����F�%+�%�y���*
X₾�W�hv!���R�%���R7A�J��)pO���9�Ӆv��r��wt���m'�y�H��E���G'���=h%꤉s���Ո�*�"��bX��D�P� �J���~-C�Z���B�ŗn�n$�&BP�y�r6`2��'К��M�� �Pc����:�D�a�J��%	��%���u��jO}�I�|�V�D���X�𻺻��}�HV��u@Dṟ�;��%ϲs��ݭ\��g	"Oa�rW3����^vzե�تP��'b��d8�����8�R���ʤyf�P�q4��`�ێ��>Pʭ`��y��:�>ք��^�X3�מ�NtwI��:��:��#6��B��;�Т*�Z�}���^G�&���i�"J�'�'V��=.ROo1���w�X���	��2�m�w/ޕt�e11P/��t�ܸ���4ƂX �Z���.SQ�LP�Atxvgr�Ոdn����v��:\����y{d'w�.ٴ���-/mN6u�`Ɏ&��>�:���%!�d�\,��#��15�`��:^UO��߻H}���x�)�~�޿-s2���e!ɘ��f�d���"��ru�:�f�A��UN��*��c%+-�X�1RM�lY�i{�+ݟs����A{g<�z�2��K��Λ��.qg�yA���B7���&�
*��dw+=�ms�Z���������3+l��GR�1�V"�E����߼�I/�}�Ḳ�O!:��:��O!;��'�`�%	����~]�3�=�{�Ǿ,n�Y��!���`p��*��e�y�a�Î:�p�5�
�Uu��,�}AfUUB���"�V]a�� ޷e�#��Q��զ���͆5��t���I�eZ�u���c��x�s�z�Y�d��e4I��-�ֈ�� ĮBd%	f	JBLDa�V$C�(��Z4�M��ePh��2#0����$�n�#}h���8c9׊+�#��RHH`�`�RP�*�ګ3���Ԫ[��C�nC4�@��eRF��+�.D�(X�%����C�L�}�{$J2��#�,���6x�:����4JjөD��L��\�b���3Y+�Ⱦ����{I��d/&Wf���{Vw]��x����Yt�֋�D���α�ީ<nZI�|F�[*�J ���h�"��X�%|zp���}�K�ɪ�*j�����3Q>>��v{ם���ԦE�2X3d���<��8�!�%B��N�L��))3zz��RF �/-W�пKu`��2c�[����gj!�,�+�2�q�CM,t<uєkF�0�� �2���E8kVZ�2TĨH��TU�������w���_�}����~  6� �               H� m��        �    m��    � �                   �                     ��ݮ]6m��H�j���v���q�$dI!�ć e�`$ �[m��p f�YIv���WP����[l.���� �/k%�Q���ʭUT���Mk�"F�+R�c<�W@U ��U,c\������ؐ�h6�6� T� 򻱨z��m�� ��`�����	 �`�\:� �cd0  H  ���s�h��&`�`*�n
�4�L�kX 7m�[ �I�2��tFX��*]$j�t�:8��5��m���T�(���N��R�7G���k �;E 6ۭ�M�*���������˖@�]N���Fٓn8�:�$� *�����RD�<�ŠI�Ƶ��6����m�  m��       ��        �              ��8   ^� �     [v�                 ��`     �  8�m��kz�����     �     �  � �6�   p    �  ��A�m��;��H6]n	 m���7K�pH�xnV�v��o
F2�՚oPL�4�kP�:��P�F�8�6��m&�TI*��N��5�m9�2dh�6��A��UU��j� ��.�JAīz6f�l �X�a�*���2*�KUVç��c�hm�:^��Ɩ2���v���
j'I$'�}�}�9y��c��'���<���[����u�u���z�'��Þ���=:.�H��Y�j�`���[8iV���T�j�V4R�pR�媭�y M���p�5*�VQ���z����c���� ����[�|��۶�lT��I'.��:�n��oD�z.�0�0,��p؇n +9�n�U�CX�WA*�b��ڪT-�9��9!��Խ��ّ��t�嚅�[k��P�ۡf�VY�[P*����pK:D�l6�� /�Y�Xm�t�i�6��6դ��@�t��v[�p�ˀ �Xj��y���h�G7n�������q۝����UWm�veUjy:��v�<QSv��A.�ڰ��j�}n��u\���+j��h���Ѱ����;���s�6�c��e�rʶ�QF��l����N��0mnl$F��Ae$�-���mv�r��+���웛n�۰��]W��m�l   hk:���$P  �J�FT���k�`9�:�� �  UU^V�ȅ` ��T�Pv���ؠ�U��
pUU�[ ;-z�H���n�H-���m���9w\9P���y`���]Uζ�UJ�V���UP������i4�,6�-�\ְH!��迍�}W��V�{lF����Q�.� Ye��od���[�,Y7���l 3�e{U��\<�����y[Ϋk����8�W8*��uR�0q���Q�2�ԫ�up2��i�ȢQņ̮�!Cf��u�9$�-����-n��uU�=��%��Q��{j��]�@�o�ca��
4�Un�u���'��CPՇ �R�T���,�;�t�.t�2KlUV�W,�\�]Pm*�-WVʻ�*�7ѵ��5���R��fZ	�Z�V�C�Ŷ�4��$�K�Uv�V�衟����rL�fհ��[@M�=��[��e�a�WM���  mۦ�cj�m��Uʲ�=/,��n�F���+��mf`	��>�>��6�|�UQ��a��T n�a"^��E0��.mm���6� �K�1�zu$�.�Kh8 8����5�=+���8&,m��6*��*Y%Ç ��@ڶ m�
SZ��m�ݛt� V�oP�v�6�yek��UT9�����{l����ր� km�zV�:Z����7	�     �m�6�3�~��U��   ���)\���l��PJ�/lm��%�"j��i����nD�l���a�m�@�,�WThV�Y�~��$�>ф�CRPpLUUUlH 0]���w[����;l|�(����V�U�l��n���\�UTn��ے� ���WU�h�$�5��-�Rg&�ʻ-B�n��N8�T��e'��u���ns�&`ٙ.�E��MK�C}u��dU������\�"c�N{5K��W�\����M�,���t��upj��rfpCRθ�M�I��ѷ]A�&�p�S��kn�X�n�|Tk�ym��}|��蛝 ��9yK�6����A'll���bK�բ�4�I/;�D��Um(�*�iI=��t�ػ��HQ�J�PV�췇�t�-�hݎ�VU�1�U�ԇR[\�H�UJ��O7����]�gEm�� Z�{+�y��+Tk�GIm�,��':�i�&Cl � -�Z�e� �Ͱ �l6�	� �`�Cm��`�amp����fxn$�M�n�Lf�8  J��.�I�qv��F���� I��Y�`�9i�7  8 �  d��l�X�b۶�m�p6Z�-��`  	a�aä`��l� 	 oP[l2�h���6�6�� p ���%���  m[�9$��2M��H  	�N��� []  $�e�   �m�m lݻ6�m�
u�U�� 
���쁃�@W��k��l� m�mq��R�v*��U� 2�p�+y  �m��i����� 2 [�e�m� ְ (��vv%��j4+*�㄀[@-�c�B@  �k �d�����`  ^���� ے��aj�5�Zl� �K!6Z��#�V:�Q���-�6D�K��ݲ�R0I�&ճlm��m�� �l*ޠ      �%[I6� [�tn<�z�i�nr�mZ� 	;m6�!*��UUFAY�]��۩UWj���\K .���L $8M�B텶Kh l ��v0 m�݀���[Sj  mm�+����<m���`s�H�,��g`��M��-�Hӗ � ݱt�� m $�B�p k]cX�m��]v-�$  �/Zpsme��h��ݶH�bD��Y6�K$�\6i;l >��$�ʪvH��U�������8Ii��m�@&�Tk�FZ�Uy����vYܱ*��C�pm����K#�j�q*�Yŋ
�.� 9u���\���-@U��Q7"�.;t@U.P��a�t�Ht��(]�Eu�8�<9t�vkG����[e�@u:�9�95�l7*��o��}j;�ۭ�^�8����p9t�h.�����;8�x���c��*���]Umu+ͧauԝ��x)V��km ;��ѕj{B�ql�c�R5\��K�/d�vں���m$��SDu�[-A�4��[��4�/u�[�`iR�C�X )�۱Yx^�Ynj�$f�k����V� AHq�A«@�n���Uy���Kj��6�^��mh����\��Wa��뤸�{<�����D:J�� 3�ԫn�,�Y����/2��Td�[R�T�^�t�g �5�Kz���X�ml�UR��"nY�#������I�t.U�0��]s���W2d�v -��1[I�-��nŮ�T��x������mK���E-�(���:�$r��UW=itݎM��J�u�]��.�N�R��64�����^�Ǜ�6���ms�x��tHlc 		ӂ���7m��*ݪ�*�1�>���A�����H�v�tWU*�vX��k;r
�ѺsU�����n�1[J�cڥ[��%��    Ӷ�6ۀ-�E�a��$�nͻ6�M��qp6ضMz� v�@ �T�uנیlST����Pn�[K5�Y�-��Rm�ׯY6ݶ�  � V�[�R]��e��^���n�6�A���;꽸�tH�����9] p�'�ض�i�J��.Z^8{05]1�4�m�U�\�.��`����c���-v�݃�lmF,v8�ݺmul��zn�l��N�v1�N��H[�u��]��U�v<���s{'g]�*��y[.�غ���&k���J����X�n� �V� ku�ֱν?�[���    �m�:C��;e�&��qJ7*��ٰ�-�(  ���!  ����r�Om[ $� *� �������ԙ�� \�TPUVP�m�b�pR��/N�5�	y��t�h8@��۠@�*�)�Ct��AoieZ�Z�	UWj���W\.�MT��&B;(��P+U�+q�5Q�{�S!
�F�^W7L�,�67n����R�hc�t�����5<�#=;�w[m����Һ�:�sA�k��A�]�ѹ�i@W[;]� A�U�T�T�    ����{�������*!�����UP_���lO�����R����?�?��W���@ ���A� B�dv� ��� 2��*t�v � ��Ch��#��PSj��SH�	�� �����ba����	"�"j��$�`� ���������HM*|">��
@�領%"RP�� >A('m�0A�'��C�ID�T0�21IA0P�P0MD�5K@P�dȤ5PR��,�2�2���KR���}P؞	� 1�ED�DЈ)�4�@� �� zڝ��#`§p�"*x�������= �FI�Ңx�>_EBE�A6�)��(`� tu�8b=���md��!҂z�U�}L1dX�J�a�e!��Y��Q�IT&�D���4 �/�`.('h�
��#Ҿ�/h��R�(�T� @�.� ���*��O]
H⁈"l}z�����S��T�4B��|Dz 1E;P�TM��E�4�����U����������?�t�p'�U��heIP
A�P�JP!P)REihp+�"!�� ]�u�ݼ��  Cm������C�   v�   �r�z�/2��-�m��4=��G&��������6���qqKh���($acm:�\7Sq3���ȁ`���3Уv�*��Ы/ 춁� �� jؽj��   $�[rIs�6� IJ�m� ���ƒ�]���[n�f8Gtۚ�k9���t7��z0�d�ڥ�7m�5�C;:ݹ���:�ma+�ݔ�Fw:�.�s�8�zprn�#v�A�mlkbwn��b�oh���an޶<v��p7jw�V���m�0�8��g]VIq�	:i[{mCz�ӥn�`.ێ�+�.��ۡN4���יl�G�����.��z5����M��8D��U���j�:y��r��.R��2�m��q��̮��!�6���=���)w��M�I35$J�Gb�72�ɂ�:���lhW<�u�	����X^�I-)��t��M�Je�����t��g��勧�y��k]V�:6)��su� �n�jRQ��>\�!N���J�v�51!��j��km�����Q9�c �� ��[Q��o4���َ{��Ul�� 8� #Z��Ą�w7i�EJ�Vwd3v��[�J�Y:`�\,E�ڔ�^W��+��]�jڌ�[�kXnݒǰdi�kӶKs/Z �J��n�:)N#�T=
���qs6��Cp,���j�u�-�,��nԱ#tHp[g�(u�N�KE��"�j(�Gg�΀zk-�\���+v���N�t���ro%�P�2��-��:��]�ֶ���;�X˓V���&A�Y�.�����8�s��<g�����1X⺻c=�}br܀�R8�����i{ez�����tU��m�l�b�Wv:6�D�p��Z79�'�u\O;Þ����+X^�nm�����岃PS���L�*����]�;�[F;���n���7n<�[���V���2�N�O]�B�������ww�ڣ���
��Q {?�	��-'�����(���0*���?��Wwe��ݑ��M��n�nێ���%����B*�۝D\U�n.�t.B����]��>7<q��z�cA�%��8��{f�J�.	�l�ѷ8lr�<���[��w4k�n���4X��I����AbkL�gK�O�vv]\i5�[����\t&�i�]0n���۳�V�^�#�Ay[��u#һ���U�^�}�w��{����"'#��N�g��v˷aU��e����a��!�cb!3U˅�?�~LI.�F;�� 7�� 7J/u���۲�n���x}�L �w^�-��=u�h�c�Ht4�;M��צ w�� ���{��^��61[
hI��l��u��ݼ ��^�k� ��oF�.ؗͻ�v��;�x����צ {�� �Q����Uݦ�I�z6�G���C�46��/9�1��>�Ls�V�����-�튄�e�x����צ {�� ���������ت�Hw.]�K�>�� �E:�/{�I{�� w}� <��A���
v���ڰ>��ş���jU`{U"���>��
Ճ�WV�v��;�x�n��צ wۯ 7J5j)�Ӣ�ZM� wۯ �����;�xo����3��/&�N.]���up6!���^nH������ƀjm�x����T'i7�w����u��ݼ �^ i�m&�+���� �^�-���u���0�v�M1]�_6�����n� wۯ�U�V�Wʹޘ�n��m��C�N؁?�m������l� �� �^�-��6�K���j�*�jݦ��;�z`}���n� wۯ 7}���]+ht��o4We��1����[�md�]E��ė(�XX���+��L)�f wۯ ���}���n�����HV�*��S���-���u���0��x�
5^����$��}���ݼ'�W�v{dx����M�v�n�ݧi7�wV�����yn�r�D�ң���]o���~���n��դ�[N���x��o ;�� ;�� �E��+Ywn�Vخ�]1���+��Wۮ�:�T�җM�J��V,ͲYt�n�ݦ�yn� w}� ;�� =�׀vͻ=�t��'T��������{u������o�Zm�
�Z�i����� �w^�y��k��J��A��n�o =�׀s�z`w��������n����e7�s�z`���G��ǀ���7�}F��av��ݍ����;�|�n���OF1��8{9�*����F1Ԁ
][�p�׫R2��t��8u�&��6{>���<�M��8���d�ǭj�=[��fX��{v9�<�&7�3ۍ^�-G��:v6��JC���q���$lj�i)n�mN�\�4��8���;��C�so6}u!��X�,=�]�\;�҈��4��S٦�E�J�g&���{�����2��+��f`�����&��*n�u����ݽ6����|��÷"?��c-�$��I {�׀���9�z`��Sj��v�i�v�x��^~����7dxf�`wu�M��hcj�j�i�M����o����x��^��މ�
���][����� ;�� 7�׀���;g��j*v�	�[L���������wƗIQh�U�m�r$Sn7az��F�z��VR,�\�:�䶵��R�m��i��'i��{�x�n�{� ww^ h{ԩX�i����7�����߾�^�#2B��bY������&)���#+$2��0V��0�h,F��|� ���������w^ o}� �yn�VZE��][(i�{� w}� 7�׀���ЭJ����`��`w��{�x��{���=u�V��-ltݦ� o}� =�׀o���k�9�v�߽�BVv�Q��>�8�wQN7eun���yMY��s-i��\gM��j#�o =�׀o��������9~��4�]Yt����o �k� ;�׀�׀���;g��j*v�	�6��������Wܪ��U�P�zG�w�� �^��-��V�[��x��x��}�L �w^ hnҥb��"��-�o ;�׀o��������=�k�uW{���bm�n�7��Sch��F�P�<�Z�k�}Ht�@�.:j��I]:Uul�����0��x��r���H�@��O��c-�M� ;�׀�׀���7���=u�U�mU��N��������u��z`{���}��'ce�V�ؓx��}�L �w^k类��n���v�N�U�0h�v��7����u��u�{��j�,=J�vM�+u���+��7�ZxQR�&'M�w;m�W��:E�:�j�v&�I���L��u��u�{����0U�{��l`�I[I6�}����x�^��� �ݤ��[LE[t[�� w�� �k� ;�׀�׀r������
���4���꯮l�`�#�����UUw�H�@��O��ݱ0I�`{��}����x�^�{����#O�U�h�/$a���7q����h�������g��'QŻZ�znۙ�q��`���wlNc)ͨN݋�������c��ZӠ%��jt��nx.V��R�N;k��!��;Vq���:mԬ툆���A�r`J�)>}k�Wc���O�X�<)��� uFYK5#���u��8�-��:�G<��ɋ��ݴh�b��:Q�v�k�����V��ߝ�}�;G}���8�Apd�sn�$�D������'/�3���mr�j*.�6;?s�����d$�M� wf� �^�צ w�׀;��;-ڴ6ě�{u�3��@�R,۪�}�VG��MMP�*ݍcM��z`}�x��x�n��z��n�&[,�m3	E�vg�do����էݭ��i���R��I��o�_Ҧ�NTء��}�[��T�ܭk�1��6!9톫�$�f��VN�rmy��;%9gJpKslܸ�O�{����o�i�����������[�+UlV]]��^���D����{���;���hV�[�l�ݦ	6Ͻ�������w��^��>�s�{�햨��N�I�������ە�j��s��Zi�i�v6[�hm�M���+�է��ws�����]=W`*ԭ��zg�ۓ��t9N6���Ӡ�+�Ywbwh륖2��v��B�q�=�ʽ���ww_���r�u{�n�-�	�6������v�7�m����fvwͬ�&�����rGq˼�~~~]o����T���*�ve7����R�aդ�vm;���ΐ�(�;�d���5�7�Fj8H����a擢�4&�@I�Os*�z9�1��&�t=�!Uk2��鷲���2���� F���T�޳e�MQ�F)$[K��f�h��Y�V:Y: �@%u-	��ݸ{��K{{v���c gݺ�b���-ە��8���
�<t�oN�7�����n�2`�Hv��SN$:9m�1ҖaD���4�a�4��:���R`vlOz���mY%� ;/�*��X�l��R(�Th�$����Pʶ)jKMf��],�S�f�XGN�6%WvY`�S�{`�TJEO�CH%��P�R�vuQ�r��H14ѭw�2�������ꔓ,Kz]!*�.m`2�R�*d̥Y�BI���VYB�!S�U]D�:���D*�Y0NXLJ¡U�!Eن�W����:@~zPF�b� �A_�@�"��� x�
������e>߻��JR��?�s��R��\�Y�\7��Yo[�JR��s�}��)O���t�)I���r���9���)K��J��b%���(
��g�݁ݷU"�)JO����{��/y�o�)JO9���}A��z-T���*��v���&��&囜u���'nE=Snr��>+dҌ�����kZ6�f�7�ݭo{�R����y·�JR����R�����b`����%�Ż�;�;&����2�$EM5T����)J^��JR��s�}��)O���t�)I���r��3��޶KjX����]�P�P�����+UP�>���Ҕ�'�{�t=�R���7Ҕ�'|��f����3yoQ�g[��Jﹾ])JR}��Cܥ){�s})BHk��Ӄ����C)'��������y�ܥ)��3�f[5�5eka��})JR}��Cܥ!>�ڏ��_s}�ﶣ�_h��kR�	�u���#{m�vc���E��5ă�`�0�s�ΛH鶭q�{����9���)I�=����R���s���˒����ߺ�)K�~�kVkW�7���[��Ҕ�'��_s�JS߹κR����y·�JR��s}4%T$V����vH�%����/Z��S߹κR����y·�$d��7���)I�=����R���r֎:ٸ���f����)I���r������R�����`�)J{�9�JR�������lC��r]�Z�����?7Ҕ���}�~��R����uҔ�'�{�t=�R�=	�i�@����:*�_~Mˍ�ڸ��˻���<�Y�0��1�	i�0�ܼ�(өR\qY���Fj���!�VyI�Y�A�n��'K�9ء^���.z7����G�����j��n&�3�[�ȗ.�Q��c��n�f۬��=���� ܯC��%��4�������8{I��p�����l�nNN��#����㍱�m[����M���ݦ��9�1\��<���QH��Q�(,���Ɠ���q�ۡ�������ԥ�un�2�3��cb�s��C�OW&�M�f��+_�{���ow��_��ܥ)���.��)>��s��Vv=�U��;�;bBQ54���AR5k:�X=�R�����JR��=�:�)K߹���)I�=����R��9�f[5�5ekn��wJR��y�9��)J^��o�)JO9��r���s|�R�����s���o3e�k7�����)J^��o�)JO9��r���s|�R����y·�JR���Z�F�[���-�{�JR��{���ܥ�@g�~��Ҕ�'=��JR��s})}A_s�r��-���Ub4��$f׍ZeF�s�`}�OdB)v+��ν����\<��Xf��[��JS߹�])JR}��Cܥ){�9���)<���=�R�ܮZ�(���o7�5���JR��=�:���f�2Fr�33(�� �1[1��=WhnR����JR��y����JS߹�])�EL�)=������ff�kz����)Js9���R�����`�)Jz�"�����%l�;�;��5T�MA4�13$�S56����4���σ��~���JR��y�9��)J}�s��JR��r�3[��՘l������ܥ)�9�])JR}��Cܥ)�}�k�)JO9��r������Q�ٙ�h���gW�����vX8w�c�ܲX׭�fY%�p����\�q�z�o�����߿��s��R��>�5Ҕ�'��_s�Hwo%H�vvo6��������&f*s[�Cܥ)�}�5��I�JO}�~��R������R����y·�JPВ�-R��0j�Y��}A�vyo0{��<�7˥)�A:�S�vRg��r����9���)<�>�5ѽfh��e�n����{���	���~�R���~���)J}�}�t�	��O}�~��R����l��5�q�f�f���)JR}��Cܥ)�}�5Ҕ�'��_s�JS�s|�R��������*&Į�6�]�B-�Af���a�ή�q�,`��R��Ɓf���]����oZ���)O�﹮��)<���=�R�s��Ҕ�'�{�t=�R�d64�;��$&4�Ͼ������e�r�����t�)I���r��׻}��P}\��&��)��M�<��R���.��)>��s��R��>���JR��{���ܥ)�}�f[5�5ekn��wJR��y�9��)J}�}�t�)I�=����R�e��*����������Ic��nE��jR��>���JR��{���ܥ)�9�])JR}��Cܥ)�}�,4kWƺ;#�1]��ӭۃ������ا�ݐ�lv���HQ���.m�ݛi)�������`�)Jy�o�JR��y�9��)J}�}�t�)I�����F�kV�l�-վ��r�����t�)I���r������JR��y������J~�\�k��ka�f�f���)JR}�߿t=�R�g�s])O�@��=�?s���JS�߷��JR�����[�0�ff�kz����)J}�}�t�)I�Ϲ��R���.��?6I��~���;�;��TԔPPL��SU6���Ԟy���)O9���JR��=�:�)O�﹮��)$�{���o3Y����cW�js[�e�m�χ��lWEqT���(�/EN�#�Xֶĭ�F7!X��zݶ��t)�(۹Ğ���I�70-�]��Ύ"|��kN:�Yю[<YTx8E�m��F�Wh�JVq�z�.Z�;�����)B��틫X?�����ِ<;<YN.�.�x8�o	tXsmu\��[��������a�.�oR���uF��B��UG��<T���e�s�!t.�>Q{C�ZK�Ͱ�⹠�{җGW��d�WE��[����~߾{߽�v���}��JR��y�9��)J}�}�t�)I��9��R��>��3-�7�����޷t�)I��r������JR��y���)O9���JR��ӌ���2݊H�r�UBUG��&U
R��3�sC܇�c%=�����)o{{��vv4i�%�5D<MLUOJR��y���)O9���JR��=�:�)O�﹮��)<�>��������faj�ַև�JS�s|�R����y·�JR�ﹾ��)<�9�4=�{�������,e~�h�m�뙹	��.q��o�D�Χc^[)v���oY�ٽ�wJR����9��)J_}�7Ҕ�'�g>懹JS�s|�R��9z��V��n�,���
�T%T/����"~<H�0gs%��[3ġ��P0R���JNs:�އ�JS�o�Ҕ�5��L��}��V�64��6��+M�o})JRy�{�h{��<�7˥)Jv��%l�;�;����݁݁�����fݚѻ��և�JS�s|�R����y·�JR�ﹾ��)<�9�4=�R�gќ��n�Y���޷t�)I��r����s})JRy�s�h{��<�7˥)JO<�,5�֞[3[�[��+Tۍ��	ru�'�i�Bh�%$'��܋5�#^�D#%��Wd�(��+UP�P���o�)JO<�}�r�����t�)���[>��h$�$KJb�ɠ����R���������RC%=�����)>��ߺ�)K���R����nŔڱ�N�Ё�x��}A����R����y·��E|xl�RV��݁݁�v�g�݁ݒ��1�l7�������)JO<���{��/����JR��3�sCܥ)�9�])JRw�^�r��[3[7�k{�{��/����JR�ʄ��}����JS�߷��JR��=�:�)O>��k,�[�7�;Q��n�*�!m��yG�s�c(.K�u��\�Z�a���l�p�CW��m�v���9��R���.��)<��s��w`wm�������	L�Ӕ0�Q�wZ�Z�)O9���JR��=�:�)O���Δ�);�=�4=�R�gќ���k-mݽn�JR��=��r���k�gJR������)O9���JR���0�5���ֵ�Vk}r���k�gJR������)O9���JSްŌ����b*��X�i��*��LE�$�I�V �	�3E'���t=�R���՚5��6�[���JR��y���)O9���JR��=�:�)O���Δ�)>|=03>������&�9:��2綼�&1�\;u/�)�WNN+m\��/�q9���>>�����Jy�o�JR��y���{��>�_s:R��������)Js���\Ֆ��޳{�{�)<�߹��)J}���t�)Iߙ�9��R���.��);�K���65c�]�/
�h��>�}��R������h{��<�7˥)Jk��̯�}��V�6[h`�WI!2�yҔ'~g�懹JS�s|�R��o���g�݁ݷgT[����	L��o0�{�ލ�k}h{��<�7˥)J? ���?t>JR�s\��)JRw�{�h{��?�?�:?��/)�?#���2���Ɋ�/�����	k^'��Ud�uRv')X�D��F���BN�IJ���'�n�BȺ���P �m��!*UH�)ЫƳB�C;+�gZW��4v�,���׷k8�`���2��Aט�Led�E�Q�powj�K3-,��fvfeإ� �f1خt�zj;0��-��X�f��������Wi���bF�pU��P��\�UIܳWu�(��9<�aJ�����b����\�7������_��a]x�,{�H30e���Y�%f��BBM�i�m��:<gFS:�e�B���`��b��� �m�$]����%uj�v��)�7���V�f�0l��wԁ�P��Zb6�螵����N���κm��Q���j�{vn�0��#�E.vP������N�e�'.R���殣�`�@���+����Dޱ;ۦAS�!M�K�>�m���  lm���C�   ky�  M�ɒ&���J��8�R[�,�i�u�S��OXh g���\ki
�#;�m]�������q[��[�]kI�]�)���Àj�� p�H��m   I��Ԓ�� �MٶÀJ�nIyyzvݝqm�,i`y�Tp�: 8�W�DC>��;���wH苧�=��t���R_<]+ǂ���1�m�y�e9�]"VM���p��k��[��]m�,`7i�^��K�&�sn݊�0)z��q
�\{švp� ��=+Pͷm���
V�xw\���;sm72�����L�Dp�_a�9M.������Uo�`�wՃM�����]%[k���1��!Μ!qs���D�y���c,��v
]��g&��,=1�F#V9��CvB}j���U�����|f��j�J�n���ۦ
��;\襗���V�os���;�m�q;&�4c]a���g���
�WG����|�������˪zc�0Doj:h�㫪1[�ۂ]i9qpQ�:�+)�sb�]��ܕU��`s�] j��nf�	B�%�ĳˌ1G���rj�j�w���%宅[{W�[�C��㊮�u��峡y�r( R�"���pw�|b���V-�UP�F2���������*��J�����}�٠�m�kXRJ'���c���Qt󥌺tN.�m�n6�s�nD��N˹9�x����rGn�l��.��Ҵ���6�A��/�Y�.�X���ۭ&�ZL��9�"u�A��mPU<e�o3�E�l���Ղdt���`9��8�[���S'd.��[��U#�qךX�z����s�M�� .�y��v�Nz�;#�^2*&�GG�n����F9���[[��[��d�"'&�Ƹ�<J�r�U����h&͵p饩s7<@ \r�
���@uqm�g��/���Xƹ�1���7�f���{��������}A?�|� 0��L�`#�1x
@	�N�ER�Y�r�IJ���[BP^��C'cc(c��6�Ku�Q���WGʯv�N˕�]5�΁$�^z�ԅ��[G@X�qR<mX���ptuѴ�n�<��n��a�;]sv�^ΞJmq�y���]%�GF-q��p�|���h�iԧ�A��M�-/^�q]�G���z	�H�;ǒ6-[n����V��g�4���Am��Q�1:��.�j��w��﻽��t���G�@M�-kKǴ�q���Q��f�]Z�����Y����e��e�E���z�ڔ�'~}����)J}���t�)Iߙ�9�;��<�7˥)JO�Na�ke[٭kV����)O���Δ�);�=�4=�R�s��Ҕ�'�{�:�)K��j��o[����)JN��y�r�����t�#I��·�JS��3�)JN���tov�of��-�����R�<�7˥)JO<���{��>�_s:R�)<�=�4=�W�T���E�:��v[m���}A�w��:�(_���Δ�)<�9�4=�S�|�"����D4l2&d�i!����"u�:�xwk������ݠ�x�y]�%����2�PKYq��X�ڸ��UBUG�:�������p��X��f����wClBHL����2���_UnbB��2�0�+)��Ŋ����0il'Vh�ZD�49�Qf��X�� f�vhh�f�vgkw��yj�vuE�9٘vh��隚b��"��ʫ���Ł６`���:����Z� 7�ąӥE$��i�UG��9�7V��;�6.���dp�6��Ԕ[`�I���7T��w�l\�8`��~�߿~~��p~Z.l�.k��%�e�bլ�ݸf䵦 ��\XT��ٖ��u��ܸS*��&I�ީ�pH�{�������3��S���J+���j���i�*�p%H�gg�{V`��X�6. Gj"ĝSI;-���������s�������;�IXB��)%!�X

I%d%T#��{�?{����,�y�TH4DSD�1U��ݡ���*�ޞ]8��Xy�wfh��]����wI����2�w�w��x���n֖��f�R,�x5�{�I��ke�c<�8sl�9��t����.q���ew@�M���t[״U��}�O������7e(�vv>��p�v��t�-�o�4����p�ﾠ�R^Ω�pH�W�+j]IE�@�)�$���7e(�3�Z�ggg������j���d��MM5���334}��Ӏouq`{�j��ݝ2e�� ��:�:����3|��ٽR�t���x��p���������K�9�6. {@���M��*|�[���f�HO�l���]��:.�19��+���t��uM$��L�=�l� ��/ �ҵK����H�3�C*$")�f��*� ��Qn��}+T��H�=��f�����g�G��jjj`�������>����=��`{�j��)E��#��]��2�ܫۼ���@0
���T�߳�`-]�0)J,�ߙ�vh�ӽˀz�K��;�VU�Wn������pvfngfۧ����ӽӀ$����~~H ����'������@l�<e��@�ZZ�yh�\����*q�99���SG�ˍ���9���d�˛ib�+�.v3G3m&��9-�b��S�M����]��^v�5��d��2�j8-�����FF��j�ƻr�&x��xg#��]���p�w`KIn0lO]��,q���v�{-���)]%ç��6!��Z��m=�L����}��a��[����-5�e� ��-���9��⚥zz��m\��5��twt���)�T�������vݤ7W~� ��4�-���ɠ����3��S��;7;���wW��� Q$Xo��nc���t���$��Uy�s���(H�GW�?��溫ߥ~�8݈WM14�D�EMM���ó<{ڻ0��>�%8�;p����Ł��9?Q �SDM5LUf �%6:�"�G���p�����Q�c���S�'n���Kj��dȁ��cq�f��W5us�{�ܟo�)�f�
6��>�%8J�`}��c���
S`rBD�v[*����<\H����;[�;;U^՘��l�|���gwp�B��9��o���f�{���W~�BJl��������ff�l�ߧ ���~,�PГ40�D��$Mf �%6}>Jp�"Ævgvq�f�{Wf pw4�'5L4AU3S`g�� gf~a��v����=�]����o����D��W�y���v�q����#�C�ˋ۷%#��]�n���s�V�^��j����T�ｫ0	)�g�wgpwfٜgh�;�8%�M$Dӫ5���z��^y�����
�*34�����`{e~�8J�`g�^SH�ԓMSY�(IM��O��1���3B��6" LBHuo������?~� ���wBm*��1�k����������\�5�_�������j���=�6��t�MA4CU�i�z�Z�s���W�$ �T��{W_�DDwt���)�7�l�*"J#��[���nC�qj�ɱ�,�mm�Ք��7j��?TmPTS�kZ[,hn�n�������\�`��I3����Q5N4�32IY�twt���)ؐP���?��wW������<����`	���+��5�5��f�����7T�?��6G����{$Ė�>��`�՗ ����&������3�u�`}���cR�]��4s��Q$��CĖ8�TE�MPI�J'`���{ggo�0ógG~�V�GM�NKM<�1Wm�`�� ����>�0{�ZX��%� I����E�Ձ��c�o/Z�痠݆�s�S�i�c�����{�����AN��
�΁.~���}��H�n���;<����p�*�����"f&����>�����3�A��Ł���0��g�W�wa"m;-�wLi}�O �T�>�Y�<B��6�ں��v�6df�n�kwT�� ��߿~� P����>�����g`}�,񿮿'i�WcI$R���6�E�v�폺��7˪���s��ШtH� 
2���eq�	̖h&�LB���Af0�e�$�"rȪE\��qpb`��N�{���_���勮��9gD�wh���V��s�2��F�v^�Y�,�5Q�Q��2�˧%��	whi"�|QvW��m;=A	۠�n�Au3�-��m�F�z�V��t�8�n��ݧnb��ohދ�xW�M2��*�=����iT㳝Z��pK����ƞ�W��j�{�^:f�8������Uգ��qۆ�B�Se�����=�c�W�j�:跦X�^����Ӥ�`{N�l�m2�=�nYm���w%�QG�@�m+�d��*�b�&���.�Հy*E�����{"�9}��2�MӵE1]<N��%H��ٜwf�;3���~��G~�6���V���;3�ܣ�ɧ%��HV��L�;����odXo����qbKx�m�S��Z�X���K����O�gf~���l�]��%H������;���}����:?�*����i"f&��k ��� �;�9�6�E�{����ۿ,A9ղ<�;�<�ɞ�4�s�n��ݧ�Y%�ܴڷvm�UBTfb�I��e]�_<O@�ߟ� �}'8�Ȱ�n��;{�D�t�ʻ�t�b[���}�;�'kDϫ��L!)%Hc���Si,&+�:�f��RQk4&�!��3E�H��!�lp�f�Y�.�R����ӉZ30���kQ��*&֜�!�k3D� �!�Ѡ�U�h!� МAPx x �;;0�0�;��x���6R�� �Uˡ_�����H0��_��C5-5D�.MV`
t�}>�8~fwff�������ݘ��L�2&�·����� �,�B¤@J8�����N��wW{�f�wxS��`�~��(��i �t��<\dp�_�0������}���t	�~Xz�b��&��Z�D��J���ۘ9��-��<�W����ڝۄ���_e>N�ce
��	[V�g �����rs]U���h�B-��s���,��"�4�D4L���V`	)��H!�hF`W+�u�~�us���������p�m�t4���;M`��S�jT�%��t�2M�;|:������}IBR���9Ӽ՚:Θ�$y�uĺ��FY�ttwc���C�q��J�m���ݛ$��ʋ<�e��|q�J��V�'R:ѣa�o0�	sf��Pc8��c1ևhD�Ymo2�A���]����C ���۳���l�}�᧐E�mo6DD��w�ݶ��tb�f�R顩v�-!��OGQ�Џ���++��GU�*O��"R����m��=<~������a���HuA!���꠭Mi	�c'!�2re��EB��;����,�4�5��%���1�[5��Ы��A{�E؈��x�B)ث�'��⒀`gd��߆fgk��ۘF�M���)�������_.���33<.����w�0�"���ꣽ[�p߶���wWun��I�=�9�6� �V�\dp�;ݗe%BUV���wW�I��2Ǔg7[:q�ΰ�u�b��>a�L�A^�w������Q][��B�Zy�6� �V�\dp��������n�� e��$��4T0U0��έظ��s����$Y��Uۛ��v��mU��x���s����$X:�b�6��*lBWbI���G=��rE�s���k�WԑIQ�pP� �!�w�~R��ʴ�����"� vf|�7T��"��{V`��U�����3��)u�꣋N����2kg`�s��n|�kQ�^���{�'�S/Jv�+Lv��;~���#��{g8ܑ`�H�ݍ�M|����>�8eUW�s����$X:�b���.SN���h���f�=�Y�l$��ݙ�ϖ�\dp�6x�荵t�B�Z|�6S`gӺ� ԩ��g��0�JHI\�w@��M`�݋�l��=�Y�l$���fgN�0�3��3�
�IP�{�>�Vf��k{��SWkv����\ l�χԂEqTes����.��GBe]�[��6�G����<u�I!��Lk��;��w����6�-ع�ݹ�<r����BX�M#��ƶE2�� n(�4���C�{v5-�[p��q���'�;����p��m.v��ӱ/F�<i?k��k뾝�����c�%|��F'-S,A�M��で�NN���*w�����www�ۮ<c��mZ�v9:���綼��R&胟1	�'=��ge�%n��}�V���Nݠ��<Z�G��9�l� ے,�^ظͅ��e
��ؒf��g8}_W�ܑ`����6G����v�oшweZJ��� ے,�[�p�� 罳�n-��-�bJۧi�
�����V�\dp�9�l� ے,�T�M�ٽf��n����u}�o�UJ)���A,;�����n���Q��`gӺ� �K7��߀M��"x�x3���[f[:9�xt]cnp�ק��u�]�qt݀�k�Y�,��f���>��.�����3�@yW?~�몹�����ou0U31/15��Jn]�ކpg����!5(K�������N崋=�Y��;C��7�g�$BYA$QB�]Q���5�X~h$
�)�f����w��T�?3�3�G۫� ���>��H"���z���3�o�w^�� �)� XAٝ��������PK�f����ڸ�����M�J�ZL�9�l�
�"�� ���R�?��������XJ�`j@CF�"fI�N�n����CΫ��7S����gh:���{M���#֮��v��Ak��:
�����.H���Ͼ������t#�d"$A��û��8��O֚hwM	�v��2>�U�$�{ڳ P��wg�q��P.�~���)v���J�u�w��wuq`g��0�lgwq���TjS`{Vȸn��r����:��0*���L30�;;8�;G۫� ���3��S�I0�"�#mXSi+_+O�^�6 ����8�;;��|y.����Ł�{g8�h�U]�;t���Cn��77d�s�S�ca���b@ѵ����Y�Mg��D�,`7C�i�������s������i�*����]U�~�����i��tV$��	�� �}��+��9���<��o��A��J�o����t�1��V�0n����E�r��>68`��1���۬���$0��s��uW��?~�us�o�U��HBY�`jdA	�=@��~���ys��ޭo{ћݛٽkz���s��?$�J�˯�wWf �R��oBb �JM�ml2�g�;r$��7mѓ�^���UpA���U��
�J�Cl�������O �,{ڳ Q�M�s0��;���G��>�,�MҢ��N������p��$� �T�����f����٤;�:a��U0T4TL�Y�tw��`�� ����l���P޳uoe�y��?$#0�g���{������6S`}[L��b�ݦ���p�� �UuUTQ�;n����6}))����7����RR���}v]8v��u��*�ص�en��+<��J���Pv�i_	.y��Gm�GN˜WD��ѭ��7]`�ɮ�C�tYͺ�7ڳ�ƞ9m@���'sѷ���ፐ)]�g�:ݲ6��G&���|m�T�g�ۭ[��خw`��>�+��+�����[b�I��=�;��]�N-��5�B��l����7YL�j��;[j���rM9�
u3����=ws�5��	��&�=��xk��$+T��N�"�c�	�Еؒg@������>�5�]��s��"��_~�����.�y�jx�)�*� �IM��J�8�H�=��fs�C3�33�������RhM�V�mӴ��/���#���g8ܑ`��!�[O���������gfwq��|X�]��Jl?�gwgh��˧ �6�9��X")�虢���՘��f٘�t���?.�8`a�����Wh��p'5�ݜ����C:�==M�MM�f�����^�!���Ճ-�J�i�m�Ω�pJ�ώ�0��Í��ـ��I%��m`��Ω�rU}T�����bU� Q8`�@���� p@N�@﻾��.���vs�m����R���;��y�� ԩ�{Va��ٛ�0�;�������{T�?��6l-,0Lv�UbI��{V`	)�3��S�3���������<��5,<LT1U��Jl� �0w�9�%�X]m�*��QطE����v�f�u�@�����⷇�(��je�UT���4��v2]��[�8ޞ]8�H�=��f���=�RT�AT�QOY7s�jT�wnq��}�� Q��`gҵN�7��M,���L�`{�j�a%66;5����8N�&.b��c�%�&0�M��eQ���Yb9��8�&U�¡�?����_�{������t�5]��wV�%B���6� �Tظ��{��� VȄ�)�mY�3S`gҵN�;;��,����$X$"�j��t�7V���RWK�]M�L#�Q)�W'0�{p�ycmQ��꫾���N�L)ff.�8`�s�m����ݙ�>��t��2�MA*�X�f��g8ܑ`��l���3��@o�]=#5,4T1U���>�%8�H�>�ڳ ��Gd�iK�r�r�%�QAA�C(Hvwwf�l�ߧ �߫�`}��f�fB�"S� <UN��]s]U�������*���������5*E������;4�38�;;�û�n��~����`g���ˏ����`*�)�v���9���R�Ѽ㱷e��6�$FF�ͳ�Ӳ�;t����1&`�s�m�Ω�p�� ٷ{wQ��wV�ҫV�8uIy��wggh�<�pK��}� MB�J|[V[���� �ٕ��gvg���f��2�2h�jXz���h�����	.ư7�ݘ���;?�Gz���6l-*�L��j�Zn�}� �fvn��ޞ]8I[X/�d���ѳ޵e�Q$�iCn��9��Ѿ�4�	���Kz�X7A�ND�i4k{á����.�1Վ�L�e$��bh��5#��V��U�EI[u	���2���D��.�A;@B��M�{����  �p �`$��   r�  �]�֗�8
{v�6�9c�a��@��6�9*T �k%�m8$HHXY�w]���l]s�ܦ͠�r&�{nX����i$�4R@�h  ��-�   #mm�e��t� �� ��m����Y�v�{o\p��R5�mV�jm�T݆Ɨ6d؀��v;F��s;�r�A^�%���v�8,y�qš:q��dTB�=9�U7kWE=j:]e�5�;�6��`-ǲs���g)�v�#�UCZ��]1�秶e���I�j�x	t����:�����m���v�m���}]��;r���96�u[9����W$�I��ί5��W\���a�J��W�ܡ���ʽ�:�����I��* ������+vۤ��N7�:�!1/%�����Dݶ��������@b��P!��˳<���C����1���yV�+�7U�X7W��crsӜbp�j�;�;g�10<vvN�n;]��O%u���zSt6� �G�	q��.Y��
�;5n�6�y\a[ti���mR�*�:eZ�f��h⵵r�9,�P�7�� %55N�0���蹍jJ�����m�m�%�q���q�ʈ⩶^�mt���N�v!�
��7b�
��N�U.��w`���Q�3��I�Ԫ����'\��nlףE�1�5�����V;Y�e�����qq���%۱l�O0:I����X£�q�ݖ�qgv�.�;G��*�˪�Ӯ�tI�9�MZ-nSu�2rN�w:��<oqr�=m�.����1��Us:���m�ٺv���&�Й�s��Zf[xYo<���/NݻC�U����2��SU�*c$�i�mer���F;%�5�㬀C,v䪕n�8۶���H��������=<�\����#�v����;&�{snw�|��s�T�=t6v8*�j�����_��D૆�)�����A�E����-��D��8�ãb�l�&;�1ܼ�+5$����d��s��z�z;p����[���t���X���銈�86��r��ɮۧ�NĻ�M�����n���Ok�ҙ)�⮶9=�Ŭ��_%��A�ٸXv�#ٶ�ph�c��grn�pv�f�m۵�:m=a}Lwn�c�i�u�*�u`�r��:J���k����JT��I�c(�Q!5'���l6�����zY�.�j�Ʋ��A�Y1�ʗ�����ߟ���l���p���gg�y,�=��+t��Ziۦ�Xz���&ɕ`{�%��Jo�ݛ�3����߿IR�SQ2���W8�������j�F�6:�"��ݲ1ҠU`�|�u��U3�����fл����Z� Z����K��F
ګwiU�O�^ȰuzE�&ɕ�w����aeҤ�]�v!�;���]����ӹ@:�-��Y���ܛ�	�O3FU�Yj6�Swv����IoO~~N6L����p	{"�;su��I�N�5�ѝu�Z�}�tu�)��F��6�v�u�f���һŤ� H��� &h�Rq�,�	p��ѹ
���V��0B+�'00LA�3��33?��������K� �j�3��zl-*�L��j�Zn���9�$�Άvh�ӽӀww[X���q����i�K�,�^�p	$��;�I� i�jS�I��&��i5�w��._W�d��;�I�/dX���ۿ,F5�)\��� 3�j�G�W)v3�)�Ӊњh�S�7:�J��z�n� Z���６`
5)�fw����N�d�:�j`����k�y,����ޞ]8���ZF�Ҩ	��ZUj�� ؤ��Sb�*��U/pL��Ɛ��cFM��N�
	��(	�h��r�:
E<D_{��=�꯼���F�b"S�EDEASQa����r��w[X�ڳ o��3�����W�[���Rǘ��e`�s�H���Sb���%]��?[t&�ݻ�m��6�CgR��^5�����nϝN�������qV���P�iՍ7]l��s�H��>��Y��ݟ�;���y���ST1v�e+o�E%�� �&V��Vg������gfi;�5E4�@L�TPT�X��ߧ ԕ��ｫ0R�X�JJ���(�jF�������ve����Wf�R�fvjfwg�����=��Xۥ@��nϚn�w�9�6$��ϥj�RV��ww�]4�!�c�Ǖ�z���9�m�M�)�:um��\Rp�V�4���ڊEUާ��m%.Ei�2f��w���,�RS�jJ�����0������PEAPT�X���?3C��q��gf��߿[X	.���J,ܚ�ZE�I�^<��6I��{����Ix:���I���:`�<��y���Č����}���W?k���9�$\d�X+}���6Qv�e	�p�K�9�$\d�X���85��L�pYl�\�$Hf�b� 3����n�k� ���:Ե[F6�&�ѱ]���a�T�P��rG&
]]t���=�Ƿ���R�8ܓ��kg��<���ڝ��v��v���S�������s�]�R���+]u��,������n��1ȹr�7;��̔u̻�m��9��C��g[�J�M-�u:�H�Y��P�m�ù��܈����="X�%�c�mB��( ��EU�
%T�A Ub����H U!RiCz��4f�fsrS��7Y�<]v�����m�=� �_7 Q��V�63�nK��X�i����� ԕ���{V~ffa�t�E��q�%KTK�UEL�VM����������D �!�}����uO����9�$\��e��T
�v���M`{�՘R�Y��zR�$��|^�}�3Z�Yfk��P�!	H���%IE���wN �V����7w�� nt��T�SQ`}� fg��;3�;wwcX�ݘR�X�����J�c�����'37m�9�����IGƭpOch���As�>��a��m���?��$��=�I�"���I ٲ��Yi\�wb�.�I{������*���W�U�W�!���w�:���5���wW��+ ��뒓�m�]��BO�E%�}))��ݹ�v���������7mJv�իv�PӼ�RE�$�+ ����E%��R!�v�t�4��M�����g{گ �)E��JI�m��{�{�����w�ܙ��Ks�=�{Z+���ඵ]2Y;K��M)z�vt�/��
�v�&�n����Ix:���l�+ ٥�t���He�V$��5JQ|�����;�a�=�����;�������n�r����ݖ�um;�9�$�u}�s��<Y���e$��	�YpR0�A�A^�:맳�b��܋eݫ���+aW�2p?;3����kwWf�R�vfx���Ӏ.]t�,T�U0T�5��{V`ϪR�>T�`���5xm���.nN�n��\d�5��m��3v����gZn��yu�۫�+����nѻUf�R�>T�`���=�j� oz"S�M�[�j����r_?U}�U[3@�u����� �:���L��-Q/TP�3Q�q�j�m`{�՘;7�Һ������b�.�t����Lm��y,�5N��>�RQ�L���fvfkw�ﻛ'=XҎ�M!ݥHM�j�Q`���R�V�k����5��=��h����s�Wfmf�*KM���u�:�w\rs,2ѥ�u�.�y�k���>T�`�[X��g�w�J�=Һ"&&)ƨi�����5j��wga��7uv`�tX� ��Be��]�*۬������;���fV��]Ȇ��;m� vmS�,J��V�kwuf 7})ۦ�V�ڵCN�H������.ưK� �:������fb�J���[����=�������`����2;76�Þ���$�c;j�	�@��f;=v�=o�jQ`�u�F�s��n����z:���j�<+��fz���H��\���ϡm��s�%"l���ͱ��6ѲX����`2��jSv��/F��7#���'N�O �1y��ks�du���r�՘��^v�jtC1;�E�-^���nv����BM�m���ܹ��/�rgu�
mN�9�C]�:��6�Schj��C����|̾�fV��9�6-��rG%��R]��| �nƢ�����Y������.��`}�]рlٕ�l���Q�I�;IU�O�b�%IF�U����� O4&"g���մ���9/�lٕ�n��p��`6-�v�[��t��Z����V�kwuf��M��RS��c�;�K���퇮�m��8��RnA����xl��}pnn��h�k��{���\���p9�
���7wV`T��%<������lGG5SQTEV`Tݻ���S;;?���T|�,�jV��������"S�N�;V��k �RE�6l��7wg8�ذwkc�i����a�&�p9����r�k$�0ۻ��`�H�b�.�t�Ut;�i���� ۛȤ��l�~�7����1$��:i:�h٢�t{����"�9Ϙ֨��뻊����lˤ���<�sb�9�p��n��p��\�Ԫ�m[��X"�.�\� �ݜ�sb���	{~��%iʈ&h.�� մ�}���ə��퓃�c�f�:��S�b�,,o�p�S���~� ��:U+�]ē�ڴ��&n�z4uw�Y�z���I3%4�9�dҘ1
RISH�Df�L�d�n�uGY��E%0JS�%.@U2,�6�����A����=he���h�mڶ�Q�gg�;��H�_00�$ĉ �Ɓ��fm�U�):�K��z�L�CSB����9e)xETY[�� l������܋d�l�
&�P�7`T���TA,A�9a>�O�`FvV���z*�h���F����;�
��آ�$"� &�?21 �"Q	 ����x�!�:S�/`���(&�> N�\@S�?�<A9��>���$^��p��J��;n��J�bL�7۫0��l[IF ����`oͱ
PU5-PIY�}��X�ܯ�>R�,����vHt�TUGbݫ��8˞��\�Z�Lh�Av+��n3q[��a�6k�x��n�*t�jՍ;�������p�'�g*���%����5M"Jj�b�ʸ�=�H�gh��.��~�w\��;��]��|�n�cL��V`l��/���۴�$^�J0IݫUj�� �/ ��%�W�}�]W`��Q�C\����ꏯj��P�[j�4� ��%�
��n�`۳������-Z�F:l��7g����>��)�)Ԛ�n��s��'n��3���)qZ��%y�C���e�n�`۳��0	�r_ ��Q+�l���$�L�'�g8}��ݎ�/�{u� ����)�t�ӱ�8v8X�ԧfx�J��;R����D�����TLLTXs�����]ӀjU��'�g8v8`���5MR�SSe����m`s3��j]��yuq`s�}�k��M@0Ĭ�S�� D����s9��3Y������/%��#��y�x' �Z�V�yYK�W2���ڧ�71����}�k�\�=�+��N��en�ɻE��#��yv���ø��ܼ�sk�<O��4;�v�GN�2��k$nb�V��<�Kr˦�t�+2��]�B��1���9�F�t�
j�;�c�>���k[�'�2��g��g���,�b�e�s�RKMݻw�AG�[��*H�M��F�)���یK�h5�v쓷\v�9eH���e�;~��*̻m��U����u�M��p�p�'Vȸ�fV$/K�	���E�O��2��["�ݙX�����
��r�Ԫ-ն���`�d\۳+ �ݜ���K���i+�1[33 ����'�g8v8`}UD�� �n����ݵJ�7X��� ��uI ����9���Pw�YU��"ۆF㇫s���V��!�Ý�v �L-Ч�o�=dV�$���ک�RS�{u[s;��;�$�0��'1T����TLLTX\�\�5���"e	� Xf�ݝꎮ�kwWf��E��L�����i[8� ����=�l�
���0uI ��vۥ�t�����`��s�wc���%�n̬M/K�	ڧjЋo��0�W���wW�u���y,�%�n���0��F��sU=[��n:����v�zc�poR��]����ظ�mV�m����Z0n�k����wfgw�˫��Q����� �b�	�� �궷g���p�p�9�2ۥD�[n�MTāST���Y�}��g��ݢ>�W��ٕ�N׮��Q�T������ک|�� �궰=�j� o���6�uc�j�l�9�2۳+ ���0�R,fwfn�:\������rp�� %�ڸK@<ɇ����ŷ]sT�ح��}o+1�1|��T%l��t��V�{g8v8e�ɐ�u��St���7wLi��{g8v8`��ٕ�IG����N�-$"�� ��[X�V��%m`{�՘ ��ĴĠx�b����kwwgv��ݜ`�������߹�u��L����4E`d�CA��L5�cP�_�ٝ�U��G��������( ��0�������0{i}�рk�� w�]��+������h(v�����ŷH���������}��qU53v�H�~ {uv`��,�U��;�}�>�B"��mR,CB�8��;�!�;�2���9ͪ���lE$��\%�m%۴�s;�4G����7z��T�i��v�Е�����L����p{\0w\��=u���J�'e1�X}����`�/�w�s���$f�j(���q$j�( �5Ϲ��oV��������<螽�L�vˌ�[q�xjRA�,�5�Sgl��I�p�99�qg�f��ż�nst9�81y�\z'n�:V`A��Ƕn��sā��8�j�H��'��p��ч4&��l`0z�T,��y��`0�:��+0��6�x�w��x���q���j�l���&y�'�s���i��G9��ں�E՘7.�=c��ܲ�'v��mgb�]yNu�ĵ�M�\���:^�^"��T��)���7u� ��%��L��vs�h�P����[c���~T�`y+k�uf�m"��P����LD�E]�`y+k�uf�UW{��0	������*%��v�j��*j�Ùٙ�y.� �UŁ�*J0�L��i��(mU���R���=�p�7��|��+ �ݜ��v����q��S�z��N:;^��`�{(\K�O�h�f���t�֊痷FT+}���%��L��vs�{�e�HF;�wI˂��{x�%����%QTiEU����G���ޝQ`oʒ���؅#��*N�cN�M���-��껞����m`$!�*jf�&dj�����]�Wt`y+k�uf )��$� ��hwi;�7��|��+ �ݜ���x�W����V�4�]u�x99�����y{�I�ʘ�V�0��A;�g8%��cYwi+� b�o3/�w�e`����[/ ��%���⶝�ڡ+���vs�{�e����I������P���&�J�� �S���s�]�T�?�B��f�Cڜs0�01�2�6�ֵl6%)�I�@41l�J#Uo ��5�$33�;��<]ou���-����DUM2�@;VӼ{&C�w�e`����[/ �T�i���;���k�p����庳 ��TX�V��������)��ݞns�]�lp�m����Ќ`6�r��6N�L���֋���$�M6��f�N��7��J��M+�ԃ�M*iXSi�{�e�����'�����m`yn���&ZfSIT��N���I��zn�pyl��"ۻI\��v�
���I�`yn��=������X�چSm;lnĬn�M���-��od�p�L�g��"�m��t|�O�q��ۚ�a���vہ�t���-�v#���#��;��:i����Г|���x�L� ���=7g8�{b��l��J�w�od�p�L��vs�{�e�l�m�����6�� ���=7g8��^��!�=u�v�O�Ɲ`����[/ �ɐ���X�����iU۠��� ����7��J����Y�|������O�Q�kH� )�Jϳ%��I�8儞	�&�-��7������Pu��6�1BN��5�%!�DjB����02����Ѻw�]��E�R��"�1��*�d����X�@h���������"��׳A�IGę5D=6��(f0��f #���:��c�8k���ی:1��1@���LN�@�T��$t�
Z!���@[5a�溼-Ovȋ���r2L`huٚ��B����cV6!���I& R�?'�6�wwwwwv �p ��8��   �   J������K�e��sv�V^�٨-��5�K�:5U���LH�mY-x4�:m,�f㦲�7m�&�m��<u�v��r�7L�M���6�8 �m  �[[l    $m��,��q�Ѓ��m�� h]ni��T�oUT�3�7m%S��q����@�ҽQ��6^�m�br�jLP\;�x	5�:��Rni^^N��qی�H�'@�k�;�c;N��Z��l��X�x�[��d'88S�)���OON�� \ut�Fk�3���Iؘ�Ug�28���3��lTۓV����[7o]��ѹ�.���pl�Q΍t�ե�I��sS۷+�.��-�`G�����֢��!��g:�=ɑ�+�P�L#�vI��+j�����cפ ) �v��n۪�#��Q� ;L2����
�me��Uk��f�ѫ����F�zl�(9��^u��N��4�.1�gO�� �
�bA��AN���ȡ��Z�r5���v�H.o*\��(ӎ�����_=uV����k��݁jP�k�u���ɫ<
����TA��K`s. ��vl;-��C���c��֌�rΛr� d)ӄ��1�F��i�Xpݨg�G㇄l���pUUX�U=.�,��&�Ql�U��l��z��>]���ZĮ���
���-[,&_5��͞b9�`9H����`d��8k���+�lp�m��4f4Σh�d�ę�]���2&9ܞ8؛��3�p�����6vE��Ai����ى����V�^������uú�.���6�c�v���<Ѽmcl��s��ym�b�Tw3]N�vأ�5[Ecgs���2�7�^4u�Q��vC�]n�X6�V-jՠr�vf�6��Ij�.�c����m�ͺ�VS��<{,���n`�۷e˥�ts���S��k�(����{wCF��K& ����w���������=��F�+�g_Y��`�j�SWG��%��� ;���ډ`����2��(���ɹ�T��)ʢՍI'%'Q�!�J�Rv�qS��ly)6�:m���p][�������.�eɚ�SP�F��Sr�5�=pnDd�W0p�C0�Zn�ud��klgs��(!��]�\�vx#k��Ü��}�i�x-
�N\�:�=�v�%]���ݹz��='\�+�Z�ܻj������n� ��6b�Y�q�W'C��(�E�/:�`':�����79���.^V�]B/+F�%m`yn��=�J,�������aV�a�=�2�M���)/ �ɐ�ꪻ7~��bN�M�e�ST��]��)E��%h�=䭬V��*�_]�4Z���=�%��2ޓ+ �ݜ�u�jۢ�(`��w�od�p{fV�9�;�%��hU�`*��i�N�bI��C�a�\n_h�H���ɐ:��ʆ�<��жNI���B����c\À{�2�n�� �od�p�z]�;LaI)�:�=Ͼ�}�S��$"�CpHdH�\Fq�p!I��1�011&H�@�U�^[/ ���p�fV W���iYn��O��R^��!�=�X��� ڹ{IRJP�He�� �ɐ��̬ۻ9�=��\���Y����8}&V�s�{�e��2 �z��V��7V w+Us�\��]Q��6�ͫG�/\���b�v�ݳ�i�M�e�`�u�{d����l��I��r�ޡ�n��!��O��R^�!�=�2�l��n��[e;wC��� �ɐ���X~��M�%0X��I��C8øó�0�U���7etX	{UTK������S�`s�;3Ƿ����ـ{Ӫ,9ٚ5wg�j��*&�ի)���`�'8��^�!�;�2��6�Qwwl�ڶ�-��*�u� v�WM���U����4�<K��$�<z:�l����SM�{�K�=��|ޓ+ ��9�6�^�T��촇v���Q����{{��]ݘ�:���%&جR�;`]�e��L��ݜ��ٝݙ�7g�,�Wt`�M��MMT�-+���ݜ��"�9�r_���>�_}��uW�=ϵj���Z�ВO� �G�{T�p	$��=�Np	~��ۺAnۺ-��a�M=�j�+Z�@\�נ�wK�[����]s��7Βc�j�	5m��RE�$�+ ��9�	$xٱ�ؾ��	&s. �V��%� �U`z5%X�-�Hv��c
�'X�I� I#�=sd|I2����R
�4���SM�	%Vޕ)V �V����{��U��IRK��;-!�m��6G�$J���$� J�g�d�40��'u��,���K��,]�m@	�1��7� +���%en��+6�����O9hݝh���9��:e�nͭ�<�Vݝ����1�zϗ�mk�l�,\[vv�����)�3K���{(y�x��ݘ�؈�vm���?}�vv�w'C�;���9�tM�sf��74=J�.LN8fx�f��c�|��a���c�5�.
���Q��T��V.W�ϋ����j}��r��"y+���y�<ݖ�@�2�ɕM�.;d�y��U���0Rq���ɟ��֊��������%� �U`z���H�����uh��� �I9���е*�J��3;4A�wDsI�TA�RL��`wuX��V �V��I��^؆����j�x�l��I&V��s�H�	�bm�OQ-LD�V\�� �V��-�� ���u)��82�"$���&*��֗ó�b]uX�]�����n�2��&L4��y;�v¬I���s�H�_���I&Vߧ޽��M*�t����W9�o�	��$�sOቄ06��s#�,Q5c&CS�1$@RA:�fq��Z0���&�MjbgZ&pM���Jl��4J���c������!��0SZ��!�^ '�^b���9r��=�`УZe�e5DD�SQUV��(�J��x���� ��Д��)�
*("��� I+k�If�$�X� Iқ���M˫E��`��� �G�z����e`�ڸX��%�$�i�7�/��]���刺$�f�N�y��9M[���R���HubZ�դ�� $��ݙ$�XvI��^؆����j�x�l��I&Vݒs�H�	�bm�e;Ut贙ǘ��e`�';�4�B����#, `�.R��8d�����B$2��)�`�RKUW�Va$��&�"�u�dC����(	�kgwx������l�S�I&V�>��BiSJo� �*�=�IF �V�ڒ���#�i��o��h�S4��"��<��
Ĭ89�qf:���^����6��b���R�� I+k�jY�����@��`z�DK��]�l,O0�I��Wg�L�	$x}�Lw�Ֆ�ؚ-�V�i��;�'8$� �d8�e`���"X���hI�H��U� I+kfwf�fw�y�u}��{bi�;Wnƚ���ِ�I��wvNpI�x��%���v��w��V�{��=�$�i��3��9��zq�[�8����i�I��Uc�`贘�0�I��wvNpI�ِ���D6���[�����>�K0w$���R�`	%��o��\��M*iXSm�H��$�X�d� ڹ{IRJ2�,Hi�o ��%�	$��=�'8Ē<�"��j�WE1�f_ �L�۲s�H��r_ &�Ʈ�V�}8M�Y����5�rc�t!�R���R�P�Jj%O`.P��2t�<�u���%�g���ۏn�u��;Ƣ]��M��vK��;��H����n��3�(��A��pK��w-�u	<Hc�+�m�=pkh6 �c�٬v5��W&G��{$���t.����ŞP�u���5��ڝ_�����n�����6�G%�#��uӒ����O�|�����]�݄�hq��q�6ֹ�=�k�'NS=̜�_s��z���qc�]���������IݎK�I��r�ޥu*�n��6$�|��<�;��|I2�n���^؆�i��V��V��;��|I2�n�� I#�'���k�ݴ��M�X�$� $��zL� 4��!��t�ݕe�X��� KUX�V�-V���3�/o���mоYg��8�)z8Q3�
眴�/Vq�wL9n��q��[=����j� KUX�V�-V����Z%�J������m�ޓ!˯�����/"T��y%� ��������R�bc���j�*���u���$� $��zL� ��Yc�J�.�橬y%� �U`{�Z0I+k�n��e7wj�4��� I#�?n����;�[X�K0�j%�!�5$�L�g������q��ѺK[�["�\��x�=QE�C���Cm;L,M�m�ޓ!�$ٕ�{�NpM� ��m��V[@�c|ÀI�+(zI� I���V��ggx�F�%T��P44�U�߿~ﺮs�o��Ba2�Iܿ��X���$��fca���	��,K�Z���i
�,0��b�f f^!]����v��=�AN��&�(3P�46@("��9r
�;�NZHe'P*���I�0�J����LH��f�F4l7��K�����kF�t	�: �����4i��HRR ���6�:ηխ��kZb�K"0�QD�����YkTf��YZ�F�n�4)��$l�M��ɦ�,�͉��]bQ@�e t���	�:�M��deFf84�+
hA�EKH��C�@:�؀�����](��'N�_z�S�@�`r�����s� �L�~�z�B�e�YI7� ���=�Z����Y�kD�I!+�`ZJ�v��=�2M�V��� KUX���ɡ�#����j9��3>�Nd`�ח�$��ϝ���y;vH'udw�'ְ��X��ݼà~�?e`�'8$� �ِ�VŔ���2��m�X�I�$� �ِ�I��rK�B%YI�ڧM�i�H�I2I2��'8�n�4մ�V�j�x��.$�X쓜U}u������mU�hM�<�RV�3;��� ]�V�a�]��~��������Sn����͑Ѯ�.6�ew]a�v�W�j��= �;t(\%�ɺ�=k:�4�SWue�X�'8�G�l�K�$��;��� *�-�ʴ�8�J�����@.��wu���%��(��-\�EZJ�o ���6I��l�s�$xūA���.�M�����5%m`y$� 5%Vn�J0	^ٌV���.��u�zI9��<v9/�l�+ t�磌݅쫻k] /E��9֢�b�:\d:6+��Ԡ,�_c"�]׎��f*4 �vv�n����.�$�]v�oK�8������L�n�y�!� ��ԁf��x���np!��=_�c�ew
�{WNR,�rUj��&2n2v�LY�5��h؅|ܻ�/f`����2�dv�,Y����3�!��^��q�ShG��EwjӖ�������)�I<Q�V���=r�|��j�a�ύ=�������#Zy̏kW0=]&딸�p=t�o��m���X�Z0I[XI,�6uISSm:��ڴ��&C�I&V�$� $���I�m�eڲ�	&��-V��K0-U`n�h�4Q7v?�5wV$� ��s�lx�&̬�O�{P��mU���	j��:K����]m`|�Y�߿��s�����r�w������\�m]�^5�iCP��N�jZk��]�qۑuMD�X��Z���K9������uX�J
"g�"!�� ��0��G[6y",BI(�1��3���3;=�KVf -J�n�FT^ٌV��.��u�wd����ِ�l��7�*!�c"%��d����gg���R�� I+��$� ۯl��vӡZhm�m��V���$���%� �U`}�cc�������Ӹ��Cl.��Su��M�㸲���<]r�i������3�`	%m`}��`IW;�@y.�0wIU4�S�T�44�۩fs33�@wwU����J��ٙ� �A�.
bb(����� ����j���D�U$��/p�2Iܬ��9�6�^�H�R��V�ӊ���vvh�]�`���۩f;��GwuX���@�R1Wf �V�۩f $�Xn�F����I�ԗWڜzS�{qsF�j��.3��͖�wf��@�x�9��ܭfv�q4���� I*�>�V�ffv������ۯ�G�)�-S��i�H��̇ �L���s�m׶Ri�i��v4ն��̇ �L���s�H�	&��k故����|ÀI&V��Y�	%V�ό����� �E�uc�1V$� ����<��!�$�+ �����ʻ�wm[Mʾi��-����ž��:�*f[gv�w\�8��E��ҡ:���� I#�;�2I2�����r��E�R���14��ِ��2����ے,dkA�nXbh��pݙXwd� ���ِ��GM�����5M`}��`BJl�U����%���vm��#���uj�|��"�3uZ0�V�ۺ� ��Q	@DTJUU����`-�F0 �N��`A�������!��n�v:ON��Q�\�
��N=r6�!z�"��[�ڸ����G�a�� tt��kt�d��s���n��حqv�s/gG'AĻ�V�x�� �؍
���f��7S����q�n�pxv��S��B�����Ͳ�*�p��-�F��ڌݧd��Q�
��'���j�wyc�gi���A�xIh*�y.�����Ճ���f�vtUN�*I�i�&]����k�zO����2���� ��$�����`�i+v�� �ٕ�wwg8nH�ṅ <BD�V���]X����9�}	)�3uZ0�V��C�j
a]��Օm>pܑ`ݙ��+ ���p���hWjRZCM`ݙ��+ ���pܑ`���T�C��tql�]�pt�ێ���	��������� �㳏����x��������+ ���pܑ`ݙ��q��wM[n'r�ė}�ߛ���PW���vz1)�7R�`����C)$PR)ة��M�v� �ِ��2�	����^��lI��v44��'vd8�̬{vs�v�E�l�6�_4�خ�M[�۳+ ��9�;{"�'d�py��.�j�%m��ixL�*F��ݜb�R4u])&���ݜ��m:�e7H��'X�����;&C��������WV�ՑQ5�ѻ���-�m`-�Y����К$��x
&J&*���w_��tu
�
��R��Z!�g�֦gf�;������Ԧ��Pv�V���y� ����&��p�R�ggx�wgm�ꪩ�b�
��V��&��p�Ȱ	���ٝ�������e~�)���Ի��	.�����D2�Y��m��B�j74���,`�M��7���;��=�2�	���n�)(�i2ڧcC��;��=�2�	�����,�H�l_9
����'.� �궰�Y�3��zt������T�L�QM$�4��՘�*��%8�L����4;�]Ww�`&�Do�A$TMf jJ���N�+k-՘���`����i�ўN�W�L�F�.��:ݫ��u��\9�N����.�L�M�� l���q�˷,��y��l�+ �vs�$x��.+u��HVꭗt��m`%�� 5%VS� ԕ����Z��ϛ��M��7�D�<O9/�$���;��4w%�`
y�z�����M5m�E� �L�M�� Ns���C���
`�F����'�6 b�9	�SF��h�4A�1��5�0щHHs	@��,&�eY����*��ED:��j��&F�`$��)��1$d`["ޚ�R��4(�A���̄titF��q,��j$�{�Y�7Ѩ! ����1с.�6f&����kZd2��{�{�,խo0g&tmؐ�I ���H� �b!�N��8�bF2���Bcj2SPQM�fɊ4�L�M���EQN����荐�# �'0,HR� ��( �Z��� (�(a`"�,�
�kƲH!6Z��{�HúBB�� HCBP%H�@T$��	B5#$�AaA8L۪�"B��2kv j��0c�פ�{�N���w{��~��   I�����    oP   7N�f^�N�f����۶���z�,�;줻��"��yڀ��j䰉i�\��ZH�+�3q��%�f�>q>gd�Fk2��H��Z�m �m ��mm�    Y����q2��T�UUU!®ghq,J��dS�ⶸ���
�LjQ����ʆ���umI8n6�*��ٰ����
�:��l����=@q�� ��;y�ܛ����f67`��l!�' �:܌9܎۷l��n:�g���>�[k)��Ad�v����5�E�v'+8�A�]���{v7�{U��Cc3rμ�5`� �8�&��:2-Aۜ�	nv�c�s��3����mV�3�4���ї����=��m�٦V�OS^��k��6pS�]6�h��紮��	&6R�A�+��!+�Z.��.%��2�UX&��n�htu��WLq\��B=t6��/q�Nܙ�c�׋Y���!����Js�켯R��l����^ۗ-��7 ��C�2�Ի��hN��tm������8����23V���̻���1�Iےtºh$��J�|�+��]�/$�0h`1�a��mUR��;� *��S�x�g����6���R[i�jU�M��ҾZ��؝����x&:<UV���㥩�,�V�u�6t��	k��'D�ReskJ-�:W�ԥVIu�l�T�]\�	bF�5�/=Ümnȑ��۱v�V;1m�m�!�^�W���K<�/*�h�r�m|I�K����+;�#�n��;X��]�m&7�yz1d�e�q��-I����ln�d젏G{^1u����=z͔��]�
�nb�̼jv'��嚺�#��{q�ؚ��O!/ъ���8(���� 6��yx�a��E�v~���}���>�����n��^7a�u-��WJ^�m���V6ޱ�?p}V����Eغ՝��:�;���L�L��%�!��wwww�=T���U�@~����P�@��>(��C�F��{�����߻�?�?�A4�UAx9h.v9=�z�x<ƈ)j�孞VR�B��8��b籱k�q����sN�O�k���Onƞ��qvպ�nnҿ�o��R�d*m��[�[��``:�w^t�;&�[�F���=� ��	UƸ"��ܴ���z�w��f:P��G�'K�דeܠk`.�k��8wCځN����-�ݪq��6�GFqv5C`�-��w����v�@Y5'\��s�{�8ԓ6^Oi���n�=:�k�"*�\ӭ:M�D�KD��� ������� JG�I�����n��c�*�'V^՘ �U`%�J0���5�x��N�n��>pI'���I��I��W/jЮԤP�����	<�_ �L�Ol� $���q�˶O�Ӻ.�<�$�X��� I#�$��|�n��w1�;n���A�v��9� ��&{G]�ڦ.wS�"��d����`�]�]6�n�J�Re�+v�p߶~� $���Z��fv�wu����e3@�Q�U����<O=��6I��I�Y����CoI<�LMEL�ISSU`wmwF�J��Kuf {R��%UT��TS�j�3/�{d��$ݜ��G�I�%�O7n�%v�HT��X	n��jU`%�J0I[Xo$�콿�1�J��;��w)Z���W!K���y/s��ks����
ۮ��X�Q5��*��%����V`�^ա\N�Bv��$��ĭ��V`����� �:�����v��b"n�0���[�0ְfk�fl("4�	��U!�ff����J%�Bс�_}_Wn���$� �G���덻i+uI�t��� �vs�$x�r_ �&V;�+%��]�M����U���ݷ� ����Kuf�:D�~e�(c˻M/h��.����-�5��G%�:�Wbŀ����dy��db^�2M�y�|d�X��� �#�=$��Ք���LO�p�e`n�pd� ��!�=.7j�$5n�UbN�	7g8$� ��!�7d��6����4����i��<Oy�.����.��"��a�����$|� �^�ա\N�Bv���`J�`%�� 7R�ϾKp?�u1�M�S���KC�a�zv1�u.q��c�As�.w�Vo�ű|����}�X=#�&�� 7dx�����m4���˺Um3 �vs��<OL� �'��+%��]�M�� 7R�/+F������;���=u�)�Ӷ�44ն�	=2H�I�9�	$x���ڦ� t�Zb|ÀI0	7g8$� ��!�6��e�cCm�m���N�k��p�5Fs��$��\��) 5���})\ea�����5t��a�����k@y�`5��������|]��]-F�Skxñf��=B�Z�xwS����:�%�g.r�u�@��d'�;��mZ��h��+�U�::�q��P�'V�	��{��Aɣm�Y�9��;������'�1و}q�M
�W��v��Fy����@M����n�瓏.vcl�l�9t/9��S�B��=�͹�k1Q�����	�0�0$��K���ٝ�������M�lGsM5R4TMf $�_3�ܯ�����j�ZmZ#I�P������L� �8`�g8$� ��[qV�n��%H�<���IU�33�%�8��F�6�J�Re�+v��zM������� K��jT�/���\�n�<\�^{7&���lw�mɭ���6^�{7��͘� �x���\�F�_���G�n��p�� ��9�6��
S�n���o �c�.��}_PUW]���vv{wk�R��<�f jJ�	$����+Jժ��p�� �3ggx�wuX�Xl6�AU065e�� �鳜 �#�=���;�ܬe����I��Um>p�#�9ݷ��0j�Xr՘����kR�	�N���Q!�^Ż-�cf�Fض3�팓^� V殺t�h�>�~��E�wu�rM��� ��al-�G֝�cX��p�9&�pvG�z���y�m[I:�˺T�f'�s�����W�p�*2D��$�R��_g��]U�o몧�V�W(wL�t�M��<|���wu�I�9�6�ڈ�+n�h��j���z��9����� ����ԫ��̻�8��o��bh���j��8�̃�,�y�x�L��`�p�g��s5�ɦ�k�n�I	 �w�?O��I�/� �#�7V��}ۭnݴ�n�H��0	='86G�o�����0�K�J�tݠ�v�86G�o�����0	='8��ں���Bn��O�,�֖^K01�wvv�Z���"��	�UZw@c��c�'�� &����� {�^��j�[��Ή|H[;���;M����,���$�v^)Gk�ꕴ�V�'Ul��ę�I�9�	�<o�Հo��M�Z�\��2��h-7� M��~��}�LOI�.���b��ڦ��[o ���`�z`zNpl� ��6�H�E�r�\lp�$������j�6��Zݻi&4�M6`zNpjU`l{�6�kK�wu���U��M]�(��g���j:]��*�0ث�=���r�;���jd�dIۯ�M��u���%<m�qɮ{]�j6�pO�Nm���D�	y�./���G��짋s�zy
ݺN;4��X�]N4�9��iZcQ��j�h�i�қ���[CۏO]�v��냳�a��N�Y��m��h$G6���u����[������ǽ���}�V�U!�Fl��{X�c��ݎ�;J��Y����eV��+�ݧeӦ� �ô������6��X�^����,$R��iۡ	��m�`�z`M��Ԫ�;�A�;���+�F��`����W^K0�*�6=���T�T�m:���LI���� ���~���צ;�jUr�t˷I���8�#�6��X��LOI�u����v�j(ؠ@�(��Ȱ��Ckk���=��F;C��Z���լ���������� ��� �n�����!q��V�˹�/Ͽ/�c�U"���"M�� &���{V�ݺ���H�1�WM6`zNpl� �/m��z`]�t鴨�i>p?}T�˺���,�֖/%��Q�j�t*o �/m��z`zNpl� �{K-R�Wq�HwV��f�4�Tpk��q[��Z:����zn���rl>;`�"�'t;�w�&�l�� M����k�k[V]�����ę�M�9�	�<ڽ��o��Nµ*�C�U�&��|���^�������lK �[&��,���e�=h@�t�;gN�N��޵�{4��]w�$x��h�o:�-nK��f����y�:�zӡƕ2d�iNsC+S��O�"�aI#:��8A�%Z� -c�E��d2f6lz��0Ѿ�z�2""cDeA�"h���,���2lȍ@i+y���$�䁝F͘d0AI@�&!')�T�!$p�1�X�V�@��j��9��͡m�C�V<:�#i�$��2�ѭ:�ғmsF�4#�2�:C�2Єs�n⊱R4�"Q4�E�1d�&X�e�:��rČ��Dʽ7��Qd�VT�C,а��dfU`cCF�$����7Q��X%��e�1��3E���+������Γ&f�:R`#0s�bB���� �0M�MԦ^��NΓ��1� ؈��CBx�y�d �> /������ =Qa �n�۽}0	�l� �^�F1[�v�m�����o��M�����$m�t�Ҳ�]�w��M��I� M�����E��+Ywt��)Y����'d���e�׬ph�OUl!�U�\�7V�$��nݴ�6Z�vـM�����^��;���=]�t鴨�v�8�#�=�v��0	�Np���n�T*o ����;���]��9��4$�l�!	������ �$� 7dxT|)(R�) B�LBL����*& 	ַ�_gU|{�-iYv�b��4��M�s��<vwb��v��?;��y�Z8�f"N����Gm�b2�BrX�>��
�=�����זF��"�LV;e[Bh-7ހI���7gv,�kNgf����Cj���b�n���[o �[��wu�I$� 7dx����ҧJ���Ě��� �I� n��wu�}ۭnݴ�X�n�m��NpvG��� ��� �mٱP�ҡ?�i��U�n�Ձ��i`$��Y�ٙ�h~�
��Em3MA���v��;q�J��EB�<�J�!�b8ˮ���#j���ѽ�-��أ��s�N{ub��>9�[��y]�'v�q�-J��J]WNp���n��=�Q���tnV�l��j}���&��c�E�v��e���,�4������u7�b�[���
��v���n�8N�h\�Jv�)^x�ӘͫKඵ�:���j��9{��fn���ۍ��uCָy}p�P���%�;���X�:��O뤂Ӧ���
�N���� ��� �6NpvG�M	0nƥ"���.� ��'8�dX�ݫ����ʩ�"%�%�d���;�w8o� o�^��r�	�Q�%V�U�&��|��lX��x;���$�9�=u6�;b�CN���׀s�ܬM���� �-PA���es��x0�Qڌn��;Xs�ba:;Q9���+�uL�%�.���������k-K0�ڧ��� �U����m 6[�v�`���:��W�Q�H�,���'�Y��ݮ�F�M�/yU�}����D���*�v�8o�, �n� �}� �d� �^�즛��
�M+M`�u�{�x�'8o�,hI�wmJE![��| ��<M���� o�^߽^�������hm���3�8�&|]�ٞ:��v�*�퇔�Jc�����O������b�zbX��b����ـ}Jl}�����n�^�ule�*h-7�В� �nՀ{�ڰԳ �d���[����X��x�{^>���"����X���a�ٝ�Z�J�f����F���t��ݺ�k������vNpܑ`_}�ߤ� �캍ۻj�Se�CM��d� ��E��׀���9_��m��}��2Y���!�J�Ǆc;����� ��m';���gug��fqmC�O��|��H�}����x���U��)��B�SI&���y���� =������=Jl�+&�*U!�����H�	퓜�� wۯ �u{[E���Ш�C��=���W����U^{���PJ�)T��A߈��u�|����Q���2݂݊M�z��`}����x����Qu{u��8㝩ɒ$�*�]�8�ng'D��E/j��3��X���]�m�:�6�%�q��������`{���'�Np_�X�H�n�[��I5��| ��x��� {�< �^���kv�ڰT�n��x��� zlxw^�����f�EKN5���������`���?I'8��rSMӶ
�N�M�����u�I9�I����x��UUk��,��a����Š�����\��;ƴ]��󵷍�8�޴{p��:��xgl�.zƛ�˞mXg���i�V����sXH�;�-����Y�ݼDc�CDi�1(/lk�<��Ů����l���;.�M�aӸ���:]ݶt�s�0p����}�^.�(�iנ������غův�L+Ҍ�s�yÖ��=�w{�{�\�[�e��;]t���):�m�-Y��!ػ����)t�pKsl�ΣO��8����'��	$���#�7u�v�������C��$�� ����z`���	���+�c��J݂m� y%V�֖�nՀ�K0��&��
���x��UUU�2�#�?I'8�#�6i���Һ[����� n��	$���� �[����;��߾��Rn�=�r�r!�ݝ8�o,vl�Ż#���'v��N���0O]*`���x�'8�#�7���{u��ݛn�lT'�4��I*�ݾfwfy��,��-K0��rU�ؐ]
��m��z`}��	6Np�#�$	+C�B)[
"���gwgh�]�`w.��n��7���=]^��e��ҫ��7�I�f���u`U"�3۵`w�e'~N�M�[=s�w=tl�+jwr�s��v�Z�3���d`ͨ��v�[G\�����lx�^���M��n��M1��v����[�����$�9�{c�6CcMWO�t�Vq;��y��W9�9�w��uҨ��]]-� ޯm��m��wmU�c�[��=$� =� ����;���n͈�C�*��� {��-��wu��Np�:_\b�e�ccd��ۜ����%Ζ^�,�Ð،v�����aiն�h.���M��x���I� {��V6�I]+`��8�H��'8�lx��k���"�_:Uul����'8�lx}���HQr"���:�v]���{c�;���wu�d��l��"��%�J!" L�T�n��{�Yn����	IX666$���F�BT��f�`�%h��ӼŬ���͛�%"f$�Zv��DTT��)S0lF&���0����oZ�=�a�9&��
�;N�o ���wu��'8�H�	6�/K(U-�i�I�Xh��m�T�+��Ayu�8�Ӧ�:�f��3i����E��.3�� �����#�;�8`��Ѵ˶Z)�����1y,�wgx����޶��ݫL���}�D�E1QD�4�5���V�y[X�nՁ��f��DMS.�]��m��V w�� �����#�7BJ���;�RL)5��y*�/������x.�>��`s���o�f�
�����TW����@EU?����]�{�u��Pw*������0 2D�h�
".J�+M !����R�@�@��ւ�/��APj��*�������������O��	����G�w���߿�X~_���������?�������	��?���AU��?��g�����������?�`T?���^`���?�����?���?�'��h�
������3�������:�����s��MD��aI��c��������T�x� � 
�%*% ��  ���C*$) ��HHBHJ�B2�!
�@��*��HB�! ��HB�� @BHB�*�H,!� HH� H�!
�!��"�� B�!��B"HB� JHH�B��J J�! $�$
��@J��*� B0��@@��J	��2�@�
���"�B�$!")��",� ��
���(H� 2�J�!"�
����$��B�� H ��  ����"! JB) JHJ� H)@� H�@� J+JB B�! �� 2��2� @�B @�"�(�"����#(� H�@����
��) �2� H�� J2�� H�,+ J�! �2�!�2(H2���`�����2�J��"�2�J00�����0����J2�JH0��(��2��#��0�# H0���B2�� �H0ʀ�, C�(( R��$(D�D�D LK($"��5�������Ҋ����o���W��G�)��������UU����?��Fo�t���y����3�q��?�UU����`�Y�<7���� ����*����������U_��{뭠�������?��oa���y�n?�ogA�v*����q��������UU��o�d��������0��:��
��������������G�E>�hYv������߁�����N�PU^�
�O�d?����{$���?���������UTW�C����?��TW/������������R�����PVI��t?O f�V` ������_���
AE **�@I%��(�E";4":7F�T� �R
���    �R�
�"�AD����BU
 �H (� �R�  QHUJ��   Z�  (  
�  �^�!��b�� ΃;w�-P�B����ށ���^h :���0m�� �����Mu�� t�ۺ��@������,`�n3�@"���@@ �.L i��Y���>�E�,���t��  X���4��(R��(�$ =�� 	��  �4裉�� z�JP1 ҔbPh����{: ��
�(�@���@ i�'`t� ,�  (( �8�)�OF{= )W>ˋNZ�YjK�����68��I�s��ܚ���咫� u�o�sd�� .��`t�=�ֻ� <�INX�Ye͗,����N�� ��c}�N0��q�KRw�ϐ�  *��h��R3k����m9e]>���� O>*��ڗ�ڹ�]��|���'ݓ��|H ���m|���[���
1jS�� )��^�#)d3���W �T  (((�(<�j��5�>�r��@�D�z�\�Ns�;����v���$� e�-C}  ��0<��\Y.g ��( æ&�c���۽�rO�    =F�̔�   �	%T ��Ǫ�%=D�  '�U%=�)��F LES�Д�U)J�  E4CRRH��0���%W�/��Q�U�����3)V(�ǘ��(Q	D+�]��"(*������"(*��DPU�AU��(�~#��F?���p�M2���!rf����������[{�9�U2���e�O���O��]��+އ�_}�W6!���,@�H�<���6���#@��%�Ө�0e���X�`K3lÒq��Y�`|`�8M�>bH�	����dH1�!�I����b2$ؖHY>&��}iB�I�!$�!��_cI�Hb�b�W�`� �#�'��r����}��<���d<K\���Y���}�xa$�� �
�$�
Ū#*D�1!�&�l�e��w�>���^��R����W�M���׃Ǘ���Æ��_X�{���KҼp�+1�u]���%j�wG��Lu��9���%׳�о��3;(m��@�2�9.���8l��7,��Hc�O{;j.뗾�������p���0�O��]��i�d.�37p�g����CH-�4t���m~+��z|�x=0���6�ᰰh���!�R�4�j�p�����;)�,~~��˄��z�0��"�=��OK���y�{����L��L�^���A$�,�_!a��Fi�U�K7����b��ᐢ�\�������]~}���/����s��S8a�3}�ge�X�d�v_c�G�X4A!�X��=��T[Ǭ�uu|����n���P�TS4����W�
��`x�H	B�0�I-
>�46��i�P^��,2��-�\'<�a�V!E�P�	e$@d
�"$��	)����5fhq=Û=<�F��쾱�D�����7;�Xx��Ǟ<Z8�*{
�P���o��X��@�U��=��X;(L�&Uݛ�:_�3�ѕ����kɪH4�Lj�*tL���6Yʂ�����)wi�=���Q�͗ͮV�׊3Y���d�����^dN9C(���^> �kCZT+�w�l�&B8�|Y���@>P8D�.�-"D"I,RP�GF��4ӛ�du�x��̳�5-YU]�GZu�=�K��I��A����f�ڤJ�f�,bi`]&��!�:x8S3\q��jF��f�SS�M�6�W�e?l��9R��3'OOM�Ga����{�ڣEkQbh�j�Ǩi06�F�M�@�*/��L�--�āi�6$��2W��4��! �j@a"Ak�~�XoR�B%4XR͆�Hl�%#D�aH]f1����f0� Z�iaau��7Fl�V�X�Yw�B֙C�!���£�!�2f[#�S8�B�x77D�E�Fc5�X��Gd*�c�@�H4�`D�H0�����I!L��<3��앯3�Z����/����������ᇏ��i�
�A�@�!aK# �1B�ȃ �D &�6+k�ÎL"0�a�?z�w~d�.n �4߮U�;~����y�\�qɮgi�����:~u�f\�I�\�r�i��G�CU<��o�e9y{f���ʼ��7f3�dN��2a���0���,�g��D�c"�!`"P�!O!��}����!V�oC�!�1�E���J�q�T�T�<OO��g�
��l=]�)�`o�"�ּ_o�\6<L���;o�7p��Y��j��i~sI��p�{1��%��`$ZȗϞ1��XCT-w�q�d7<yba
/3z_��ȇ%vn�<�{�$�W�mUm��\}ݾ�ל��xᙦ�}��QOB��,X�m�!��k�w|�@���J'�,0	S������	���k�s�c=�vx�����K��]&ɽ��X3c#�ץ��h_�6�ݜ���^7��c%f����\P�xQf���{L]�x���!���))�c��%�mH�B�n�l��}�5(�{�Ҿ��ϫ��yq�CXaI4���S[	u��4s��b%d�y��}YU�J��L��,wu���d){&��:�&�*��Cc>BB+F����پ�h2%�͘p�<|#Gc�O�1�.�KX�q�0��^O��_}����3Ӿ�u*����᱅-\p��$��H�y�SR���6MzÇĂ��JW6i &҄\�f��-�w�ȞSy�5�>�j����3;=^zD5�/t��^���F�Y��&� R-&EI��e���g���!���w����lٔy�WS{1snU��1���ˬާ&����5ЁDҌJ��A"�8�lX��7��@�)��l��%K&n��p��Jp�d�!�9P�zs�V�
���0ф���� �T C�T��綥$ �� !	n��=��@N>O��� HB(Q�$bU�|s^y�o��M��ʇ̛����0�����S�p�tl������H�h�q����P���v�J#h��8O/��=O�O�Q�FH4]E
,di���0���
��4-1B�/	��{,�ŉ2U�6�U��J.�y�}�8U�ͣ�|f�}�0��Y�]o`ϋ/�&@����9A�|B	�BD��0t�b'���!|=%8|��Jk.�tf�}H�Fn�dp�"F�	2-!"�k�$!N��
���sU|ϊMW���2.�P���\f�6r(��K'��`QR�0`6�^鲤�<�aI��ǲ��~�î�����y0��{��/�$�Y@�ű�n{w�!0��:���������X�h4ӕq��=�_C
�|m�&?Paf��l�{v�g�%�k�,�`���f�\�bIC��~aBPZ�HP$B%:�rJY\ʣ5°��MoV{�	\�u!�0bFP��
a��0�伤 ��j�bA�>����oxC���֋��ʨ��84��-f��M����<���! ��w�!/7�8|�*���v�ᷦ�Z�M���Dn�00�n�Ys����
kB���S���Ƙ�M `�aC����PL�zJ5�l�fT��E�!���]v�y�| �#X�����cl/����e�g��zz�O��L2���j,@Ɠ@��uh&��Lʜ���L��5��B;Jj�`��s��kl��Ɏ��2�=�mi��U��
���H����BH� �W������!W�ok�l·�G>0`B�c�%љs�ɭḵ�W��c���=%���4GEO<3�F�B�s0�Q�"�#�L��ƨ*!�Q��E�i���v$����/���Y�'f�Y�U�
�P�B�s��m���h�Mj�e]541J� �F�+C[�5���eZ��T���NB芳J4��e�l����1��%^8����V�c�Ѡl��GL�pu+d�iy���6Q�FTDQf@#,1��3Ai��w�Lٌ/8�ga�C,�k��[,�X�#	��$`2, bF (@>�}��=�-w�X�]���k��J�>���UYs�ϼ6k�<Z�c-ц�*F���B���(�LbV�Ę'p��sg�����oƍ@�Ԁb$��C@E����q��vr�20�7/<�ƭ�V��D��e�i�ǚiyl�G�^wQ=�ysoL�h�E��fws��SY�P�Q엧���X86!1��<��=A��M�F�<7��=<�Ĉ��VJi�34w����p�EE+f����v��Vw����o���j�i���b��bl�š­�⮭�}Ba(���q'
���n�RJ�͝�Ŝh2U���;��0��Ss�J���uC�������]E[�.N�¸�K��e�FIBH�c��(����|{Wy8^����3j�q&�^i�M�Ղ�e�[x'(��梋�K^�>��he�B�n�f�l���!I6�E�|�(�V���V���,ϴ��ݛ)��ٝ7�����=~-R)3ʍ!��¥��?���4dbY!�!�
���#CKl"�"Q�&��2@"D�x�鶌i��2.��p����+���zA������X�_/uvqy����yV1��
�;��ϯ���P�"c!s;��m��m��m�� � ��  m     I�amk�[�	��]#+X	�j��
P�Um�m���m�A��жJ�]���l��U&p�`jT�X 6� ��/n�k�0 	kk��m[�H6�kl����LN��n���[\�hm[ ���Ym ��� @6Ͱ��m� ���  �` �κ@8[Vs���h  Jpi-��I�.�p	� QJK+�U9K����J	äԝ,�J�m��V�6��   [@	
P6�                   	    ��+�>     �                  $   l            ��                    h        �>    -�      ?�>  ����                   8p                     ~�       @     6�                |9�6�|>m�o�  m��qmm� �[L���(k�gf��R�l�cm�F� ��b��Pm׭۶�l[N $   ޣm�9%���T� p8����m�P��@$� I$ ��=��l����m��n�B@ �     $H�t4�mSF��0X�7ki�v:B�o[W�4�j��u���4�6�z^�ધ���@��)�Hݰ�ƾi���H�m�n�g%�. �V��v�a -���p m&�@�U)�UU���69Z$�u�B�[V�{^��m�sZ� $m�eU]J�8Yy�@m*�$FF�8qu��&������Mkkmۧ'F�ƾ�yz@&�I�vI�&�R�R�:��� N��=����6���m��X {)���R����+;�N`H$6�JH�۱'��Prx8��
�ۮ�G�m� Xa%�-�o[p8e+;l��j�` ӷi�V`y&�áuWZ���UT�݋(z��όb���S��-�=���-a�ʀ�N��<���T�.��5�-���bɴ�'[�m{gZt���z�׵��m� 	)���r�U�s9݊�ؐ��:m� m	����N	�y�6��-ŷ��72if�9�ĀH�l	5���E����a!Y$` I�
�� m��,�����p����h8�n��vj�{<�T��4�l�i�ӥ� 	-��ŵ��U�pl���r�ft9�_��u� m�n���� ���J����x�\��冓�D0$m�ڽh6�y/ YJ0�V�ڠ�y3��
���Чp+E&+5N�;;;<���`)m [[m&ݰ[R Km�mWinm� ��a�h�n�I4Ό7+N��ke@^��j��G[% �M$�im��d�h��  ���t���N[m�m�8r��]e�^Z��Wj��e[HH�� .���1�Ēr[Ug�mV1�PZ"f�
� ���8ۍk�'�Au��6TnGtzm�Ӭ���됇v����*�@�qӲҭU���r��3X��l��H����-<f� �Uq��*��������e]��)���y[��*8tmT��P  ��5-�
�����~WφI+���R��
�U@@]]�i_�|y@�UTګ`�u�;�$�8 @  vu��   T˶���f�[Am � N�R�ci7m�0�j�)t� $6��� ���q��	�l�v�M� k;0   �,�oa�@ -hMl��l����	V�U�UYUd��Km i���7m� �`�Ykm���j�ڥ���0o8`<6�Zl-�)Jl;i6$8	e�`	 ^�b^��h�8�L������CnMJ���*5h)��?S��Y~�[�Kn��8�cݞ�ZV
|�@n�ڣڶm[<�0;c�� �9ol3mnl�8�]o5�i3��Jk�8�R���J=�Uʥ��P��퍄���=u���)ۑ���|<��u��� �Ƶ� �/]���ǭi�i����)25WPt�tk�H��0�+*���@��J���*�N�S4�t����� T������5^ m�^�P�n:�G�v�I;u�vƼ[��UR���J��
 m�u$��٥^j��jU�Q�jU^` ���`j��ȷ6�m 7m:ˇ-��rG1��k�N��ցͷnr�IO�� 6N,�V�!&�d���hr�J'M�'5ؓ�l�Qt�+d�9�����g\lr����P6�������v*2�0�K��N�R�9�͝i\�lr���p.�m�f|9���j�L0��r�BB�n�j���UX:;E��h��R�[��۶:@ ���td��]X^ʶ��AcWLl	 u�-Y.�u��� P�J����Xv���$�Aj�  ���I [N�d��ڶ:���ZhC �)l�V� nM�]6M�t��� �   ��\��m&m�� �q*�j����vUylx]��&�	۫L�I���h�ր�Jආ�.��r�i.��6�oP �`4Y	6텶�,�tA�t�pr�PU[Us�3� ].�,����,m[�IͳvZ���n��kzޚ^�����.v}���7K7�g}J��y��YM�k���]���T�<�Y��UVQ��u�nX餵L��H��n��A��/X�S��q���~]�]�mqiF�燰����,�ul�޴[R[BH�:ҁ�F��@���=l�+l�KS{ m�c= ��m�H�]�6�}��w�I�����i���k�=�ܣ�W�WUe��`���Tһ9���T�ڤO����<` ���c m��&[�v�@.���  l $8�d�m�'�^Չ�촑�lӔ �ѵJ�e̓K#�Lg[#m86�5�zu�m��� �������e[V�]6 ֛kh� �l �`m� p7�|� �n׮���^���m   [@��K�1�V�j��K%H���k5�6�!�V�F؍k$��m'�6�Hk  m���m�,��� ���t�;I�� �M��m:�lk�������	�"�d�MXz��:�h�����v�Skz�p6�;A�v�  ��Bm{v
QT�e��� �P
�TH{E�/J۰8m�k�>xh�Q�i�rÆ�dݸ��#sh��d=�n���n[�-��5�n���+��ٙsFùN���^�b���4���s�Z��:M�]�9mU/�l�*�Z���z[us"6��49$sx� �Ewi��G�J�M�  �`k�2��q�NC6ñ��T	��st$ԫHL/cp�;�dtf �lDk@ lٺ�f]m�f��:Ľ.   ֘�$��I��m     m�Fl�:*�GQ啕j�W��)VWgm�[h
�gEʷAذh� i6�Mf��H� n����m�z��X�+Dk���)-�+[p ��]UGk���9xݶF` �m#��]�t�2��Xl�6ܵmvQ�s����2.�t���j|�;J۝�G$ݤ��s��]�t&��[*lG&t��"��4t�n�qmI#��(�$��hz�kpH٦�tKN�q8�HlN��Um@n�n݀89i��IĲ��5�	��קJ��u���8mRl.�Hpn����z�
�\�U��v��B`*�kk���iV����Z��a��cn':VĖP5���n�ѳ[��   ֶ�l[Eҫb��ж� �:���������٪��06�)@ v�՛`  [A���� �E�  ��+` 6�� �|  ��n���P�$�i#`h v�[ׄV�!��   )C�  � ��ѳf݈���%��  ��`�   �@-�  �h�+Im� l�{m�� [�ˀ  [NM����n�F��۰�@  6ۏ���|p ◤�`n�i\-c�5Ͱ $     p��6�d`Hڶ�UC�`�{-�UK��,$S����$���,��� ��ȴ�h�Jvij���o6�U�Z�qu�s�d��M[ Z'��lI�p�mu��ﾭ~�ק[�$�$�J�J�'.� !�%�-K�r�P W�s%���s�%�U/0��wv{UAĻ�5�����8��N���f��u���d(@��[S` �8$�����9:�:KoK(V-��!k=[m\͞�k��e���|���� �<���  ��٭`�%�g	gvŚ��1_`�SX�y&�f�m�'�p�B���ѕ��[��YV�6 ��9��B����m� 8���^�{���*��""�U�^*��GbE�� ��O�TN� S��6��ľ�0R��"!�)v0T8�Uد�j� ��&�J��"�LE]d� H@��	H��B$a$�d�1�	�h�T<Qv� �H�iU}H
F��IY��>��
0
�<O7�~P�r ��$�!	��HF ���a2@�		B�`�R!�B�p�����Â�
&�R����:Z�E� >
�V	��@"i>�� ;D]���I!1`@X�!"�b�0�ڀ���X*|�
 ��,Uh � ���c$CJ��T��O f �UB z �*�a�
����iG���P(Ib���]�z C�D�*)�%� �+�/�x���O�S�@�`'����ւ��_Q0��@J�� �A\Q�`���O�S�B(h��b��h | �ӈ(술��G��B$�$G�����A  ZI��^�j�U��6
�UN7L��Dۉ�8�d��ɮګ@�ͦy^�pv6���kc�p�{m�l   H��    l �(   ���m�m��   �l   6� �`H   ��Z��5��������X֌ie��H�0"`imUR-A�� =;M2n9X0�͐�fv�rc�5���*��	Q��v5���4Oeҋۮ�I�)u�ە�`�`wR����.�QnF�c�G2n\�.����z��iy�H�d�u�W=��",�ki���):z}&��Gyݺ���ͫ�/9�W$���qgb�z
y��v4��;s��c=�՝Ƀ��]80)�����ck�sGni���#�����
����}b3�� �H�޳;]�Н�sɺ�,�v��V�c�n�;��Y����I�	�n7[`�ٖ��d��&�.&�L�.��;l�h9��*&��a�9�g�br݂�����HӴ�[���<�e�a�k�v�^��e���-m�{<�v^׭�':�̆����qg��/��s�m�e�.i]�Z�cu���ݸ��U�K89wb&Y��cctG �Jl���-�끭Ѭ�[���5�6���a��Pl�\U�u�V�!��G��&*�{<r�S�F��.��vS`3�9{1��a�V_hܹ��:����:Y��vչ9pt� h��-��#F��aݠ٢���'����˸!�y8�Ս�ۭ.ܭ�Sm�����:��jӻA7nم����/F�C@)���_+N񶱆_�c#�C��y.6��Y�Vz�Zɕ'�%���\:7W.ۍ�[m[c���۞���6���'P���V�M��ɷU�ke��E��%^W����M[6�V�ۘ��'N��-����l�0+m�#�,�x���c�C�v���si�ǭ��طn��b�n���p��v�/V{kP]1�����^I��P�uh֠�.�n�k&f�\ֳ�q��"��ڡ���ȧʄ�hMl (? �U���'�Z�5��D��<X���ҭ,�Z���VVV^{:�2p�]q�ש�G�&�ݮ>x��p[��=�ad�a����w��n��;G��۴�q���6m҉�V8��S�:��0>ۮ��Gn�$��-�����Ń�[WOi�KϣP#�˓r�=�lv���j��S�롮��׃��ܻ���OU�+Ƶ�Ȇn4��7;&�n�I��[O��绮�{1�;�<�v3˹6L��^ɇ����9����r��'����m��m�NW�h����rz^��<�����IH�qh^�@��������Z�X�wF&��Lq���=ޔ�/;V�U����Y&9 R"5$�����yڴ
�W�U��jY0N��$�1��^v����{�z�)�z�Sz�o$S
Ƙ�p�k��yۮ#B�*�<n5��ã��v����١��&r�|�}>��t
��=ޔ�/;V���u2eչ�2e����>�{���qR���4+%4�ՠUz�ޱ�"��JT���sVg^v�&���������˯��--��G#RA'�h^�@��S�-�M�ݎȱ(�)����U��
��=ޔ�/;V�וǩ`F�	��byt�A�qnu�su�F0�{eX���W6��b#��152`ӏ@��W�[Қ�h^�@�Z��Lr`%##RB=ޔ�>�ՠUz����@�R	�v�$���@��V�U�B���Op����; �2jk��ꤙ�jji͆��ͫ'�k�z���Z���ɍ�c�DI���W����ڴ��i����{���6�D	��%Y���۝�bۇq���n�*�7S�`�%:�����rB= ����ڴ��h��z�R�q�qE#q�W�h{��9w�׬�>^�uł�bn�[����;��;=�f�B�73^����Z.X�wF&��Lc�h��ʰ�q�ew&ð�!""��zY�yuX�#$�#�M ��h���٠�l�=�:�?^�0&�t���cX�:s�	�ʯ��ql���ù���kZ�5�@�Ϫ��f�{�Y��� ��Ӳ$�6��0jE��� ��f�^�4y�Z�!�Ɍy1�I�I4�-�{��<�����@����%1ǋ#��{��<�����@=�٠�-�7RUT�v'�ʰ5$�'{�� �M�`���fq����i�@�$7q˷6��f�- m�ej�V���y�G�v�C�?�Ϟ��~r��UU�d�9.�s�cl�Iҧ^�}]hv9�:�ya�+��#s��bc �����6�5�nò�#|�wþ|�d�����;b1LkOd6y�"�������мGiR���ݫ�7��2ۂ�lJ=�N��<�/Om��g`���9��s<�Ow����������������bњݞ��ɞ���rl*u�;���=Q��^�Oq`���x)"r> ����x�h�@��W�r��qdbj&��݀s�c�B���nf���ڰ�f���cV&��&8�c�@/u���� ��h�[4�LJȡ"I�9&���@/���� ��hw&��N�,s���٠�l��f���@;�u�gB��=���Ti�U�O$pz��W��z�=����%�d�f]��o/��[4�Y�y{��/��@����r5N�4�n�3��}���JeH��, �m� E��vJ&����o*��c��9�1�}ܮ'#n(�m�&���@�Қ�Uf�u�4]q�
)�G�I��zS@=���f���^�˖#����9��4ު��f+���W_�@�Қ��؝Qc����B����_n�t�ۇ�)�j�n,tc��ۨ�J��N�R�m���߳@��@�Қ�Uf���bVIcs3#�M����^�B�3q�`��@;�� �ri���B�0�@�u�`�N;$�D(A�I�+u�]=������c��H��Vhz٠r�W�z�����5cj�"s	�w��/uz�Jh/R��b�Q�m�
cM�P��ۚ����Yi�.��k'(��s;�غ'�����RF���rh����)�}<�+b#�;����[NQ.Zt�T����)�|�J��l�9{��<�b9�Pi$��9��W��f���^��Қ�U�Xړ��L�(��w��/uz�Jh?f� @��I>U�`w���)�c�$O�$�/uz�Jh/R� �[4��;��6��&8�lQ��LIͻ�6�:��܆o����e&�6�C�G�z�����+���@��@���b�bh���R8h/R� �[4^��^��>�F�mdɎ"s	�w��/uz�Jh/R� ��V<�1L&9nMID)��mX�zXO0ʰ�IL�w^�U���I8�rG�{Ϫ�>^�z���/uz�u��22E�Cq���igmjG�ۉ6�9��Y&��Z��\�Ƹ]��"��F�d5�����n.v����m]<��{>z����W>�;��1���ծ_<�ᗨѓ���{IE�C�7;Z�I��c�������Ű�Nf��9S����j,�۴���s�b�J�y��Hk�f�vO�|�B�[dfNBaD��gk2�lP�'T@ږl�֦ٚ[��p`�.��{V�\��������v� �7=��h���c��N"n:j?v�O��t�[4^��y�Z�U�X�'���m�lu`s1��IL�=ͫ��ՠ|�J����\�$�?��h��������~?= �~�4�ɧd�m$9��zr���ٿ��$������$�;TԒ\����Iz��ejch���M8-I%��U��I~]?~S�U����$���Z�K�J�q7�6�i��*���/6�Ѻ�Ӷ�s�C4X�r��p]���R�u͞���?���~�/�����K��ũ$�����I#+ⲋ�NX쫺�W/$�z��V�/&!�&4�M��w_a2I&��>��$}V��$���\X!H��H��$���Z�K�J���=e&�����K��~�x�qq�7 ���}? G��Ԓ\����Iw;��$��U�X�'�q��|�G��Ԓ]��}�Iw;��$�ޕW��%mJf�#n �n�ź2D{-���ڃ/���p���nO\�-:��@mq4ڀ5�| ?������]��-I%��U��I��RI/w&��N���H��$���Z�K�J�n�#��y$��~�n�UO~n�:s�&<�����O����=e&��|�/�6�P�ZE��f�1��l��$���D������K�t:����� j[BYNF(RR�B�.��06�� I�L%�B�kH���+l+4f�]Q��WK����M� �"M�h�h,(B�J(B�(B�����iD�j�Fo5h�X�J���v4�h�4b�jɬe�b�
��.	�K�tB�3f���
�]!����H�BB���!X:3��flك�ґ�V�j��bE&:.�4�d&��	ef�0��$�,.��H��I!ăS��e�^�2l��	��a@(Fi�WSI(F&͊]`J�i˘�J��
jSLH��4Bj�����!NPA��f�m���0#p�L��(�,���� �a]�SD�ŗJP5����jC���A|T��AT\T`��&"��@⼂>*��T
"��h���������ֹ������{��]���ݮ��ɓD�5�$��)5$�zu_|�]��-I%��U��I_�"�S	�F��Ԓ]��}�Iw;��$�ޕW��$z�MI%ϰ�",\�-�q<<V����D�g��)��-�u����N�e�q�3�6ۆ���������$�����d����� 6�I����t�o��;��4�������]�$}���$�{��M�$���&~URz��?�5�3T�O������� ����$���Z�K�J�����b�I2D�'��)�$�Ӫ���wqjI.y�_��[q�<�E`@��d	�T
m���'����Iw��N	4�2(���%���ԒW�����$yڦ�����$~o��~Z%�S������v=��[lC&0m�:�<���ݍt�>�#8������d�$���>��$}_}/$�w��?���}�~�d�N��W꺐�ʷEʱ�j?�I#��5$����|�]��-I%��W��$e|V<�20��&⚒K��O�I.�w���ʫ��<�SRIs뎸�Ĝ��C�Kˮ�Ԓ_YU|�G�U5$����|�\�G;��[%dn~ �o��������q�����I���6I:��S�$�Ym�4�1!		�RABD�U;������lд�Q���ӵl4M:��[p�6َtN�e��u�)&݉�õ�=]�r�+�n$Ĝi���e咟l�.n��۱����8��GhW��<�a�G�3��{x�nu�B�ϵ�k%�[e,����_Vh�Bw\�Y7k���g�n ]����n�ݘ���w��d�M�[���n����#������t��P�:wGe��j���w��ߞ����r$jH��u��^�q�:��n�����.�N��rI��`��=st9�(Gg'�q�Ԋ?��K�����v��KϮ�RI}eU��IyT�b�I2D�'��G�$�ݴ����Ԓ_YU|��>�jI%��Ӳ	���ȣ��$��]ǩ$�����$�>�jI/wm>�$�A�1U14L�1ɏRI}eU��I}TԒ^��}�Iyu�z�K���8�\��n̓������| ?�w���ϺI=>��d�M���V�I�=�tFޫ��ܚ4�p1�j7m����Cص϶rm�[;��:s�:v�@�|/wm>�$���=I%��W��$y�SRIs���c�H}�Iyu�{�-��0�
Pm*�ă+H*X��0�RPah�m��p�#�d�]��[�H�_~��I;�Ϟ��UT�T���B�T�t�]�Y$��_���d��{�y$������'O}������q���i���? ��5��SRIu�������$��U_�$��H&+$�$BQ$�jI/wm>�$���=I%��W��$y�SRIw��o�KԦ=�� ۇ{]�j�ۮB=�-��o]� ��K	z7rR�Xl�p�o�I/.��RI}eU��I}TԒ^��}�Iz��b�bj!�#��$��Y�n�H*�?}��O}�~{�I��aY$K���DɎ	�$j?�I#�)5[o����9t�lTZ)�_/�l��Iz�U��IϊǑFF�$�&�?$�^����d����VI$߯��n�?(���^��fg+��r��9��cm�|�^]w���ʫ��=ғRI{�n�� ���y~/l�mvz�ʷ���rv���:���E�n��9��:z{r�Hi����k#$ǩ$�����$�t�Ԓ^��}�Iyu�z�J�����O�8ԑ'_|�G�RjI/wm>�$���=I%�������d�d�J##���K��O�I/.��RI}n���$�t�Ԓ^}ͧd�m,NdM��Kˮ�Ԓ���>��H���h�HAo���݉.�������rcԒ_[���I#�)5$����|�^]w��]��Γ��}<$3�d�V'7�6�%�{p�u�VN7#��La�a��3�u͛�"_|�G�RjI/wm>�$���=I%�����3��EFH�p��K�����EUOO�aY$��~��n�#�_������C��������A�Z�~~ ~����fg�˜�����5S�zX�zX�#�œD�&<rL�>�*��L,w���)������U;-SpGr4�@�t����M��s@�1�M��B��e�SaM��EM6�S\�P૥奝�UR�"@ �Ο�W�iU�]�MmgOm�u��ˬX��T�����5���)�swF����X�y���gF��3���d���&䮎pí�ۜUغ��@��N�k:�pskS��U!se��qs��=�{:60�R�b��n�ܗp��3���k�`.�9P�I+�.��f��/nWգO�������~4�Nv7�6R�m�;��g�N��wa5�d��@{Wa��mqT�$@�dr�?׮���U�w�S@��m;"N	�������s@�ت�;�)�{�S@���2rZ���1�[Vَrl�=�L�1�`ssmXg]e:�ԧL�h�(��Jh��>�w4�����T�"�S�N��4�]��b�@�t��y��Ē���ؠݞ��@x#��� �u�s�x�F&؝ �4��"@�I!$���빠_X��;�)�{�S@�i`�c��M:CmX�u�{p!
%%$��RF4J�!@�*�`J�)D����vnI��g�@����rʪ�㘄�A���;μ,w�6)�nm�{��l�H.+$�$@�dr��4�]���V���M˹�쉸�hc�#p�>�w4�Z{�4wJh�)@dM�8�`��$��L<1��a��.�I��Gc�E$l9m��)ƺǌ��3@��ՠw�S@�t���빠}z:�1L��872%Z{�/a%'s�76Ձ��Y6Wk�5L$c�FH�p�=�)�}z�i1fd4�RQ&sd��^g�bnd2%$��׮�}c�@�t����Mդs��c��Ɋ�4�u�`l(��^��ǥ��w-Xb���G0sێ�u����+ki�1z��'N񼻉��Æ-�dۜ�s7jk,�@�t����M��s@��ՠ|�AqY$�&,P29�Қ׮�}c�@�t�����vD�I41̑�h^��^��?��J����Y��>�Q
�)�2F��د��П{�vnI����rm`� �V�� ����#H$�+�w�w�`fk��B����UN�s`w�xX�����{����u��*��Q�(c"�B]��5�������v�˹�v�NQ��a���D��žO�]��e�oͷ�����;���\��_Hgq�`l��Z��
bs-�6�`}��W�2f�zX��hzSbG~i�Lq!1@�f�e���Қ^��>�w4ܲ��8�!9$�X�4?b�w�f����;��=�[�x�;>�)�m�ڕ,���ׅ��Q��o���k�`w�xX
�ϧ�p)�R��+*�!F
hP���4�˘�13�(����`�T�h&q��pbA� �א�x�O#��X����e23����N!�!�!-����X��(�p!A�T+���S�]��hR'���i��l�4sћi�h�*2h��4dX����᱓���&ך%Mbɞx�M��P���)vq��4˦RR2-y��V���Sii�fp�6�X���%D�I�i�'E	Ҵ�%X�E�#2f�f���J$�Ś��d�a2h�l�`Je`s�c��(t5��m�;��ƛ�0��49W�Ui�R�malc9�����˦f�.x��
%K�D�'(r�'+yQ`�������H�l�\�]v�U�Tsh����:q�Y�#kc���"�4����K�[�����%�6��`  �ڶ�  �`   [�   �    m�   ��    6�   ke���$[,�7��i��*�c�eA�(�ĭ�UA:�B\�ݺ�����wI؂z�nm۷*�=����]��F�q[�j�v\��ϫ6{1.��X[���0�-��V�zL����$QY��(�>��ݧlN,[���K��u�ga�7���k�?3�J�uf�.p��v�:��k��'#Ǹ�-�]h@톎�0��@p{U�E-��Ü\u���&(��5Z@d�s�rWn����k��0F�<��3<y�����u���p�Mvq�X|�����𫇷��Z����m{�bS��v��qԗ*��q�u'�'�.�[�
MwC[��ss\��랫�$�"z�-<���u��v��8��i��v�3\p�gsv����4�͝x/5�s��I�u�#���9�ce��v:l��=7j@�Ak\=z8%vҼb��D3u����zHnM!��9E����:��N��{$��wU�/[�WLű�Nv� �.L��P���g.�N����jklur�[��-�ܭ�F�<�U*��hy3���.9���mro »sUi�4�n�ͳ�h��]��nR.-��'uK���F���	������#�F��:wn,����=8,���j��#�/�?{4��v�^�s줦{��U�T�
LfW�'j�v0�v���I�`{�n�ep�䞲��:/J�h�Oض�M뇇��r�cW%�k��%.s��Q�]�l���&�m�t�KmUX�c
��0-�mm�n��[E�u��l�E���&���v�@N5��sln��檪ٲ���v�z}m�1slb����g�d�v�{U����s!lknۤ-j�v�n���$ ���{�]�w�^�� �P�`����P�Ңz�ӊ���w���ߧ-��K���L�:]q���H�m�m�WUT�9��<E!�{ZR�Ƴ��Þ"{G\e�[s�-�1�J8�2L��X��<��ֻs�NeðNuug�-���vNX�����l�'n{i��]k��������s��^v��W<��MؒIga8�[3��lg��ۓ��6]��gk<�[��n�۶�b��q���H)d�<r� ֠�VLר�j�7��M�S.���\�&:�9n-�Dm��6�n����GK��8��ѻ;Z&����jۚ�355*�n��{�Z�;�����R�C7�5l�$�����P�U2��.�/aL��zX���>�)�}z:�1L��I���C@�:�;�xY��y���3V=,�묚�Ӡ���e���7/K��K����Js�zX:�V��B��-�l�>μ,If��>;�K�JhYn+27��&�!#"q�K���������:��
�l�әzݿ��������`��tπ�X��d�$,�^��,K���o�iȖ%�by߷ٴ��$)!I
{��vZ�m�m�J��ND�,K�~�fӐ�;Uv�xE����HBHȮ����J����E�D���Ȗ'|�}�ND�,K���ͧ"X�%��O�ٴ�O�U��&�X����~/���3
f�f�&ӑ,K������r%�bX�w��m9�K������r%�bX���~x�h��4}_�����U\��J�ff�m9ı �<����r%�bX�t�}�ND�,K�~�fӑ,K���ͧ"X�%��Nٹ,��K���ֵ�iȖ%�b}���m9ı,O��}�ND�,K���ͧ"X�%��~��"X�%���ޙ��z�DLnqP�6J�b �h޻�n�a]C����j����{���ӫ�xv�:�iȖ%�b}����r%�bX�w��m9ı,O;�xl? "j*HRB�-�����$-�n�5T�	�L�n�m9ı,O���6��bX�'���6��bX�'�>�fӑ,K��߷ٴ�Kı;��5��S�cm�����$.no��r%�bX�t�}�ND��z�>E0Q������Ua`�Hj&�gy��iȖ%�b~���6��bX�'��g��K�I�L�&fm9ĳ����w��~�ND�,K�w�ӑ,K���o�iȖ%���B��VBA�䭝��[A4�m���6$�H���؛�H
{����v%�bX�w��iȖ%�b}���m9���$.�L��`��)bd�c&jY��˘x��76�<�a���b��PP\Sm�ԧHN�.�)!I
HY�z\/��,K���m9ı,O�}�ͨ�bX�'�}�ͧ"X�%�����u�˭e�WWS��M�"X�%����6���%�b}���m9ı,O~�}�ND�,K���ͧ"�bX�|d�N�5JU�7p�!I
HRB���ӑ,K���ٴ�K¡D�Ow�ӑ,K����siȖ%�$.n]ku*ZjSmU8r�M���$)<��MD�����Kı=����ND�,Kϻ�m9İ84������>|
!� `&��ڛ��
HRB��[5T�h�M��ɴ�Kı<����r%�bX~`����i�Kı;������Kı=���m9ı,N��}�-�SS'������q5ɢv]̧�g>��m6��@eN.�gIt���L� ��w��Y�ŉ����"X�%��~�uv��bX�'�}�͊r%�bX�w��m9ı,N�%��)p�0̷2۬6��bX�'��}��r ؖ%���o�iȖ%�by߷ٴ�Kı<������7��������rWl5U����%�bX����6��bX�'��xm9ı,O>�xm9ı,O���Wi�
HRB��d6Mn�s-	�H�.D�,� u�߿xm9ı,O{���"X�%��{���9ıJ$�����|B�����ܪ���rj��a���iȖ%�by�{�iȖ%�b��{���9ı,O~�}�ND�,K���6��bX�'����/����Hʘ�uj�.�� U�s�ۉ6�9��R�!&�3SKo���K�+�I.P�(��8zz;]v8�ڑV�U|Pj�y�f���\�݊(����[q��9�8UT|��b�X��r���e�,��Z�hƀ�E�u��@��֔�ۃ�k�tn+�Y\b�9��3u�ht\p��˹�[s���0|��x���8e8ol-5�OZxZ�/R��ݤJn��Ѻ�z����.�nぎ�v�y�r�m�V.��R�~���q���?o��ӑ,K���ٴ�Kı<�{�a�) CȚ�bX����ND�,K��޿fj�)����\�]�"X�%���o�i�
�%�by���ӑ,K�����ӑ,K���ڛ��
HRB�1e��UjZ)7����ND�,K���6��bX�'�w�6��c�P��!\��?o�WiȖ%�bw���M�"X�%��zt�Me�k#32�e�6��bY�*�'����iȖ%�bw�����r%�bX����6��bX������߼6��bX�'��/I�I�����iȖ%�b}�ﺻND�,K߾�fӑ,K����"X�%�����$)!I
H\ܝ_K`¡����[2�Y*��=��[;�g N��rI��X1�O\����������~���e��4�=߻�oq��N�����Kı<�{�iȖ%�by�{�a� ��5ı;���j�9HRB��$='��NF��L�˅��bX�w���>U��A^�cbj%����ND�,K��w�iȖ%�b{����r'�*�Pr&D��������T.��1�m�������D�����"X�%��{���9��Q���j'���M�"X�%������ND�,KϏ��f�s%�
��a��Kı;�w�]�"X�%���o�iȖ%�bw��fӑ,K�A�Ww��_��$)!nmכ�R�R�j����ND�,K��fӑ,K����߹�m<�bX�'��~��Kı;�w�]�"X�%�~����V��O�c����d�δ�vm��m�l�;���:��ܽ���]�`s�b��N[|�~oq��%���}�ND�,K���6��bX�'}�����CȚ�bX��w�m_��$)!z�O'Ls%1n[e�"X�%��{�NC�G�h��L�bw�ڻND�,K�����ND�,K���6��bX�'��~�L2L52�[s�"X�%��{���9ı,O��}�ND�؈J�ApU7Q3����ND�,K����i�����oq��w��rWl����r%�g�  %r'�߼��ND�,K����iȖ%�by���ӑ,K�TY�����ڻND�,K�����t�jS`Kl�_��$)!n��6��bX���_~���%�bX����ڻND�,K��fӑ,��ow�ݾ�+���)�7l�����m\���:���8Ɔ�	��K*���)y}
"��������QNJ��\.��$)!w���iȖ%�bw�ﺻND�,K��fӑ,K��{�ND�,KΟ��^�K����iȖ%�bw�ﺻNC�@ �&�X�}��v��bX�'�߿p�r%�bX�{���r'�"���bw��_�5K���Z�.f�ӑ,K������9ı,N����Kı=����Kı;����/�RB����.�j�)��I��̻ND�,T,N����Kı=����Kı;�w�]�"X�ȩ���%�`aB1`�!�ES�����'{��w����$/Vx�ꆊu*Fܶ:kiȖ%�b{�{�iȖ%�bw�ﺻND�,K�s��ND�,K��x��)!I
HYY:���T����k/7J�\T��m��l�og�qq�lR�=��g�rŉz���ߓ�g��u�����WiȖ%�b{�w�iȖ%�bw����%�bX�����r%�b]�?��NJ햦��|�~oq���b{�w�i�~#���b~���6��bX�'�~��iȖ%�bw����9�BJ(�D)!O�O��t�jP�T޲�9ı,O߻��ӑ,K�����ӑ,�MD�����iȖ%�b��7����$.��UV�.�%MM;5u�m9İ@�=����Kı;�w{v��bX�'��{v��bX�bw�w�ӑ,K����vY���p¹�5�m9ı,N���ݧ"X�%���ݧ"X�%����ND�,K�{�ND�,K&1!1XĎ��Aa�a�F�T� aBEJ��>}��?������Cû5 mRN� �[q�l�j�u�ֹK��[\p��,����N�D!���n����bs�;C��m�zm�,!��{�v.�N�v��'8φ�^ѧ��渒B&�"�ɚ�8�*�Ա�ݩ�ҥ�ȒL���$y9��pm�]��F4q�6@��qζx�5"爭h��矁����D/�N��	�{[#jy�i �:N#i�@��͒��&�9�9[Q��7(�����0�M�~��w}�5��^s̫��Ȗ%�b}�~�v��bX�'{�xm9ı,O}�xm9ı,N���ݧ"X�%����;rɬ���-̻ND�,K���6���"0GQ5���߸m9ı,O�~��v��bX�'��{v���@D�K��{?֦Y�\̺ɚ�iȖ%�b}���6��bX�'}��nӑ,K����nӑ,K��~��"X�%��g��nY�.\�2۬6��bY�*�D������9ı,N�?��ӑ,K��~��"X�� 1WQ>�������oq����������j���9ı,O}���9ı,N����r%�bX�����r%�bX������h��4{����\����7*�`m�e.�(�ٓ�G6�Tu��v��=��p��������)�p�����ap�a���]��,K�����m9ı,O}�xm9ı,N���ݧ"X�%���ݧ"X�����}U��tdF25�=ߛ�o%����!�1$Ⰺ�!B�d;�h ���H1�@��+,eH	j���Qi�B�'�qU�W��9"X�����iȖ%�b}����9ı,N����r����&�j%���M�f���p¹�5�m9ı,O�~��v��bX�'��{v��c�
��MD����m9ı,O����ӑ,K���w�����)��k�\�ND�,�"�"+��}�߮ӑ,K������Kı=����K�� ��߿r��ND�,Kޝ���Y��&�%̻ND�,K���ND�,K �@�}����Ȗ%�bw�ۿ�ӑ,K����nӑ,K����nkW5m���{[�ڜpHO���+�s��^A�Eؔ�&�5UCALCni7M\/�RB������ӑ,K������9ı,O}���_�_"j%�bw�p�r%�bX�����e�fL��&e�Xm9ı,O���nӑ_� D�K����Kı;���m9ı,������)!I
HS��uR�m��u�.ӑ,K����nӑ,K���w�ӑ,`�$���$#c� ��������:���N��QY`ǘ<� '�,2U�ԥf�p(�ExK* r�%��Rq��<�ּ��<4n�tl�Iu�ʰh��/&^^*�꫅a==}t��h�]>�B��}<!]6�m7䤤�b	���($Ji�c	�Ytˡ�@�B��ᘳlٻ��8�� ��ű��	�T�5'
(bL~��ǈ�߽
CP��{ǀb�(����0���>t�Ip&h!� �#���֎'��9�Le�)f&�ӿTSV���tDK5��c�f�5���K.�U�]��d֣�3H�RTb@�a��!�
|���&�}@��ꠞ��
!�A�@p�D"
������P�4 �U*�'�3���iȖ%�bw�n��9ı,K�{5l�f�a0�f3Yv��bY�P j'w��ӑ,K���߸m9ı,O���nӑ,K�s��ND�,K������hȌl��{�7���{���{�ND�,K�{�۴�Kı=�>��r%�bX�w��m9ı,�~�}��gB��[]�R�ӳEӎ���ݍg����t���[�V��p#���Oφ�8���3Fk0�r%�bX�{��ݧ"X�%���nӑ,K���o�a��>D�K���߸m9ı,O߿]��sT�e5�k̹v��bX�'��ݻND�,K���ͧ"X�%����"X�%������r(ؖ%��a�\n��X쫱ʹ�ֈ�#G��}�ND�,K�{�ND�,K�{�۴�Kı=�>��r%�bX��0�UC@����e���$)!BV'���6��bX�'��w�iȖ%�b{�}۴�K��q�A��`�"nD�{�M�"X�*HY]�59�ۖU73-���
HR%������r%�bX ��}۴�Kı>����r%�bX�{���r%�bX��ܟ��S%4B�P�+6q[���l`�u�퇓�s������cM�vߞ��5�%Z�+G�w�����ow߷]�"X�%��~�fӑ,K�����ӑ,K������9ı,K��S&�R��mKm����$)!I;��6��6%�by�{�iȖ%�b}�w{v��bX�'��ݻND�,K=߯��_�#FDcem�������D����ӑ,K������9�K�����iȖ%�b}߷ٴ�K�F����?]9r�ˢ���kDh�,O���nӑ,K�����iȖ%�b}߷ٴ�K�[�{�ND�,K���n\�.Mf�3.]�"X�%���nӑ,K���o�iȖ%�by�{�iȖ%�b}�w{v��bX�'�U$GI
yM	�����;�w�AYV���`k�ZY�AUU*�[*�uU^y�R�����'%�M�=�T�E2��v��ؘ.�a��n-���]h���[¡v�8rra�8��<��6�H'�n
2���Ͱ������P�����6F)c�3��k�c��N�"e�vU�agY���������*�F�W'v25vM;n��=���I�%a�3������67]�"W\��������w����J�&4����v�99��ٸǓsv��/*��d®Ѯ������|)
u4��t��7�)!I
HYݿ�,K�����ӑ,K������?��MD�,O����ND�,K��zyUS���4�l�_��$)!s��NEı,O���nӑ,K�����iȖ%�b}߷ٴ�O� QTB�W��' �&�d�s2ڸ_�K��߷]�"X�%���nӑ,K���o�iȖ%�by�{�iȔ�$)!OL�55Cm�dӗ7��g�1Qu���iȖ%�bw�w�m9ı,O=�xm9ı,O���nӑ,KĽ��V��j�,&as3.ӑ,K���o�iȖ%�a���D���߿xm<�bX�'~����9ı,O}ϻv��bX�'{�ާ{1�ci�ѵ=�\[a׮���9�`u��c��p�ݘa��bnjeY�ё�Zm9ı,O;�xm9ı,O���nӑ,K�����h�~ b��MD�,N���ӑ,K����˫f�ɖjC4\�6��bX�'��w�i�P6;����0X$Q:��@��@xȚ�bk����Kı<���m9ı,O;�xm9�"PT`ș����w�\��-9T�bl�p�!I
HRB��~�ND�,K�{�ͧ"X�
$5Q=���6��bX�'�~����Kı\��[.�K*�4�)�sp�!I
A%�T��"*�O�����A>����bH$��O�7�?�}�}۴�JB�����UU9�sJ�5p�!LK��w�ӑ,K�� ���ߧ�6�D�,K�g]�"X�%��~��"X�%�O~/�2�!MB�B�7CSK�F����g��ݎ]wև���ɯ��s��z݇3�6��u��W~{���7���x�ߧ�m9ı,O�ϻv��bX�'���6���bX�'���6��bX����o�Ћ��+o����7��,O�ϻv��bX�'���6��bX�'���6��bX�'��w�N@�,K�ߦ��̷0�Y3��v��bX�'���6��bX�'���6��c�
5Q>����ND�,K1�����$)!I��UU�6J��j��a��K���������r%�bX������Kı>�>��r%�bX�{���r%�bX�{�캷��s5n�3E��iȖ%�b{�w{v��bX� ��ݻND�,K�{�ND�,K���ND�,K��m�ʽJ`@�FJI�"���ܼ�k��:��&����ʚ<$1qts][�#��%�bX�{�v�9ı,O��xm9ı,O;�xm�Kı=�����h��4w���.��ꭻ.蒮m9ı,O��xm9ı,O;�xm9ı,O}��nӑ,K�����i�*%�byܟjt�̒f33.�f��r%�bX�w���r%�bX����ݧ"X�%����nӑ,K������)!I
H]��6��L�i�O5.a��K��=����ND�,K�s�ݧ"X�%�����"X� B$T�QX �s"ss~W����$)�5�5Cn��n]e˴�Kı>�>��r%�bX�?{���r%�bX�w���r%�bX����ݧ"X�%��~��&I�ֲ�ź�����˻7�r��o���x����9�Z�a�,�P�{�'��u�b}�{�iȖ%�by߻�iȖ%�b{�w{v����Q,K�g]�����$,�mUW�l�54ԩ�է"X�%��~��"X�%�����r%�bX�{���r%�bX�{���r'��?�*dL�bw��eտ٩s5n�3E��iȖ%�bw�ۿ�iȖ%�b}�w�iȖ%�b}�{�iȖ%�b{߻�iȖ%�bw�﹙�B�S3P�˗iȖ%��X�{���r%�bX�{���r%�bX�����r%�bX����ݧ"X�%��Z�\ҖU0i�sp�!I
HRB��xm9ı,�$�a�w���Ȗ%�b}����iȖ%�b}�w�iȖ%�b`	����]arL��j���jU������m�sm������Řvp���;c+�s;kv�!��vż�2^-k�8�m�y�U�vz�[WZ�XNv����ƚ�wnP�f�ڑ:v]ܛ'dڗ3�CY� �z6������lS��Vz�mY���[d��v���p��޴��뭹����dAa��ѷn9��n��d�4�m�*�:��V�^�Ϭ}�S�e��'�i��..�Oi����w�e�ƣ��k)��*:�u�`B�tK`S��4��]��)!I
HY���iȖ%�b{�w{v��bX�'��{v?�D"�B+! Ț�bX����ND�,K�w���rA�M6U7D���)!I
H]�����bX�'��{v��bX�'���6��bX�'���6����" ��&�X���~��WZ����s%�\�ND�,K�g��iȖ%�b}�{�iȖ%�b{߻�iȖ%�b{�w{v��bX�%�M[{��4e�����]�"X��3� B`��H�?w���iȖ%�bw����"X�%�����r%�`�Bܿzn�)!I
HY^ڪ�P�95uu�.��"X�%��~��"X�%��$D��ܿ��Ȗ%�bw����9ı,O��xm9ı,O=�
�D�JbK���2rm���k�ۃ�	t��/hJ��MŻ�Q�)�8M��fND�,K�{�۴�Kı>�;۴�Kı>����Ed �&�X�'߻��ӑ,K��������.u0�5̹v��bX�'��{v����C�@!���� ����PpQ6���D�Ks�6��bX�'���6��bX�'��w�iȖ%�by���˗VeֲL�K��iȖ%�b}�{�iȖ%�b{߻�iȖ?Ȅ��2'{���v��bX�'�����r%�bX�u�F�-�N�ҧM\/�RB����w�ӑ,K������9ı,O����9ı?]D�߿xm9ıRB�o�g���eStKj�|B��b{�w{v��bX�'��{v��bX�'���6��bX�'���6��b]�7�����ߚ�J���;��zy��iI2�j� ��Q.\L�Rr6M)iͯ!D+���ʚ��M̶M9sp�B�������9ı,O��xm9ı,O{�xm9ı,O}��nӑ,KĽ��ou�f���0��˴�Kı>����T�,K���ND�,K�{�۴�Kı>�;۴�Kı=�r��hl�54ԩ�����$)!I��xm9ı,O}��nӑ,w�3�%P%
-(5����U"��UJ E� P�V��OM����!��D�����9ı,O�w��"X�%��n˫{��3R��4\�6��bX�'��w�iȖ%�b}�w�iȖ%�b}�{�iȖ%�b{߻�iȖ%�bw�﹬֡�2�a�5L̹v��bX�'��{v��bX�'����������,K���߸m9ı,O}��nӑ,KĿ~���d:��Wv4�pD6�nR���M�<)������r��WXݮ��/X�жՎ��v��bX�'���6��bX�'���6��bX�'���u��P�Ț�bX�}��]�"X�%���;��R�Bk�ˣY�6��bX�'���6��bX�'���u��Kı=�;۴�Kı;����_�dD5R��[����4�T�L���)!LK��{�[ND�,K�s��ND�,K���ND�,K�{�ND��7������ �UAC��~oq�Y���?� ��;�]�"X�%�����6��bX�'���6��bXqET�QL+�'���u��Kı/}�շ��3F[I�\�e�r%�bX�����r%�bX  ���(H������ؖ%�b}�������bX�'��ݻND�,K=߿�}�W��Sn���/mp��. ��fc����Wn�ךWa��+bE[��)u�m9ı,O=�xm9ı,O;���iȖ%�b{�}۴�Kı;����Kı<���uosV�Yua�3Y�ӑ,K��~�� ��  ���'�g]�"X�%������Kı<����KĒ�޺uB��Rj��m�:�_��"X���v�9ı,N��xm9�_�PD�O~���ӑ,K���^���)!I
HY�-h�j�5I��R�.ӑ,K?�B�~���6��bX�'�~��iȖ%�byܿw[ND�,U�����}���ND�,K߲wS��̄�35�F�Xm9ı,O;�xm9ı,?����{�[O"X�%�߳��ӑ,K��w�ӑ,K��|L�"r�Q��P�o���5&i	zJ�sAR9�SD��(Jt$0d	���`NN: �ѪK4:D)Jg��*�*@����R6S<5B۴������	CXL�B&,�d�%����b� ���&:@�
�y��
H�(R�3Y�3{`Di�i��B�p"!Jq���)�yM��U6 $h��kl�	f��p[�f�v��6��^U@H���M���,�I�ti&�����   8��p  6�   �    8    p   l     �`$   �֊Z	{(��(rŚ�	�i#J�dh��"�� ����ʝ�����kV8�ݮj�hl� =��6��N�E��L�������!H��d�M��*ڮ��͹7ah�l�-����פ+m9��&k���ny%z����\q�ö�Pk����l�ezc<9F:D��n�t屡);l�l�2 �A5�㢽.Q̔��`C[n�J��l0�{VwWX���νG"�ׯ�SF�I�p�N��y�ln�Šx��ņBc�Vj��Sی	��lv�m��E�Us���m�ۮˈg�P3ք�CӞh�pv��i����M�<W%θۆ-q�L\n��00��i�^�8U��>�ds6p[v�P�zz9��Θ�ښ�%%���[r����N��iݡ�\kf�Yd2t���ݞ��ňx�,;�v����b-�r�m��i�rI�PhKW6uL��Bn$�m;�'���󦬡u�1�p��/�6�r�����E��㤎-�k$Wm]�cus����8xr���\����U�`��ݔ��f�1����m�	\a퐶v�qyG7l���Q;�Kv���� Q�Ẩ���2,s��̻��]�&q�n�{i�q�ñ6�vB�8�b�f���э�z�uj�ݮ�P�6�j�؎�Td�6��`�WvS�ۣOY���f�zT\��7/ml��9k��}nf�лnr8;\v�N�s��k��#�]�vF�U�Gh�4�{\��6�7m� �x�T�d���YN)ۆ�`�6⨷Ӳ�KLR�	����� %��MwT
�5R�Ñݹ��Ң�u��W�OgVx`�VC���ee4�P�h��ݺu�7�N�3�u���
ڂᘋ ����D�����@������\|UO<6�Pt oy�̓Y��fh�.�o;��R�N�t�uM��M��l!��X�IM�0�g�B��,�t���n��[p�::+\��=��W�ٞ�����p��v΋d�Wf�mqp����{G�m�{�w5e�n��ӝ�r�֙�tꮦl��$�+ŻN��sk���v�ݞ���{s��Cs���y���c�^75'����I��ʼ7�M���%�+ax�r���뇁�H]*\�eN�t�g����ܜ&�K�����.ĊS)���fj\é�Kı=�/{��"X�%����nӑ,K��w��C�,K��w�ӑ,KĿO��dXJ�(b�����7���{�����"X�%��~��"X�%��~��"X�%��r��m9�CQ(�$)�iS3�`�9�Cj[nn�) �,O�w��"X�%��~��"X�%��r���r%�bX�{�v�9�q���}��f���p�|�~oq���GQ=���ND�,K��{�[ND�,K�s�ݧ"X�%��~�F�F��;�dr��u%�r�.�w�ӑ,K��~�bX�'��ݻND�,K���ND�,K���ND�,K��~�ML�.Y3L��V�6	��=z�n@���G-^�73�m�����_�3i�͹���{�'��u�,O�ϻv��bX�'~��6��bX�'���6��bX�'����iȖ%���ޙkGST9�`�*]9�_��"X�����r}0$!���"��Td@�P��D�(Z� ��"2�B�� �#	�+!*�D��!t��F*��&�j%���6��bX�'�e�u��Kı>�>��r%�bX����N�\�Mc3Ytk5�ӑ,K��w�ӑ,K��{�m9�ı<�>��r%�bX�����r%�bX��ս�d�2���[W����$.k�ڸ_�K�����iȖ%�bw�w�ӑ,K����iȖ%�b_��w��kN�[m̷4�\/�RB����6n�X�%�'{�xm9ı,O>��6��RB��v�f�Ϊ٭�4�Rn�J��t�K����\��A�2d�9��^;���������"K"��h��hw]V�]��P��C�Y�`v{�ۧM��5SM
[j����W�2su�ٰ̬́=m��>��M+R!4dx���[s_]�9���x���$�F#� ���JJ\�$e!�� ��� ��wf�w����KldȞG܎8�?�ٟ��_����ڰ>�rՇ�N��l��h�6D�	���=m��>�:���Z�������Q�m�J����n���	�^^y���ܦ�Fg�c�r��!���dhrg�z�ۚ�:��]��DG��ݛ��T�9��ˑL�-�ՠ}Ϫ�=]�@���o�$��
�0��:��U-��[��Nl������Z��s@��V���
�4��3)�N[sa�""{�vlfm�3d�uBR�Dw��9<�mӦ�(�Na���z���c�@��R����XJ�MѨ��TS�X4J���%��oc��a�x{m4Y�[�l7jȏ���$��I��tKtMH�)m��W��`{�)�Uz��[��^��0�$�*�n�X�^�(J?	Cg����`_���nhW]z�t�F�"n���*�^�����>���{�4��(t��j�"[��
=B�U������^��������X9�NS�ɑ�9#ds4�����M��krNy��7$��z@	1"�@`��""�E��Ǿ�6���J�F��M�Ò9�ll�E���  �Ή^;[t��m�5J]�7)�lmn䬉�ʏWOW:v{L�+pq��K�a�m��՗������q�F;�j��[=<�l:�Sp�Sķ<s��:��rkkz� f�k�nW��<�IiѹkՠF�5۷��ub�M+��I)�@����]��nC�]A�'�ȽBtm�T�bcd����t�l\D$��J�� ,F0X�  � b�D�F1E H��I�b� `!��s�5���B�P�Ǧ���
��6/]k`x��{���!�v��zݳ�Fۍ���8�|��������k�(������Ձ�����0m��.5�7$�������*$`�P$D"�QTw=�V}S�U��u�`r��GɑDڐ0R=�[��}Z�����ΐ
���>�K��	�]h�:"~"�A" D"�!
��;�`{5��2{ܫ�<�����׮�QCC���Tۖ���:�=�G�@�����p�j��*s*��:���ʢ���U#k�vk���8�r]�.�m�F*{m%���k�팽i`v�`��
���>����v���M�g3(t��j�"[��fZ����J��Tz���u>���ܓ߻�������F��2djH���̫���͈I/(""�ӻ�;��� ���q�"s��G�{�)�U�^�����>�uz+����L�rԺl�2yܫR��ww��ڜڰ9μ,Зw&��S�j��:Br��]RK��H�&�z[�;����+۳<<�3��V�8�L�&ԁ���������W�{�)�>A�u��~��O�JF&��KmXeOr�b!%�J*��~,No������/Yc���G�D7$N=�����{�1���iL�4�R�J�
���}��ʝڰ9í`�j�5L$�l��(Q���X����U��Q=�^�;FQ�:r��5N��Ձ�3-XI(�ͯ��r~4K�\�b�bL�$,�����t�ub7Ò�t��ֺ.wpj�����݇6j8�&G) ���~u�zwJh��h[)�p[N4�NcPn�Ձ������D(UG�޵`w�~,����A��	"K"����3����jP����k�3����s&Ej@�$��e4��5�'���M��0�Bjp��u}�6��9RW�%�9Q�I�e��WqՁ������77mX[)��*�o$m	4
!����o-�f7]�qv�\&�<W6�<�l���:i�:�H	�$�@��M�w4���g�(�C�[�������aL�e���̵{��%G}�����u`w�t�;�̬��&Lq�&h[)�}]���)�[n�U�U�2S�-�]6XlB��(���u`n��`[n��������JD�5
m��;޼,�%���D!	B��������?�}]���ȓU4HI�K��L�u�m���@ 9V��j����vH�����D$ݡ��m[k��ʆx�W��|]D#k=��E�ys�1bα��<,;\:`y����j��eV�v���燫�N��>�K3tN-�[�۱t��ɂςI%�l���v�N۝��i�J%�^�6�����x)��� �r��&����i�iAݥՒw���~|�;涕���X4B�Ŝ��ݫ�����e��Mf�λ/S�\�A���p&H�Ȧ(�>�n��������Қ���s&Ej@�#Vُ��%��BID6g���Ձ����4m��>�!4�iH�ё����V{ׅ��S;���n�,�ǎ�QCC��M6�ua�_��BP���������V9���Vq�)l#p$�@����gwoO������ɰ>�I�d��*���o���tF����ynwnܽv�<�[B�k��k^e�yBJ?
;e����S�m������+1Ձ�Vd����7wmX�ҧi�&�:R�%�e��Vc��I%*"�P��+2l���ǅ�(_����$�Pi��:*�̷4�Km����-�w4z�hWlz�ߦ�WY&��i������@ E!B�~��`n����V9Y�`}>�H�2(�S'�f��YM��@���@��������BMob���v6׮�ZNL%�s���3��ڭ/Wu������I����R'I�g ����@���@���޲��,j4ɑ<RrI#�=�j�-�s@�����Vc�Ԓ��3kA�U�aL�s`n�ڰ9�xYȌjx��L��K��A�g��[h~�K��H�v�f���!I7�Y*K!Rf�4g����G��!e暤�x:*I|����.�ѕ�7Z�z� Ka ��0`���D�2��Ц�S3dB�vc)9�hH_8&�
oa��DY؄���&c�H�<�p8k�9��������<��$���K5�K����莔h&6��	BT$�(�*F)D"�H�������! �&�! 4���#<eF P7�P��%���H��l[B�ʿ�@
+ ]"�b- Sj��U�Et*�@t �� t	�b���! .��g����v������a���f��YK��V9Y�a�!DN������:��y��C@��c�=�j�.fZ�9�xX��:�:���CSEJ��G5�k2R	�^������gv���7O�B�v@�cq%�8��I#����h۹`s���D%�!BH"9A�W����W�E:�h�rJ�i˧6fe��(Jd�wmX��u`s��6����:i�.j���V9�j��+1՞���
IUfW�6��Z�9�rML�[U4�t�mXef:�9�̛32ՄDBJ*)
^	�}xco�����R�;��r�m��9�̛b�	����^����3=�V�YYV�L�)�D�^�T�6m�4����;����̝���:�0Jx��F��8<N	E�[�s@����>���yڴ�9���$a����rO<�>�蟖) 	�$�
����3+ޛ3�j��s��2dq�r9��@���O�!DL��ڰ;�zXN�c����n��h���nN���S� V(	J�߿M����Z�9�xXeeeXy��q��,jdQŠ[�s@���
;ݽ>�[[V9Y�`8�$��
q����_����l�3j˺�������86��I���V(v�.�ƙ+<we�Lq����G�ݮ0:�v���קX5O�% V��>l�ܱ�y��lmn�L'���<.�,+N�nC����=6![=Y�]�du��y����Y[����Ay4��'=:��ey�%oCvw<V��\��m;q�[��`��p�.�g�gՁ�xۤH�����������6�U���Sn����6��s��M�sXs۴f��j��$��u�_���@E�EH�^g7���k2�֮�]3�Ł�VVU��Vd��Cw6Ձ��!4�F)�"<��@������ń��j��1��P�B��BP�
�
����Ժ�`�[	�ۧVc���o]�޲���^��t�o��8$I�o]�޲��וa���$�� D%Y��M��F��dqa ��f��YM��@���@���W+�Ս�"JcFF<��V�س�C��ɶ�����:�޸�{.�{9Q�28�9�����h�h�e�Т�$��!������<x?~tM2e7NJ�Knlr�����"Q
���V;�K�c�6�|�#n19�L�8��w4�e,�D(�ȈM�������`}9�ۧS&Ejd�RL�>���>��-�}V��n��X�ұ�Ɠ�G�}�x���	y(Q�Kw�~���~�j���S@=R��25� �do�3V	��۫6�
��/K���Sg��M�k�^]4��&69���E�{Ϫ�;���>����(J>��u�pǠꪐ锦�26���s-_�$�
��y��;������U�z��YX8Lq�&hy�}7$�g�w(j�Б*B�����!j�����w$�}�f�NaS�̉�N�����В��w~e����w[��}�)�p[��Cx'!�{Ϫ�;���>���>�e���DBK�O&�\�uI̲f���=+{mV�Su�r��96ygs������͡L�kw��Хۛ��S�i�UKN]9�����YM�[��=��h+l��2dQ6�O�$��YM�[��=��h�韐
G���J���ʺ���K���{�톁�>�@�s@�zנ^�ƣm�UE4Kc��BI(��^l������DZKz�G �U
a	L
�])R��e%Md*Ń�֐�+��*(@CF�S��W�=�|ɹ';=�ɕUHt�*�3#nl�2Ձ�P�ݽ>����@��U�w��,J6�M�
7*Ыpv�1s��/2<u�[�gr��x0�F'�VHGjI�޲�޷a�s�ܟ(��f����̊�NS���s`}��e�B����ٰ33mXyڷ��䃌����4аM�y�Z{֙�Q?r�&����,�]���S�i���Ö�$�V�����ޛ��a�wt����s$�5?��4��h����4ϲe���Y	ry��j�Y5s5��t���z4�� mRN� �[p�6���NGY� ���h�Ş5�&�S�d伺�똎"8a^&c�2�{f��v�؇�wx��9۠ҏh!:��@9�
��e6�:�@E�3\���6����R�Sōq�+���8l���jDI�$x�
y͜cJ���^n@������e��ht3�����u��r�4/ʹ��оcK��#���n����6+m��r����TU�������&�щƓ�)�P-��wJh�w4
�W�wYcQ�c��cN�)�{���*�^���B6���q&Ԇ��s@��v~�P�D~o}��,߼�2�є6�M0CT�m��;[�Vs^�g^�������j�nG�s��?(��o�8o�j����XI����`�qø�MTkk��M�������\m�ކ��n�N����l����oJhW��>�)�}���;�W��KW.�6����D�	|�$��K�
����X�~,�^���F4�d�93@�z�^��=�w4^�&ӭ'�RK
n�?~���{�?�y�,w�j��z��e�F�"70sp�:����u��9^�@��S@��XR���9*g6�'nk����h�.�q�1�b���"d�a�;c-������J,s2Ձ��ʰ9�x~��B�u��~�g���ls4�6KmX�̫�ǅ���ʰ9��W�%2rw����R�鲪�Ձ������eY�G5.��+��5���h�JJ -T(��I((QRP�aR @KJ#, �B�U�.N��ڰ=;� �L�rZ�dʩ�	�h��@����9[^��YM��Yq	Ȑ���@����?�ٟ�������������eX�D-ݛ�Vc
��=�;[�9�[a�v�n���9��hTl��j]]�zQ ��f*��u�7|_�~zz�h��@�빠r�I&��8�x������ٙ��W�ߪ���ڰ;9�W�P�~!�ٞ��:�ۄM�Ɯ4�����=׮�������>��y�Ǒ�#�@�w-X�̫�ǅ�$���@�O���2|��P�曙Cc�Nf��ڴ���9[^���s@3��߽�9��:�^-��t�[P��*�wh�z1q��W�~|Ͷ[3q�Kt�F��ߧ�@�mz�]���hd�w%��Ȧ�'D�e���ʿB�� �D(EQ��Z�7��M��c���k+(���p�E2D��=�w4�է��=�,�ݫ���r�t��j]M:j��~J U��zl�?g3*�����9z�iؓQ$���N-޲�+k�=�w4�ՠ<�n١�#m5IQ�"K``oz��%�NP_�����e��MC!C)��SA�h�*�@���O���A�	�0ٽ�I@��*A�XZJ��a�&�!���2��j@-SL���XE�B����۵�l*J@�l�KeD��M(�A��th֖SU�`5�r�6	SQ"E5�
.�>��$��*h!�א�0��H)
D��&�!X�D �&��
 s�w��??����ؐl�-m��]�k�I5��Ā�VUj���Jܲ쮊���M�A59�g;l.���[l�m�  �kX  ��  -�    $         8      �   ���m���5��0���h
HJ��)W���җd��u��\c����s�m ՛@��t)��ٚ�H�v��aa�v3ru��A��;h�ļ�p�gbA4�GlgEŠ�iI9���v���WT��=
���u��Q�t.�p"�p�%�v���uڳ��K�ݞ��y������{Ih���9�������퉘"ڠ�O �s��کTބ��wb�g�kZ4�w�"��Un捲�gD�Ѵ�x��3I�Z�S�,]
��]H�W]B��u��PVp�Oc��&�ke����
Ɲ���Ӓ�,�,������ܽI8J���۰�R�^�Lu'm�vq�A�.xpm�rAF,�$^���������svE3�
�KX!z�ݞ#mF�v�n�F%��I����tRn�uǚ�YԾ�q�-���-і�v�[(�9�x.�n��'nK��+�h�q��= �85m���8S����M�;;�l��|c�c+U��6lI�-��B�zc<��\�����EX�v8-Td�ͧ�q^���ڍkK(�o@������˴&x�鈂܆v����ɣ��Ok�G
����ss�q�n��L���밦N��;;g�x��R�v��ij��;��L�\�"�l5[��UE84�ch�NG���!�*���\�"n�i���(Ƿh��\k��t^.1�F��[���Kci���\����٩'5�L :]'f�-��'em���@�T��m�WW"��[�Qڶn�@�L3�j�U�:N�DU�&��k��H�\��WlY2;	�C�4Yz0�k	,�;vqػv-��%��wNt�h�W�tλjӴ��m$���)�">!���  ڱU=}�}�w���?~~w�:�h��V���`k�ZY�AUU*�[p�{v��i��M�)�8���8���v5
��́a�s�6Fy{:�F8��ͮ^b�.ڼqvI�ݞ@�ny�o-����3m	g�vN���:2欽�3az��������tg�=�u��C��4&��1��;>v�&����a����ԧ [����[�M�u[s�v۶�v�n`5�#r��n�~B@\	�.M�wR����J�9fH�A���Bcgj�o>5ƺvx�S�xᲠ[�M*6�Cs1����z�n��Y��<��g���k�:��擢�6�q����Wj�=�)�r���	L��9F���N�F�ꥵ`f�l��<,��I
EVϷ�`f{֬��u�_�8���iȴz�h�W�{��h_U� �+�������4W��=�w4���/�U�~}�{涕���[�*9�˒Ě�ۭ��v]ՍQRЪ��U1�3�PB?����8�r$H���������Z��?�/�2w6�NmT�P75R�ji�[�{���ފD�@"��`��AE�*�a$*�b���RDB��g:�;9�Vs�j��!A�6s�>i�S����K�X�~,�Z��JhW[J���Q�8h�k�/��h�)�_t���:P��D�1�E#�/u��5%�,���{<�X�fU��*L�In9��Wv4=�&���)�ynwnܽyGV��W�����L��1�Z��|��zS@���/Z��w4��똡�s�*[e��ǅ�P*�g=�=��V3� ���)T�M*UT�`vy�Vw�j�G�( I$� dB�Ūn��gf���٠}�V�i��"R2F�����ٟ����;���3��Ԓ��y�U����m����6�&)�ץ4�)�w���/�S@�ũ�r7�6��?�	Mf�;n�x�m��KG���{u�۶��[�ipj8��AG��4���s�I/�;���9��S;TʚST�EM2��3-_�(IL��zX�zX�)�{��#i�&<�����^2��f�DBJg{�K;�j���2�B) �"�'�f.�/�~�;7$�Ͼٹ4
UA4 �o�{�M��j������r-��4�^�����g�@�}V�o+�@�Hvs����+p���u�I�/�ƍ|q�>v���7O"Ln	a��b����>��ۚs��]�����=,�N�KtԄJFD����4W�h�)�w���>][V8��j"brC@�}ɰ3�xY�9��V��O&{35F��'���h�)�w���/�R��%�y�`skj�v��4����%'�n�}Қ��h�)�7�#aR��ZXJ���д�Ŵ��Q��$���Z#%]���~�w߃t�Z�%U�s:��f�!�m�ۉ6�]*öS����y��L��ّ�7�c��1kv�!�`�ls!�� ��h��Ga⣦z��1� ku�$�]v箔|k���L�rl�F79:
��x�)t:���,V������1�h�Zț��&�Y�;a0��<��9����őˎ�hC��C��A���������Xܶ�6�:'� �%�:��\l�W.U:��6٩ ��ac��b���s�;92N�լ��f�l����������@�v���4�w4
��Y2BL��&�p�=k2l�^{�j��:���9;�[ML9l�M�5Nl�=,�2՞��n=,�ǹq�N)M�M*UT٠w[��}zS@�v��ҚsW(*[���2�f��>μ,��z������4�w4P���#y#hI�����.!tc��.x����{�����ָ3pzI��q�&�D�䆁��Z{�4�w4�Jhy.I:5I<b�WYw$��s�A�>0S��`�]JhS{���1e�!�� ������Ep�`meTRD�@��%	|}{���^�+�o��H�W��pi�Nbpp�-ݵ`}�xY��v�f�������x�dC��Lhnf���M�ڴ�Jh��hw2�d���li�@�Vd���^���j��:�;���ӕh�t�p={.]�"v-�ݞ6爤���Rsu����]�����V��E��Қu��ץ4Wj�a�������m�����Қ���;�)�w5kiH�&Ձ�u�`s1�e"�B��$
��U����H��U��,c$S@�Z�"�QL���ύ�n��덫ĉ������������s-Xμ,�]I:5$I6Hɚ�Jh��hg^32Ձ�<웰P�b\����9�Z�M7fѳ�n ��t������3�M�i�r�q7�$�)0i��-��s@�����̵�	%Hgk6lf=
���j��j��:�U��;Y�`{�d���d�	1��ӆ���ۚy�Zz���Қ���1E�*]5`w�ܛ�̵`}�xX(�$qb�S�3����rI�	�����bx�6�@�[��}zS@�빠w�U�}��'TNF�%��H��-�[q�Ӑlqɳ�;���[`�y�����vf4�I���}zS@�빠w�U�w���>]q�c��(2BcrC@�빿��/;�h�~��>�)�_�N�IO�I�y�Zz���Қ�]���P�pi�Nb��Zz���Қ�]����������L�pI���>�)�z���;Ϫ�;��hzeiɍHG(�����l� id���������M�m�9}8K.����(Ӎ�wV��1j�1�F�'`�q��AOPtnX�jx�7k�`�`�ua�3�j6A������݄�dy���'��n%��pTc<��v-���Y����l��bɭ���qw=�kGn^y�dwL%���V�űl�����1��s)���L��RQ����slV��w{����,iI�!S%+I���s�{�༾^x�v�8O)�g�Đ,O	.�1̑�q�6����nh��h�w4����똰�C�I	��w�ܛ����ڰ9��6�̵����~Ŏ'�#nH���s@���@�빠[Қy�X5#j@$�������w4zSC�����f�u��/�7�!1�#�=z�h���;��h^�@��F\�!@��Y��tV�Nd]�j�q����Txw^+���Nd8�pj8��`䙠[�s@�[��Uz�׮��s�u�4�'1H\��~��)Ao����m�����ܵ~J!%2w+M���\�j�nf��~�����s@���޷s@����ɒB8��z�]�޻�y�j�ӵ��`rwB���7Nb���tՁ�ܵ`y,������`s;��m�o��~��8wq�c���[g���[�۬q��q��s3��;��mfMn�{vi�6�<�<m��;��h^�@�빠u빠w���R6�0�cbs4�Y�s;���rՁ�fZ���
d;�jg[��,���i�`wsmX��) Ch�,�N��e�������HL�i��P1�l�#� 0�/��� ��f�HBH��q��"�0�
0�B�(J��+
���8�@.ݕD#N�����SFjs�a蒒`ƶ!�h����\¬��������F�#4�h�X�T!BU!���	)���!#XBj�.�tL0�
D�2J�
8��D�>�t�j��T�3@ d.�	*G@&ۦ�WXJ���)A����5���ׁ4�*&�S�!4����ANs��U�Q4�PCb�LP�6��4�@�������H
b#��h��}���'�{�n��$��q�F��f�׮�޷s@���׮��WP�pi�Nb�"�f�޷s@���׮�׮�ͷ��������b�U1
���\��'b.w<\knvv`��'57n����67l�ͨ����π����^��^��z����+#&G28�n-ץ4�w4���W�h+F������9#RC@��s@�[��u}V��Қ�a�X�!�	1�3@�3-X��M����¢!%����-k��Hڐ�I����:��@�g�K����f�ڰ;���v]S�j�6��-�ݭ��\Of1����n1�z��K�::n8m��=!R�:J�Gͷ����u빠w��hzS@�>I:Ғ�j�n�i�,�r��(�2gsmX�?ץ4���[�Os�s4�]��Jh^��:���=Ε46��cBs4�)�}zS@��s@�u��9z��L��8�i8Xg^s�j��;���^(p��������c񶹦d�Oi�״�ppl�I6��n8 �c�tJ�\r�v9���gnX�-�tW��D�*�*��B�p�c:Y�f3�o����!�Óm�[b���)�V����o:�=���nL��6��h�sQ�X�ě�ᵣS�nc��^Hy(h��n���g֛���=Z��1��g[��k��,�A��sk��C�|�؊M�ks�HO][O��w����s���lt5,�[c��lʼ�8E��l۬����~|H�ql��D�ITQ��~��4�]��Jh^���a��I�#0�s4�]��Jh^��^���/5���mH�#��_�~4�]��]���s@=�ZVF���Ԅ�䆁�빠u빠w��hzS@�>I:Ҋ!��S4�Vs�j���/no���_���s@>/%X�o$m
8��45ɜ�ǧ���6�Fw�uc�����a狴wDf[#Ĝ�&E���s@�Қ׮��?�G�����i�RUK��RmT�L�߾���+��) ����'��`w��W舙n�54�N�e:uS4���j���r��I%3�͵`f�����9MJ)ӕT�5MXjQ��=����u�M��s@�=�T��#�̴�X�rՁ�f����nhzS@�Ԯi6�4d1�/.�wW.K�țz�pe�Q��;p�u\�"��H���ɍ���:�����j��u��>���ڰ�ڙ���u-�M6���Z�I(Jd�ǥ��͵`w:��T{Jٙ�T˗554�MSmX�~,�rՉDPB�B�%$���?��[4�-�s@�+�u�4�'����B����X���3��V����`wkM���\�j��j��u�`g;���^s�j�؈�Z�����n9��Wv4<"F��jV̺S��m�/\�vz㦋m�rv�k�l��m�F를���3�{7֬�^s�k���C7'�@�����H��$Q��^��Jd��ڰ3q�`g;��H#��R�����Hh�)�u�M?�~��s@���h�Z��R ���!�vu�`g;���^�H�!	(��Jh{+J���Y�����/��hzS@��M�Jh�jo\��ȞƝMf�;n��-�n�myp����>�Q�dy������/�"*U��6��ߍ��4�)�_u��>��n<I�RdRC@��M�Jh�w4�)�z�TЇ�<���ץ4^��/�S@>���1�T�:��e���7�`f����u�a�Nn^�gt��r6�T�ܺ���)�_t��ץ4�wd��|L��zӅ�]p�I�6۶�I���7<�̝;�R����m][hŰ���s�}�6
��ĵ��&�<�ș鸴����i���G
�1�-�	!��-ѣu�a0.���w|,�6��;�y�u���ru��j�Y��ؒ^dݙ�1\n�=�'�E�j8�q���h�Z�*�E�c���\鱆�N{�N�]r�����֤jH��]5��V��d�v��4u��o��mȶ��]�;�"��B3�f�9�	�]���O�u�M���ץ4�`ԉ� rdc��:���}�s@�Қ�Jh�+J���Y�����/��hzS@�빠w���x|�u�ME$q�&h�)�_u��;�xX'{��8��JڦT�&��ә!�_t��޲��]�ץ4��}�ݝ'���3�.8�j͋��nva�n8V��쉐��^�g�И�������w���}�s@��M���o�?�J�˪�WWT�[�����<���_DB�p�*#g�7����fڰ;�xXV�Y!��F�h�)�_u��;�S@�빠v/��x�%1�hm�s�j��1�`g;��6{��+�5���MI�921��z�h�w4^���]��i�$o$m`M��uq��]��.x%^���h���`�]�X/�_ͥ$o �%1�C@��M׮�|��g�;����I֔�7��ㆁ�t�}�Ɓ�t��}җ�J&N-��fh��Ke6��j������1�ga8�B�B�(I�(+��>�w4WJ���c��;��;�xX����{�zX7M��i���tꉦX�<,ws~_ݳ�w����|�eX�r$�4A�r��X�{a�}ѹ;�s��RcQ�m��0��H�9�&ܒG!�z���=zS@�YM�e4�_�uŊ �9$�h�)�w���޲��]��ڂ)Ra�#jC@�YM�e4�g�Ug�֬����T�7T�)̵I��`w��9��V3��|���A��2!EWg|�nI�&��뺷,ME$q��z���=zS@�YM�e4�G_ᑯ��LI�∬�C:��َ�]:^,�0#9��M�i�r��e�O �ȣ��z��@�YM�e?�!}!�͵`wkM��JtK
M�%ӝ�e4���=z�h���zѦ�ɑ��8؜4���=z�h���;�S@�ѫ"A!#nG#r��s~Vv�f��1�a脡NwoM�/��ر@�$�����zsy��ܵ`u7�?"QA�)�aF!�P4F���[��&�2D���ąaP)�ւ5 ā � (1�������!cP�HRXFQ#!�������B$cRD $�	+B�*.��IM0b I�P�0�J�!��'4R��]CPXk�h�HB0�����*D4���1�
B4b)`2FFI&�f���"��q��D�!4� !! �%D$B@�W3l�(�+�viQưn̽UM�����+iT�H�cD���`��R�`�bㅌe�0v�m�  m�8@|     [d    H  l H   ��     �  �5�Nqm��^�n�wŶ�J�,���T�.��\��a��UI������hQc��#L��ƹ!�����T�F�V4�<<Ʈ6�Kv��t9�smm�����a��uf�mI�j;H���+��p�ݻ����	���,{,m����u�>`�V�[#��1�q�s��j�q������n��l��Okb���|�7]���f{t�����5US�]���'۳��n�O��fz�;����`ˑ�b8&��H�=��e�V�i,�)@Hr���ڠ:����@z�ɸ�m���T`D�n՛*���i2�Q�����v�ø�v��v�n;r��W%m�l=�j�6;I̯(lbαŴm5�kVۃ�Q�*[c&l��ԋW$cp�ϕ�ir��͆^{v�r��r�e�BEm:��C����]��jM�H�"Z�:'��Mؠ)6-���0�9ntSSp��N�n�u��5n9ƨU];sg:�%jy�q�;d˸�z���/*oe�[6�Y�5���- �YS�1c+JO��%�����A�v����Y�B����gT/h�N�TbP-IY����{mŠ:��{o[y=]�n�O'�ۜv�X���*�8|;�AO3�ש{�a����NNUʶx�����3m�����]-E˳uFGd���[e0���;=���kb8b��[z�q��p!�^��l��ohI9���;U^tW)mUT6C�M[T�!�{%WPqU/m�旖��q�y�A9�n�bP)�c��,���8�y���[���`�Ѧ�,�Z��V�vE/!lGI`�!�gw=�h :�:�]%����[Ekr�u=���{�ӻ������ q����E3@���� H#� >	� }���]f���V��,�k� 6i'-WU*[*�t�;m��Ω�y���d�ۮʦMHk{P�#�lsy��KNun������m:Z�<HMه{X�xT��6�p�����g���wbv�g��]�᫕s��yz .�mM�xH�������	/v�qy9G�p�,���ޓ(��`�uqN9�롡�������9��Oĸ2�p��f��m���t�2p��ˬ�h���0k=wn����ˎ{O<v�Iݷr����P�5��8�(FI�8L�)�ߺ~4��:���*�W����v�ȔǑ���4�w4
���zS@�>I:Ҋ&�r9p�:���*�W�u�M��4���[ɍ�RL�9�}�hzS@��M�]��Ҧ�N!@y&8ӓ@�Җ���^���j�3��`s(�X�Ғ+�iȥMK���L�YGv/'��-�nA��k��q&Ӣx����nfPm�c9ׅ���Z��q�Q��zX��5�D�B(�nF�4�w4���;�xXμ/aB�;f�R��T܀�� �߿M�Jh�S@��s@�v���a�$iɠu�M�Jhz�h��@;��'cY�(�9!�^�M�]� ��hzS@��F\n P ,�4�H�؈�P cW�m(�(���lEm�X�*�&R$E$R8�u빠���Jh�S@�+�u���% �ȣ��ֻ�ׅ������u�z�Q2wkM��M9%�&�:�݁��K;ׅ�-(�dd���H2,� #!!0�!#��0��#! H�H!a	"��V��@���UCz��g�rI�}� �։4�L��q��p�/t��ץ4�٠u�M�hՑ ��F曪l�;�xX
""w���3q�`^빠r.qD�X�X��/�p�Nն�Ŷӻ��^ݺ�f��/��ht�ݱ�ڣb�����f�ץ4�w4�Jh��B2L1�$NM�Қ{�4�٠q���1Ĳ
0�Hh��h���f���M����iE�H䙠w�W���}��o~����g�Q�0`�qv��s_o�|7$����U���%!$���_[4�Jh��h��9���o$m��B��sR��c���2�[u��l��������v[�'�щ�($��h^��/u��;�)��� �Z$ә27�'�]��Қ��4�Jh]F���J8����{�4��i�%
g��K;�j��L�)R�M:�Ф��}z��Қ{����M�ڂ(FI�8L�rM�Қ{�Ձ�u�`gq�LJ �!
,�{���ȶD�K��A[�OZ h�t�kn`�ٯW]�B힝�[\p5�8�k�nz�ܦϯGY鍧f�FxRf9A�5=T<q�9�,��;r<L
��^��q����{N���u��nIȝ��.V�k�SŅ�[x̹j��m����t&��':<c[!r&�oU�S�x��:�(]���8��X;Y�9)���1vv�� �eʄC�5m �c
��>�u�V��mt��x����չ3㳺n��Љ����' �,��$����`w�xX��~��#�n=,²fkje˚�TܷM�`w�x^��L�75��g�@�u��>��o&7�HI2D�^�@���@�u��;�)�{��4ъD�Ly&Hܚ��Z{������T$�y���37J��i�4�m���6yܵ`l%ܽ> �����˰�"Ō�p�HDޭ�X��d'y�g-gu�.c�]�^��߇�v|�P�̉FG$ng�^��^�@���@�u��=��C8��RC@�y=�7�AVA
�VYϵ�Z�����M�)#$1�c������`w��Vz!D�w��_�@>�+I�2$AF9��빠w�S@/��@���@�|�n���K�n[�L�;μ,P�zf�������Jh��݄Q���(�?�̑uH��G&��T�C��A�+ֺ�l<����o&&%!$���_f��}V���M�Қ�n�M�IdǒdP�h^��;�S@�t��_�����[���NdȜd�4�4l�h�Ϧ�PJE�xE\�j}�h�)�|��Y2%��h���٠}zS@��M��뒥�SN�0��`�1��B�������;μ,JY�:�:�rg�c�^����ِ���F�p�״
=`�:']Wg+sDThN��4�O��������;�)�ų@>�+�,�IL$�wJh���٠}zS@;ܚn��&�n)$p�;�)�ų@�����Қ�]C��R�F�Lni�;�u��zX�o�ќ �
�뿞6���
�.�Y1�$�ץ4��;�)�ų@���/�d�0DMdk�F�hr��n�ͱ��N������f3����8�$i8h�)�w�S@/�f���M��jȐ9�(��C@�t��_��ҚwJh�Xw\X��Q����٠}zS@��M�Қ�:R(FHc�2)$�>�)�wt����M �-�}LLN����I$4��;�)�ų@�����y��޷���q����������I�6۶�I�۷M.�.af.*kk:v#�F��bȶ1y�G�|i�'E�]=z�{N{%ԏ:���Wmp�6�Zs����϶4&[۳��=N���V�6ܻ�Iգl7���$HD��������u�/)۵ne�nѣe��.�"�ZA\Ip�:���P�	�g�4��&'p��py\OV�_w��}�������|�iz�ȞƘ�p��*s�\F�.ȶ����}I�Y���D�r��F�rG޳�ų@�����Қ�]C��Ńɒ88�4��h^��;�S@�t��B�S'{�j��R�̦��卻�g�@��M�Қ|[4�Ѧ�I���$i8h�)�w�S@/�f���M��jȐ9�(��C@�t��_��ҚwJh-�q��J�ힸr-�Ƶ[]��q��:���8�m�Q�릾���f��^�Ӷ�$<���{Ӎ�|@=��{�9d���i�t6���B_/���P�|�IBL�~xXw�2� ��&'`ɄIL$�wJh���٠}zS@;ܚn��:��9�N�a�B��^��3]��vS@�t���WP�y1`�d�' �:��Қ{�4�Jhy+��:N#i�B�	��%Z��3nva�n%���Gp��茥��-r&‶z�-S@������M�Қ|u��h�S$��c�$�4�Jh���٠}zS@��5dH$�#�6�����3�c��.)q3�!B��[�^(�)|@�M��fPP���r��4c	��	tc
kui��UY���_��h4��@��&�����p 9t�3���.��<`]e�g�H�`lA�¨@�E�9C�9E�­BA���Xlњk�����;����;|�/��9B���E
ZB�%�	X��0Ch	���3�F)C��*�$>CD,R2)
��0d�\�s��<��bI�	��D H�|� H�!	�H ��a�IBbol���Z�B�FH&��aD��J��k),��b!X0*P-I`�6h�M��J\76��Tt�C�)������E�b� !�'��衂�}(�|z d}$��/YM���0��`���_��ҚwJh��/��H�2d��c�@�����Қ{�4��h�Z�֒7�6�M�8���b�#��nyU�����{	�V�M�LNA���I$4��;�)�ų@����wri���#q8ㆁ��M �-�ץ4��>��o&,Lq�D�ų@�����Қ{�4���4b�%��ץ4��;�)��x�i! "W!U"�b���� b�3���n@���51�7�'��4�L,8f;�������ɩ�eL�`\���Ӓ�l\=�&{OX�q�aY���)\j��p���rT7h�4U�6�~���3�c�>μ6!%�f=,ȃ0���r70rC@/�f���M������B�7������-��94~��w�S@�t��_f���#�0�QG�Қ{�4��4�Jhw&��lQ��7$p�;�)��Y�}zS@�t�ͷ����?^����՚���gU� 4�m��I�ʺU�ns٨y嘀W;6[�'���?ӧ��>qL:۫�m��u��ť�.yӮ�6�ȴ�ږ�U\5]��v�(�qv��' ��yڰ���箋�;��CŷV���.`4Rȓ�@���nt���7c��wi�bs�ԁ��Me����t��6�Ri�r�	����<fuf_Df�|ƞ�se�Ւ�7O$v#�jȝ�,��m��4�9zc2��g�8�p����>�)�w�S@�t����q��I@y&E&���M�Қ{�4��4�
�)�DێH�p�;�)�w�SO�G�/�{���˨Ց s�#�9�Қ|u��Jh��<���?�F�Hh��h�)�w�S@��M��uLNF��BD�B�ۊ��#���ix�<�N�;��]=o&ж��r�DXLs �Dr6��/�S@��S@���B�@���9�)�Mk(hrK��5�rO<�>��u�JЃ�#�b`BDO6�=���埍 �����Jh��M܉�q�#��}Қ}����4{�4�C���&Eӆ�_r�@��M��M��4����H@Y&E�@�����t����M ��f�Ջ���m��4�[���gg�u
����Wbݠ�9N{\�c�6.��(4�9N8�I�@��S@�t��_r�@����˨Ց!��(��C@�t��_r�@�����t���`wk$�L���Vh^�M��F�HB!M0�Q�C��Ł�u�`ga��5M1H��mI�}zS@��S@�t����P�w�:�n̎BkYC��m�,{�4�Jh�+4�JhyF^΅cb��u\sA��Jӈj7lmv��ۨ���tv�^�I�[��v&Z��;�)�ܬ�>�)�{�)�}B�Jʤԅ0rɩ�Xs���D%'7�{�K����B�9��i��]<I�F��=��Ɓ�t����M ��f�wZ<mLR&�rD����s���:��g��!B!	!@��	a �#��S����
�^�W�vnI�ߍw2�sXWQ�����M ��f���M��M�\]r6ȖC&bBF(Ԋ�{V�́�wc�������V����'im��\I�9S$4���ץ4{�4�JhΔ��)��4�Jh�Jh���VhZ�'a�(�L�8h�Jh���Vh^��w&���%#RGQ9ܽ,{����:�9μ,�C���X�Eӆ�_r�@�����t����M�g�Yr���I$�2����t�l U�s�l�UҭU�\b�)N�ܥvݮR�o`3�b�{Zy�<+9���mt �
�!{eQ���u��.p��x�v1��w[�(-�U��^wS��%Lu��h���Z(7m׮��p]%��J�BJ6�.�;{nWlj��cc�φ�WXzI;6�W;	�U���սG����	������r��`���b�;���{���p|az�DLB"�K!�9�͆C�kn���G��E��-�cBXݖY�$�{]Wͷ����|��>�@�t��{ܬ��*LR&�rD����>�@�t��{ܬ�>�)�r�ȱ(�'QƜ�@�t��{ܬ�>�)�}Ϫ�<���yD�r��-���$��{���������U��@��)&9 R"9Rh^��>��h{��{����.��±�O���";e�҆ջb�m�ƍ���\�rzt�.�5�k��u��#���>�@;�f�{ܬ�>�)��M7r'�0JF�R- �u�fg�!%�IE��s��vf<,�]ɰ>��o& p	��@=�Vh^��>��h{��>�����c�	M�.��IBJw�zX�͛ �w&�{ܬ��*LR&�rA'���`jI)�激;ܝvs������A��u����ա��OkG]�Nwn�7I�u6��݁��/��8��A��d&jH|����+4��>��<�����s&194��f�ץ4��Z׬�=�jȡ1��GM�Kvs���rl�dvb!!@ E��P��5�f��=�f�Z�L��B&94��ZW��{���)��M;�8�'ڑh^�@=�Vh����}V�����^�1k�I�&:W���m�d�8�κ�c�9R����B;�،�� $II�{�Y�[Қy�ZW��>�G\dj1ǋ�jMޔ��E�-��= ���@<Z�q��M��Ny�ZW��z�4zS@���bQLN4��r-���nmX{�������⨅DB�]��a�Ą$<��2011FHH2R0$I$�I�8 �_ %o����t#��!t楔�EM:�s'���z|v�f���zw+�@���1&��za��M\��p��x���5n�I�-��j�B+2��)��4zS@�>�@��z.ꞁ֥��1���G�]ɽP��6w6��͚�3:�Q	(�wf���iS���DԷ6��Ձ˸�@��4��hp:�[Ɉj �%$z/uO@��4Wj���N��Ձ�㭧C�tS�*[T鹫3��B]�ݞ��,O��Ձ�EW� �
���EW���
�PU�AU��EW� �
��J ��(�X*X*B
��� 
�"�A
�`*A �A
�E�������� *
�V
�D��D*
�F� �@H*P��E@���X*F
�Q��D��`�DR�*T��D��R�R
�`*A`�DT��DR
�@`*@��`**�P��@
�E��`*P��EH*F� �AX
�P"*Q �A��A��@T��AP��B�H
� **�A��AH
�  *��"*R���@
�T"*Q�� ����EQ`*�D��E��AD��E��AF�X��`* *T *@b*`*U * 
�P��
�Q`*Q��@"�`��B���@����E�H�� 
�UH
�A�T�"� *E`*b�� *D *�"�"�
�P ���U��AU��"����EW��
�PUx"(*����"����
���_�DPU�"���"�����
�2���q�8f�����?���������[��,7��U@$�I��        �
 PIK܀� *Tm�Ɩ�i0m;t�I�f[p;����(�L5�飓�. UE�k�t��(F]ƅ�dp�5���lv*�w:f+;�tv��  jB��t�@،�6� P�`;GNݍ(�'v6�u�-�, �:E�Փ�v�GF4�d�S��9���l�$h�� P�cNd�u�v`�#E)�YJ�tt�4қdi����@
J)  �R��S��'����@        4���@a0F@4�S�z�B%D� d�&��O���I�0� 1 2	"&�M 4�biOș�M��h� �E	��P  2  p���-:���h�$��7j�?�`�!��b�(�@���%�6|>��0@�$H�Bzq���K����3@���;����ʮ��{W��c��<'y1+��-{rB }�A�H(
��S��1���%~s�?DT�P�>��lC��i~���_et��|`q�pDQI4FfJ%Υ�uG��[�t�z��\���v�ݶJ���Swo ��^"�h]h�DM]�^k@�racģ�4�"���TJ-c
�6���h[jb��-)��ah�Zl]�DDF�O'9\��y�O1^O<�'�UP� ���y _"
�U|���ZL����,���Zl�6%l���e�-����K�ݪ�o#\	�n�:�Yk��k��kZ�l�f��Ұ���W�_z���wh~@��6r�Jƞ���C,A3rrOS�BUnգ�V�gk&��������Ӑ.�Gfi�
čͩ�UW�# ��o��u<����о���D!��	�;��A�$uC�a
�	B���	BiM��Q"a�<!8e��x�uN�ąX�M�kBzj͈(��j.idؠ5F�0H:�n%��5�(Х�z  eW> <֧���4�<P2��&$�̻eY˔!D,��
-e��Nr�H�hF@`�1l�HU�J��k[�oG!�s�.�R��I�]6m F�D`T�XY��E��x�
	Zo89��R�e�i#!�5wW����y��k(�	��D# �E�2b�k�#w��h�&���9�cM�y�A*�V�
��"���%�hd	�ssF0�M���� ����&����3�dP�J(0�y����u}6�Q��ݼ%]&66+S�L�I�ͫf�y�R$ݒ�0��:�"�ЂP�"$"�n������d4oC��F4ـ��wk
���[4p�SF��i,������Y!Af#�l���v� ¬�5�F�p6 ��15c3o�a�)�ZB�0�`�L ��RE�ѹV�CL�$T^\c��E�t����B�0�4i)TL# J�����5����u[�Cp�=����;]���Jr̦�m�;=ҸmsC��&��3�F�s*��[�jUhy�[�4�&��΋nؑ{����e���Z7��l�li�ٙZ�s��Y�XpP��D&�Js,�(L�9���Qh�v�v4���I&�*X�2+J����EAb���Ut�a�b�-����7�IXX8�m#-q�MY�:M�?�Qn/��j/�_�_�]L��             m�    ���                     �                                                               �                                                                            �x                                                                             <                                                                             �!�                                                                      ?���<�U��Y�$� h�WiӴ���m̴��M�&Yd� _V��u㭡�i=k�nÚ/'@[M"�����6H��'TTn
��@m��d��-��m��5^Ù�bY&�u�#m��ECj�Ö�ӷm�L�	�k���M��m�nѭ^p�$���n��-��|�x � �  l(  �m ���  �6����mU� v�H ��  p 	6� �k֏RY�:J�	���/�e�*������r(����-�u�&�[:<q�p6��ڽWi����u�xv�[��l8�v��mm[&��mf����ÿ�y/������(��8�z�6�n��[��"�`��'���d m� 텑�Ui�F�v��n��)[��hZÛl���Cm��m�u]��M��m� �t˶mrD�(�i�6�tmk��6��29�N��:^����Ӛ�<��ie �Y\m�[@�6��	���Y�	.����t�o�$vd�m����ە�W(��t� ���'+i)��kY& 6�m�qm�]m�ە́ŭ    �6�mn�$ ��` m�$�����컗a+���V�^6��v�7극���6��rF��e�B4Y0�.ƛ_�y��Yg����Ͱ萓����<� �e��$TN�d�ݮJ��H:��rlLP:3�hܶ�6�U�[R�Ry��w�1����V;lS�{$�����r�M����Ppo�}�������k�Ve���f9�ln2e�-��E���і�,��(����찳~��d��6J�C�b&Q���[(6��Y�H80�͝/����<*�ԁ܀=��9ٚHua�9H0���6p�#D�8��pژ]wy��n��
5`�hc���Q	�dJM���ѝ���qG�������we��n1���"dy:�4��9H�A�J�D�����
��c��
eW��ӖF`���m,!}�f�	���K�"$�w0'x�:u`�^طF���ؿj��`FH�~Dp-� `�6W�Px�
 ����������5��'tQ"�I��q������i� I  ��6�  	            ��              l              ��              l            � ��"k�	��ܖ��zu4*����хi';'[��m�����`a$�P�7m�����[�j�MR;b������B��iUR�,�@�^�K"��j޵�K��YD����e�j�T�+\t�,�X��K5 #m�Rb$ň�V6,�ֽQ�W/f����Kt���ڣ<�ȦP�
(�|V(o�=wi:�o���Z��������I  m� m� m� m�  �Xʙ!eec�;�4��BI&�P^p��rW?���{݅�ň��j�m��m��ml�KM�	��m�j���;��EYU�ai�qM^˙�z^����<	�32�_~���?w� �P���*d��z��/ԫm���4#v{:��������*׆�K4��U���~��~���<���  /
��X�����v��=qKng���vO��l�{W��C ��׀�_���f{����˶�O�=����y~� \"�G(ʴ�-��a�����ior�0��Y<94wo�.�§ե�e�;��k{������3|Y�گ��`   �����%��7�E+�ft���ـ�C=���y*�[x���3շr[���W�n���-�
����:���Am              mۖe�ǭ,�ݲ��ɫՕ3��Y�MsD��]E�{�y^]|  ���F,JY��ro�벹�s����ςin��^�޽	��W���u�r�=�w����u���<     :XT���X	�j��C����g;Yt+��z���{��.�[1r�d�]���3��}����-2�����~���  ��/Z���]�Mnн�8�kКGv�.�{nAL��4���K����{�V���9��n��l�>�y�{����Ϡ &eζЂ��0�bZ]��^�7�}��e���X&��[{�Bj�o'j��%����+�{˙�����    X���w0�g{�noe��9�w&{�r�\�vjp�)z�fЁ1�xrh�I������r[n[n@             m�o[��i��UѴYwh�2�c���¸�il+��<��'��;�;z�����  �Ze �e�-0U㫩�|f_�����y�5/kЙY�7�y絠�_����{3�no��{N����{�    hL!d �&e38��i'{}����y��M��ݙ�=|Ze����~~�κ������=���j�  @YBWD
ZQJ�{�w��f�9]�[\����V�K������
��:��U�R�L6S+
��4���PH��@��H2��4)yVVJɋ`��p[(�q �X͸��=���9qw������X����R�q���F=���<"��r|cY<3��\���r���waV��d� %���ϟ>����g�w�  &�[wD乒��=�3�]��"n����I�����˙�ςk���;�7�?����~V��ظ, �ݿ���L��k���߿� �F�ݩ�jt���5��f�m��nWN���t�v����U�Z�^w�&�>���~�i2��>�~�ޟ}���'��l 	                 6:8���&��[Q%�`G�-v�:���"n'��haM���S�����  D�k{8�c��?_��ݳS>ס2�E^o(��~��S/������Z���ʱ�;���-�����{󯞾~�<�@ M�[ۛ�JS�媽�ڢ3.Oxrh�)���x� ��|g�t��ϚL��]׺�h�~e�F�׽�}�BeXݼ�Y�9��7� �ILl׵:\_r��緾Ŝo7�����_z��Kr��M0�@b�� |��s��.Z� ��{�� $n�9޼;�e�DK��  ^����^�X[�19�>e���=ӝ3�|+{�;2�{o�M��zx*�4cv�j�[�E�w�߽����    R��`��Z;I�}��=ò�}��fϮww��'$>�W�>���ܴ�W|�e�qh�=����f�O��w(��/�w��d����             �n]���y�gyW�5�LV����k �����l�R��$��Ǻ   v��^YW]|��m�����^�DHa�~���Sj����'��I�ZzmƑb 
͑���/�[�c�B5M��d�8B�k�\��j3P�$���� M�u��T�MC�qQ�CH:���I��8�>L+ٳ�Sx��7X���!�_�̳�8�պ�J�#&|܆��N��ƛ?jf>�����Y���S�q.���ɿ�  ��q2t=����GS2��(����f�\^���nU#�" �]��(�e�_�\�wP�^:D���"H�߇�
�o(�$r�$ߞ��s�ܕ~K}�{��y����    ���:�ؙi]{\Iz(�{h=ϭ3�m���mF����#�6��rd<_>1Gu���ffd||��Pw�nv��,F#�ƞͻ�7��y��iM-����q�Y��ܒp    ;�[��on�km��o�miB ���ɢkrp	+J@��XB�z�iȣ�!���q5�|�44@f!܅�8P9U��6��D�6 �`��r7?3��|���j�o�9�n�*�g�B��y2���C"�c"Ģb����H$Bx]�(�gr�cF�,!,�Bـ�7��#$	A
aL�bB���\t��CY�)���΋:Q�L G�Hf��-�  ��  p                                                                      ��x � ��%ݪ�sջ��3D�tӦ树�ln��L�7B6⎩t��6ٵ��L��mi[-�9*��$�*�Sp@R&�~������"��֯Vu���;cN��9[+e�R�;��k�2j�-�:�d��,�7e����9%�)9'TX�u�λ����PH
�IO˿����K�ɭf���:�/o�s���PqѰ�������=z����y��y���x� �@�           m�e���a���hYj���0dz(��HP��v���\X�ߗ_� Utf�C�OM��X?5iG�A>[����S���<� SQ���#��۸[��q�&� ����isP%�	��sP�Pu��Q�u�raP�Q� ҇3��mh  @��nK�z��|<Ҵ�'P���	3]�̳Xx�?Dl��FE��Qzͺ�NAJ��r@w,7���0���o�Ne���1�QH9�V{�-�Fݵ_���]sϝ�    4&��L�� �T�Lʻ���:��� �(�����;��@��&��0��g�zj������J-���Rcg�
P� E��sw�`k��9�IUx3� ����7;�7��su���]{_5�=ik��>��\��ɀ   j���8cgm{��{�w���� 0Dj����j�r� @D���.A=�S�[n4�$��ܸ���"+��-�u��B /�#���BlJ��� (�
i���h�1:E��&�>O?��  &�[t�&ѷJae���C���3��e4�Q~p"�r��:j���,՞"H�U�܃<GU|܆г����w�b#�"�o�M��� bG�#���{��ޮ�?���     ���      �ʩJ9XBR�jd��%vEn�v����u2�K@��{{X�I">=�  =4i���5:m���?j�fc�|v��k�\�y�Ļ�d�A`����8m�4״�h
Ն�
�i� )�L,�D�q�O �/��!=L��9��sG�$� �\P�K�3  :&#K3���׬y��Oz�3�V %���r@n��  �K�L�D8�C�{tګ����A荸�d�N߱L��d�"H7C"3N_�!�T8� �T�r�6O�����  ��{vɷy�)��7P��1a���Ʌ4$�/�#� "���nϯ�M9�4�f( /q�PwM�5f��^ �8��GכֿS�|2�����%V��ۯ4v(�G���    5 �2�[��]P)�c�(���A��k�g�~���{>���}���������-ʡ���8\���-ހ��㜡��I��25DΪ�,k�*�L�5�m���v�e��    DБ��h7��,���r%��zꊿ|��4<G� ��;�i�����t@W��Q�Y�h{��2���b�9�g�=��i��7W��������;��޼�y� h          ?�<   tu�:75�2[����f䒍�*��~��n4Uh��K��  Hۉć�z���x[���&���a	��-�� ��9G��BlMv�54hv�#H�b����ӑ����r 7f.���,�f��/�ʾ�k�֝}}�   1��R�j�28@:n�-~>�������xJ�y��TA�]�J<D�''`oU���<�^IW.����Gau/��c��V�Q @�E�t��äM%�-�����DΘ�yE�^��  ��[59u�/TaG#1'��SNcN� n���g���hi��)���£���&�Hp�Oz�II�0�2�e�p�`T�D ��*$" 1$H ĉ#H�by{ɽ걎依�ٚ�Q���6D�eA8(AMk�7�8  `x�D���rQ�9x��<9u�)�C�Fb�yG�4}mz@ f����x�y�m�����3F�����P�@M!���?����Щ�
�,#
�ÓF���y�|E��s���ޮU�xy'wϗ�����=����@ PJ�7%�2ܲڱ����|F�3n������f�F�p����t7P~�LI�C>���G�D�/Mׇ�r���#�{�]j�ҚZ��˭���	               mۖe���M�R���,�u�e���[��v�C7��;y�x  rA,�@@��_�vu�My������c��\ #O������6�8�1`� �ۯ�=���,�c�O��C5J����[3*�V�лk�쓓�  ʭ���o<��{������é;9�9���K����^pRD m<� �f2��V ����&�����~�G�S��Q�Z"x��G}��ѦwQ#� .#��6J�t�� �Mt�%֮v��^�� �36"�QU�2�"�
��Qg�*�܆�u	��" 8A�����]D{�f!�7�7֟�q�hZ�K2.�%���{�    4&�ZS"g��7(e�&����vx�x��.Z�>�b�#� ���ɢ(w(�OB��Q^�6�}�.#ș�� �������Y�8�芜��i-/�  ��1t�?;�y���u
���g�t;V�i1}�]�'�[n8ǩD�y����ɵ���_	^A��ƀ��:X�d��is+k�<z�*�kK߻[�m���              d���5�9WE�n�^:m%�)U��]:EJI!i���P  M���.)�nJl��Q�q�3_�Am��8l������>e���zb�#�Tے�;�5�yT���}礫��{�{�W�Yɮ��w�    �Ie"�Q�;m�5帖a�vMo����VN��ʒ8T7`:S!*��Sd&���h�&��DC�y zz���ͅ�?<�w�n��S�b�~������� ^�ifr}�ӦY��
�`�"�|܆�1���\qE}���]�Ÿ ��:"-�F��Ԟ��`�"A1���|�ZM���w�ޚ�:-,��  �l�p�n�rf��~�6�x0ǎ�Ϥ���E�1p#=|i��"L\A�C1f{ϙf���@Hˏ�!��D�p����|G]sf��{"�I_$�su�5�,����   z����o�y�K���-��w.п�<���7e���q��<ܪ@r�G���HM)���M��p�y^�4;�|5 f #�o�xzgr5���h8݁a ����wU4'k�f�6�1��K)"@IBOBo���     p                                                                       �nmhi�n&���Ҳ+,�Ѳ����)�l�}��km�6��m6ӝ��`I%�PVUDڒ�b�Fܶ)4�4ȭj�c�������Ӗv:�Y�ݒ��洕��n��*�5�i\��.$���2^em�m4�9������Ҹ�Iiv�W�����XPe-�=�֓KZY�k�xzp���o ���(�QBo�������m�-�             '	7hѫ���,�Ymޯ[3[�9�m+C�d[��   ����Q X	�`��[k�{�&7TU_�2ʩ<@W�w(�_DD�k�|ܴ��h�ψ��ڰS.�� ��#ƌn��Zz	i�A�g�f(]�� ̭��F����:�U� 9C�E������Ku`�&�I!#��]�p�n�C�+[󲭚�uQx�wW�St�u���o��Y�<c�Tj��.�����|�7� В鮫V\]� �'{IpI��ĐI�J�H&�$D��뤫���A;۱$C��%�$�(I�9�K��J�w��t�wy0�$�ؕ�MQBH��)# �vt��;���.	 ��ؒ	"s^o�U�SPI=bYK��D��.	 �yv$�HH��PI�]{�x�2$�H��&1Bb�=���ĐI���$�r�RA$OP�w^�1� %ʺ�qEɬ���pI�˰9
�H���	��PI[��$�M�����F��ND�$�j�A$Nr���A7��'��$�����r�SPI�A$Mn��
�y�ؒ	"n%A$yϷy��"H=�Q9�K�H����A$NĨ$�Yɜh]�l�$D��	W/)�$�w�bH$���t$�v�D�J��R\N���]��{�����@ 2f旉1���%UԻȒ	"y�fE�ue	 �'{IpI�.đI�=ߜ�Uu��A;E �&3IpB���ؒ	"r%A$�u�e��Ȓ	"w�7�L��I�9��	�)I�1��캚M�$���X�	"v%A$�(I�9�K�H$׺�.$D�J�H����rĐI<��$�s�f �&��Ҙ���w}�$m�נ@              �sn�tvg[rN���hX�J	�E�5`W#h�����sKZ\ĵ�t�K�ο?^�   l-��8&ZW_t�֓kK���[PIvR\A=��>%LD*'"TA9�{w��Ȓ	"w���j.��bĐI�*	 ��RA$O}�^�^SPI�nĐIq*��{���=�*V;�*	"��I�;�K�H�y�X��TOy�zUc��A<�A$.5A��$�w�jI؅D�J��oJ�/��  ����$u�X�1u�K��\Ũ$�甗�Mf�I�;�K�H&ꄐI��y�u2��H'{v��w�i��m11���PI�A$Nf���J�M��Iwu�� �'"TA5E	 2'9IpI��ĐI9�ۗ2��H'h�$D��.	 ��ؒ!$����M�>]� �'9IpI�����D�.	 �����t���޽<�~_� ʭ��0��N�!��&֗�Z��ZM�*	 �QBH$���\ND����s�U˹�*	!��%�ԈTtP�	"y�K�H�ʻA$O5��U]e�7�N�BH$��R\�'����`���"A���!�H;j	�ݧ�*	"y��	��xr�TdI� TO<��$�k�bH$�Nĸ$����(I�<�+�%��j	 �yv$�HH��PI�;e	 �'9IpI�e�]�1� 	6kn�ӷ#gM�W�H$�ؕ�MQBH$��R\A7��$D�{���̦��	�+0}uN �&�IpI�˱$D�%A$��ۼ�ё$D�).	 ��ؒ)"r%A$tP�	"{�u�U��:�I�]��3bH�Z�ؕ�O(�$C���o>��~�H��K�H&9�t�r]�j5�9� �(I�9�K�H&�vrS�t��~�O�@ N�"&�^.J�
����A<���I9��$�y۰�P �D�J�H&3u���Q�$D�i."�.Đ�	�*	 ����D��|�S)�$�w�bH$�ȕ�Bv�A$M���A&��ں�Ȓ"v%A$^�vP�	"_i.	 T�$�H��|�ܸkI �	�(I��򃝤�uBg�,I�1ۭi7�/�z�i��۰	           �    6�α�ݵ�CT�],Y�ʢ���+pH���kZ�}r�/� �3�]3�lb�eTВ	"st�$A5�v$�H��PI�$�f�{���^SQʂv�����H��PI��A$N����	��%\�Ȓ'�*'bTA5E	 �'{IpI�.ĐI���*��)�$���]F��&����	�݉ �'"Q	��R ��+iӤq�no�  M���.[���W�#c�B��q�wTo�Zrҍ6�b@դ
�2�MVy�,׏y��5�$�#&u�mE���C5G����9SZ{�u܋m.�.7׻�    4R8剙�'�e��n4�RA�3z��$� 9DyU��NR�	�?:<��{������BYn!{��,�6;K�'��bF"� � �5�`c+ܺl�`ŉ��XƬ	Va%Y�YX��/��h��j^�W��ѽF��*`�i��e���:��њ�V7�_\�30q������\ib�����M�������~�����|���  r�\tB%�+�mcK|ʞO�fE���fL�@w/� [�<B�0�}�SIЭ�x��>�z
e��r@�T}�Q
"&��]�hI���
�Zc�Q�g��P  z�:;vɷݼ��J@n�5�J2Fc���hv. ��q1Q�56��y
1�+���O(�ߟ�f��@�5yF�s?72fP�t�X�Z_����>�8���I                ڲ[z#�]����t׶�9cw��kΊm�1��Gn��z��zy=�~�� =RFe��}]P)�b�\aG����z��d�<h���b�Vބ��� &��Q�&��9H�f������-�#���;�|��ׯ��@ (�^H��uBS)	�"���*��̳C�\"/		!ܢ�ɟ7!�<F�B�F���Hߺ�ˡܢ���CӏL��X��ȗ�d�����     �H�0l,Ig4�ryi�ؚ��� 7U�[H�#x�KF�j�<.�"�*��YcSFD�!7P�Q3�\����/�ڽ�kt��?�@   _�f���r
8Z+b_}6����������S/�w(�8������)��H�&H�BeF�_�MP��	�;�ȼ�P�~zixtv����U�����;���~}  �idD.KE�ѩ;�0�#�7T_��r�ƚ$���ڸ"��ґ�	��r�#&|܆����/:D�G�vP)��v�MÐ7�0�T%
2A�k9��� [@              �stY)wmР�u��9�br�rk�uz�lDb"��5  U�E`��@nW.��i{�s�^�y�#N��&��Q�����k���Bm�.�8���x�h{�3@�VA��cqEƖg�&����    ��Ӓ�nYeR<@�CuE�U��6�ݶ�@7T"!��Gv1��|
e��Qu�i�:���q��7U�X�u�`I�CHHV��Uc�x������ =$"��k�+�6��~�%%�aC�]��hn(�^<`n�����*�a��wr�W�;��ev�b�5��YT *��(KW�dߛ���޽������{����|�@ *�)]Xr�v�&�ر�>�/o.6�N7W�+ w!��}~�2�qiGr�.4-/�9H冱q����@#�K���v=��|Ǚ�Y��9��   $٭�Zuѷ.������zMՄʉ���YT4�V���-;y��m܅ڎ�0��kAL�Zn�ȓ� n�ӏIM'z�؁#�q�Q:��#7ۚ�)��FG��)AƎ�b(�S�#!
�J �Ƒ���,�%2�	RB�PF���(�:�\h��0`ф{*f�fRS 8  6�                                                                          p Y2��6˦�ٝ�f9��F���n+G�F��ƫ��m��ѶƊ��.��m�ם3��ZȢq�ږ8@n[!�h#n(��X�!%#��8:�#nT�sE�u�G��2���f6��­Q�կ6]�%L�\��m�Y��/�)ח�#k����R��֮��Oɛ�Q�X/�D2/���^��;�d���d����             6��f[�wMMv��6[�I�v��̣$��nV� Ԫ�UK
xDb��` �L詩�Jt��G�]�=�0�!T��r��] 7P�?s��-C�FbE������-k@�B�C�笲�i�v��de�����  t�uk�p�rB��C1F��i�o�M��  �S �i��IM'��r@�B�
>��2�Y���tDU5���{�gyu��.|�ɀ    �R5T��BTQͮ���=.�'�jaLn�l�F�1��s�YT4�v�� ޷FTw!�X܆�h��qGr��
������xƐ3|�_,���� ze�2۵�%4��
 n����oAL�G� �����Ʃ/5-�܅��}�4���nS��Pf��5K����^�A7�E��b^�Y��׳�    Pe�Q��uͬis�����w!�7!��W��i�W�T7T+�4����^��N7Ub���:�_l��t8�B��Q���q a�|��             nKn����p-uv�[���V+�V�]�.���wz�4k�   i�'�l���o�����N�Ճ\�Cu"+�@c^g�rh��{�a�'�aꉿ�ZL�@�CuFv.�Z+bY�M��2i7���v    ��JKNډ��-����b�9��;�^��%[�VOd�&�N�P�9�G�pU�v�>�2�"�t Ҍ���y��h��0%�����qfLk2լȹ�=>   �L�^8���=}�}i�����&��T#n��Q��Ukr���ꊦ���Ge��1C;�h�wY=��iP,�B�w�'fS��@7P�Q^��  �[q	&�Jˠ�S\{��R�U���$�͘�@U�寅9)P�C�����38rh����1���Ș�C��i2�����fMw�{I�Ǘ�   ���@�-5I%Kr@w!6��@$��M������C�ωS)�w!�]����)�CH<B���Ü�7PN߯�oz{���khh             �N�d�+9)h!�� 
[-QId�t��I������=���� �s.�CLի�/������.�V��ј�B7P�H���i2�ER����Usru	��G�?m�)���ϲ�����=�����@ �b"�M�7,����"�#k~�z"�t$�r���R:��&R#��j���H�;@��U�rU��Eڊ�,�3Y�k2��Msoϗ�    �V�e�,�ݭoqw���{ܿ7!����;���/���T7P�qWi���JCx�cr�eح@�6n:1hB�D�b$d`��_����2]o_G��dh� ���X&��ʑ�Y�}�@�e��ЀQ
�U���c�S)�j���3GuD���uM�c$"E��n�3  =$"��C�W2w~~^v��B
����f+H,@�uYxke�� ��.�Mu�I�C��7PV�ƣ�^nC0N� �$x��2�*�� �m��ƣ�����Q��}��ӯIL����3zv�ˡ(f(�A�^r~ w!�����W�����>�8����
�W�/�M��             �n�Ѷ�YL��Z���n�"��q�1���[%M�r���מ���@ &�m�RM�6��;�?oF��&�x�ff�C1E���ru	�(��\
mP�Po��;���\�̋Y�����_o�  -�Н �
+9]�m �����b7'����k>!p
p��t�B�K9(�ǹE����ᩣ#� �.03+�Ɠ.�1���ݶ<j��� әͦ��f���5�U���D��J��Sj�r���	uX���'�S)�r�Hb G	6.�}Ux
e��Hn�G1��?/�km}��ܚ�������     n�r*����qfMo�6�A�/�&��r��3 E_�ZNT�3h=Qv���܆b���Qԃ�$�� [39zl��Po��(����  ��.b��jItN7Twy���Y�,���C�Fbg�SR��AҍԌ�p�%PY���}#%D_�94f+�$�.���9��O�h             n��淴�2q��٪��޻�X���JttԻL˽u�j�  "*�&�%j�Z��~��%���2�j7P��������A�=�>%2�����C1|A��i���;�׾/�~�n����   ����v��JȖdT�̋Nnxc��f)zH�9HFj�xjh�m�]��^Չ�@"&��PMZ���V�dG&�"X����    ��RZ�Q7j�Y��]ȗE�C��Je8��G���C���S.�9W���`@�����I���;Pr�uE��R����vt��C5,�� ���KĆ�.4���F�jz�˨�7Tf!�7!�7P�C�9B�:
e��Qx��0��B𜌞�M���N7P��.�?��߀ ̵����AL��r�b��L��ɉ n��7P��py)*�+����ɣ1ܢ7e��s�֓.�dM!���J� ���s�Q"��LfqpdH2�$j�6@�$qL��# @`��u*��@e�!�� �@5���}[��h� m� �                                                @x                       �nZӳ��4�X\v�%����#Q�,h�pNJI�4�m�Cm��4T��Y�P	#�*
��DUZҍ8űn�n�5���$+%Tu���;!&���IeCm�DcQB�[b��l!B��6ں7H�nh���km��D䳦������ָ����'(��)sm�oZ��5V���a��x|*#TL�w�����|���Cm�l             ����-s��m���S�[��B5"6����<��<���ם�<�  ���]f�F�l��{���!t��>��S.�b��"�3��IS)�hF�j:���4?i�kƎ��Q�z�nkދ�.��    $�J� ����Y��rD�5�Q}��ј�V�u!�� ��kI�B&��Qv�Uy���s2b�� �gA�o;����>}�����ϟ�_�  �
DV	��7,�Y��;5���̚�]�)�QM1��1|v �~'$y	�\4���0�y�q�ŗX���`���$�!ʋ��S�|Do!��<����  t�i�J��&]��3f!�7!�;�wN7P���u�)��n��Ի0�ݮ�M&�;�|@�A]@ח�'#�w��]r�����w�d��� �!"�a��D�K2 ����Z��唓�����Fbd_�L#1��~܅�^��t"i��z���`���[����Ǆw��� h              %�nn���puFV�����Kz�[���v "[�  0-�k��r���Ms�/���A}�%4�w+03U�J���S,P�(n��A���䁺�ʍ�= �/'�)&�d�%�Uk���s��    �,��%���%��"�FW�L�Á,��&��:��ַ!�7u��C�!v����]�>9�F`C�k�Si�� ���Q��gϟ� ӵu7jgjt����h�Ó��*7P��p�)P�QX�� L��7TW�raLv���.�:��I�B>�cuFcc�;�  :s9��9
l� �B�t�+�v
e���f^��䂘kޮ�NV�~��W��&::��99=�������_�  �[۶G2�LK��f�}���&��wf*�����us�Y>s��3�u;�~����S/����K�m�3Z����$                �TK�����[f��]UQ�V�:��Nٽ�)����γO7� II)����)��]�,��`)��oك���|��zg�YT�\��7�]���Y�3U���|�� ��ifs���e��e��<ކw@�u�1K��2�����ނ�~�~��x��4�=S_~���}��  뉲M2$�bS��\��*�r�d�˵}��Gy���gs~c��C��$��}�5T��!E"�I!�!%�BP�	R^����=����ѱ�I�Ȝ��<�S�(`��@b��Y��'�v�w�w�o~�ʿx�d�����    j��r�-2�L������ւ�{�}Y�=ۥZl�ϯ�|>NI�S��* � oB���""�rWÜ�]����w����˯�  ��Kǧ��=��َ�z�e�̻����.U�fuY�N�Y�yw����^�n�΄#�o~��'��}��             nKz�3Nz�:7V��V�u�v�bI��W�崵wz��x_  3V�d���m��Ϟ�����ԪktvK���KۛcVb�xjh����;��I�7�}ٍb>>w333   k��ڐ�;��E,����,���S+/��h���{�6��ͭڳ}J��9̻�����U�R�r���  r�.�-r�j�%�7�m�p��ۿ��n��֓/f����7y����&���O�9{��NS���ϻߟ��_� V��C�L�3 �^���z�h-����ul����Jrw\拤���%/�k��D^���-U�����c�>���<�   ����ܕ5�o�>���o���&��<׹��i)��V]�mX)�������`-��������JfffR@             n��ٵj�m.N�����&ٵ�.s&����Rs�z�c�  I	kB�ܧ��7>]�����s��G~_J����ي~�-2���׋�u��v+u|=�����z�� �k��r��S+2���3���S/y�sA�d��e}j��9�+��{?|S��";�]�����e$��ZI����g�    �9%NQ���X�/3/&��]��Ȭ˶����ݫ�$l@s�W4Jefo������'+���p����    B�p*�(݀��t�sٛ�o�Y;�w}� �������[7��������]���
��n��g��W*o|�翿��  :&q���-ː���ͫ=���W۳y�>���L�]�~���[{�Kw�����✚�r��7��9����dƇgffffa���hR��@S�����*(,v��=P�&�lS�M:~��,�2;� *��`�\�j� ��
VD�FԊf+�	�� ���� !HHD�=���T��	Q��� �vH&�$"� �`�
  ���@@P���qA�t��S�b��Z��8B��������ce#����j�P�cdPt�2}��(TTR@H@�#%D���uO,�%Q;[ؕ����R���湅���Ǽ��q�0���/f��O?M�}������+���*B3�����,���1����Cl$^ҁ���xy�D'm�$e���%`�S㞪����2��0�fy�jG��@$\�U� �(a�(O�������O�r5��:E�]+~����[��}V�XO�rB[�̿����zm"��a��! Cb�W�"��Dqo���_!��s�ҴXS~ƤB���h�R�3���5�U�ō#��1w�/g�qֿ�;D�S��Q[��J��MN�6����}ۢ�qf}Q�$�I��#k��TPo���C虎������ȋ!�# ȬI0RD� B!��Pc �Y
T�VB}�II		�$TF�a	$Q�@�$�I@X�E$F$T�XDH����F�V1V@XHE1�� �1FEBQ$C�CdI$VA�F@D�Q�E��I I ������H
,��B�", � (�`����B����*
� �F
����, �B
� �����
��"�* Ȣ,�"�", *� ���D$D`H"��3l��VW��S(EȒ:������&p���=���.��! �RqVAa � �P�1�2 � �����0
�-�h[Ʌ�X��U���A�<��+��+L��L��r���h#h�� <n)�[������6��~0l�z���f�$�I��E��i�4EJ�;_�_R��#�
����F�)���D��Zɐ�	q瘍�����6�����֛�����L^V Ϩ/:ڡwc(��&���r�SS7 H���T0��|V�}�Rf�k%Q��V1���g��~zC\���ʂ**�?4B@$�����$�v�x�#vp4��+�`	�Z�=�(��I�N�!wP������3Dc��PYw8X��O3PHHC��&1���1^M?	��TB'N��I"HxRe�ʅD�(�S�b���r7�5��C&F���fW�>��\������HH��t�џ)>]Q�W��"Yd�5�H�yi� ��F,�t��H�vt3e��+v�?��uO�6���A�y�)�1=H7�A�G�`�t�KL��[�8�`���)���Y=1�!����_�~ަ��(	!��,)�3�C�d��_��pt���X9��h$8�t��P<�a�?73/L��>Mʠ�rL	������`d���~)ν�'	:u�D�h7�㉨�ҞL�V2�˦sJ�z�AAu�h1E���͆�c��y�qS���M����{�:��p�/A+����&�I���29��25l�]��&�c&V�sf�Z�Mp�EAXA���W;���zM�!���H�&A�����Jَ�n@�n��S�3��Y�4А�H�6�Z���	�@N#�<+��ƭҤ�+e��Iz9���p�؟PƱ�Raw��q/�m3�w$S�	�Ը