BZh91AY&SY��wc �߀py��g������`�=��Ls�     � �.*�����hI �MOI�<(�M���h4�@%)$2a a&��  8ɓ&# &L �# C �H�*dS��    �H��~����'��2���4=�h�@h��A&ʞ��j<�覙�4  ɠ�Ղ �RW��r���E]D �2�g�K2D$d_j
0*����?s`@�X����(�2)8p�˗ ߎ�6����N�������]����~7���<x�Ӻ�û���}��#��q���;wwv�}����Ǐ:t�#N���_Os��8�$8���t�w\iӧwv7ww����Ǐ#��x���$"<����ﺾ�qP#ӎބQ�]�e)�����Y�]��U�\D�E觱�o�gm�eƭrb�ӎX���c�bR��` �d��(\0lsvJ�N�I�2N���J�6ӧ�7/U>���&.���V�3I���9�,�@�����[��ssv�ܦir��Җۍ��aT˺hݻ�w3��&����{G���l��P���A�2i���
��_8S���3��t���)������&8����#�\�J�6��Z4]���̓����ե��IQY�שՒ M6�[� �061E4y�Q��q��i�x�P�f�Y�u�j����ffff��iѻ��[�����wwww/3R2U�1�� ��*%e�i^؁:���6�4Y8�(��ź
���@ө5��$�ܝ�t<tEP�n���նU��2	��B������$bsv(���_-�3sm4�?h\�'2P]���	{�@|�U���+��YS�� 55J�83D�$ϡn4M�]���؇�9qb&�s�C��}��%Is�Ј2� [0 �`L=��fh7�Yΰܪ�f���d$��[�oO�,�{���E�.uß�x��@�ӧ2X(�J�4Ir[���c��&�
wi�����dDI�+��e��c��zu�J@#�L����Y���2r�6Y��'�y�N`����bp�j-����߾%;��#1+�$C��	g�QP^B�X�B�O�'���j��������M����C8.p�r@Qa�f!�Z��,�E0��e	#��q$x��;ϓ��~O�J�� �8ޝ�"�c\Dqo��n,K�a��D��� $�>�!@�5����(bX�B-����vؼ,�2@�=�]#�Sr,dȝdd�>�qw�W;�#�Ns~�	B���#y>�$�~��26�;���3b��duP�i�Hz�k���bt??�,4�r�_�h'R)���k7�1"��%�32.�$�Lߖ�v�WA%�C����AA!�4�V4�kƂ�$ﻓ�h���`[�;��Us����K��� �,�� Y%�@�+��"!�f-B������s�9��͹xB�Gj`t1�#>���ޚ�LD��M.h�6��Q�?=½{�e�~�x��#�zӰ�w��������|�/e� ��{p��s|�Dz�O�����O�Z-��6����  �ܐu�'7�$=�U��8/��AP��|�E�<�8#�Ͻܮ��Bk���^F���Q�me� �3����f9��p�sb��N-;�:�Ճ�C�o{�r��l��0vf}��3��
D�}��Z��L�m�0�k4��=B��A�sP���8�gJ��tŜ�bߟ�`���ⱻ����G=j�\�J�w��d��υ2��n��aL��L��	�W<�\O�0H"�JЂfH)�Wų�>5��R������O�r|��R񃞨�?�����0�ȟ��$�f���{����+~z�e�J&=�Kan*<n8Y6D*2	�>��]�1�z�3o(sýX��=�3b(�ӥ�=+յ/
j�� �!�y3�����"���7���@_?^��[o�f2_N��p!�fE!^���0?���<-���/���˝�r|燀�E���Ub"!aE8ǳ���t�$+�&�oM�w���#���3��a���E\�QU��y�q����k�-B�E�+!XJ�M��3N��b�(��%� ꐪ�9d��1���s̒�SL^R��V��$�0��2�I�MJc'H��l��d�Y��\�ї$h�4ETa(�*�i
�d�9�p�ta�A�:êl"� ,�,��U��#�l�椼�'����ȁ����z��OB�g�7bX"b<�q��O�A�����P9��u)ݎ~W�]����!BsLQ�?�m�ɗ�?�pu�j��?� H�A�t��{��w�F��Hd,��	u�UR�qn�4*Z��jt'N�z�{����'_�d��Fz�$��O|G��g^BY�!j	\Nr�sn�u͛�k�ĤgV
�`UO!�q�8V˹�]�Z���<�<a�A�Z1E��E�PV,X���)"��X����E�dY�1�b���@.�4���.���=ߔ�<���c���G*��00��Y�,"��� �����f1ߵ��q6����.�G[�I�\%����a��'RV�w�t���s���(ɴ�_(�iH�P髩?g��6�(��&&�j�㟈�I��=$bcݑ1��F��n3��k;˨z� �P���o��[�y�1��7o$�5��(	�
?gk�	�`|�;a��A�4 �ژ����j���+agI,l����M���Cpwpϼ.V��i���)�h��4����!�cE�Syd�b�X����gI�Z/!fu��{�P�o�(􉧔����Pe �����r��gD� �veJQ��)F��;�c`ͅ1#��q{ceÄ�E5"y_�s���|oUKϯs�1���tМD�<K�N���!z<��X�E6��S*����K���Z�ez�
�$Ty�D�$�k�B��t�ƳOt�*��ku��	mR���l���`AX(��$���M�H���,̂��Hum�D��x9���b#�U9�iq8J��0�M������D%�.��8~����מ��A�m�s���H�
8��`