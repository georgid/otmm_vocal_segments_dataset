BZh91AY&SY�� !%_�Px���������`}X� C��� {`�$UR�T   ��  u@<d�!P�T�J*h��T��hh h���  O i�4 d2hi�@`&�M ��Ъ��Кbh C#C@ 	5�*�������  "Q#M&50L���&��='���Si%&�O�?Td��)�OQ�F����~� 
�@�S!]B"�A��e�,�I"��PQ`R�ԒJ�X͂8��B�
�A���i.��n����ة�]B���Vq�d����&J-)h�]"�IH���E�"��D��g&e�̼���t]�IH��j������Z��əu�&e�e�"RPj��轅�R%%H��t�KJJ���J�k��Xj�������)��ґDJD"%"E�"Rd����2�-���\Z������-��f�f�My[�uA�Ls��W��1|55gU�%��;�谮�T��DI��¬a�y1y�r�!̑Bi�5p��Y�v�ЇV���FZU�VZB�[�؃7f�U�n����	Z`Ȅ��Q���{��T���P��UE�M^p 5�y������T#j@���#6�5�"��͇1u�z�x�e��Œ4�-����nQ5����]�[UN�"��nv�w���vQ@ꈛ��D7�*ьu	E@� �Ӄm�1�$���r��nM�u#%B�A6�,�%��!I��0��o%�������`"�b��ݩ��h��	4m�``0!~k�1�(�b,)�~<�b�'{>���a�U,�h�f9j�+(QX&;c�m��\u��
�̑"))IH0�N�J���DМmD�y[��+jۑYI-KI��ӷ�����H�5v��q�N��n��ٳ\��(�	ݟ�p~����� �>��7�;��r�۬ƛ�n�owm��w�����Û{�x�ffc����<Y������˼�ѭ��{�7wwwq�����u�����u��m����m�m�ݶ�m������c�a��m��y{�Vl�a1z�%W#aQ��1X�����8�bԬҀ�Y,姰r]�:mکB�ٸ	2k*�V6fDX����-�CA��R<I�˓fV�}���zu��ă	��0wk�,\ŝ��)���_�p��:�`
[�T ��@k��w������9G��w��&`H����DL��+�d�"$ę�%ܻ��9ڪ��m͒C�պ�,��v�r&�Fd-5���&�	Fz`en���pz`v�5������L��;vhb�@p)V;1��؍47x�>v̷��\����M��9���ȉ���֟`�=i�{ۨ��͐�e���t��=��S�7���EuE�a0�E�������ј�]H�\��בS��@���[�pyw;�� z�����6�v��P�pd�Q3��Jg��s�O,<�%��׽ꪯn�ggmQZ���ǎ�Fez�:�L!�f<;�5��"�{o����!�!v�@�a��Q�Nu1Cf�j��,����L�;��X�vw��z��I�����֪��;�>�+��f�vQ�'}�3'�3���]��=!�09�;����zx�0;�P��:A4p�C�>���#����3]�7�7��s�=3i4�pÚ�b�H_=oYǉ���(m�M�g�ܴ�f���q��4
&�<0-��tJ`z�#�@;Zg��'�H�s+� �;���<I�[ʝ&2t��I߽
��<y�����i�9�s�!�l-�	���hr�2�T�����WUUu��]�L��Vm7��UT��d,4���v'2󌮹���VQ��ewePt��� v�I�e��<rm���w6i�7�;g��.냿#O �|��S9*��Ɛ��wP���saۦj�f��<�Z�{��������mm!g%��Q�XE���z�'��G8 ��Q�⼅���Ϝ�&����C��:5
�1�s��S�ꠠl{�:� �7���>�:d�|��6���y8b&�H|�><�CR�Y�He���Z8�z�c��l�j�Hs�CI�Q,�k�0�!�3���54�F ����WO���.���M������yJ�����)�yg�!�nv�ٝ���n�bwz�s5G	'ރ�v1�>d'�{��wDq ��r� ��hm{$ޗ�	s��z�D�xj�,�����$WP
}s�ȥ~������D8��z����=ڸ�C��z�nK��&���]��������ܮ�� �(P*,aT;U. y�Jha�_u,�ڹV["N�&�g$�%�W�+�P	�j!˘3�(�kg`az�:F��(s��1.�-+�Y^�Y�/UȸP`=T�n�C<�p�(r hJd�reD�̩�
���Z���N�Ǒ+3<��3��<�53j����'d�r�קT�f�c2e�� Z��{$Ҫ21\T��L�ܧ�8,?\���F�t-��Vp	ݙ�9�̊�T@��EW.B�"�c����M����
}��X�x=�����Gv��p.J�����vf��=��/ֺ�6�LY�w�o�|�w���^J��Ֆ����"y߭�\�ۈ{�X��gOTk����p>q�����*�����ȩyjdH�bЀh���gEZt�]�W��u����t(���͎#�Ó�9P"�����I�ا�};[�Uwq�^�)�O-�[H�EL ����������<z-�<��v��GK����IT6��zio�у�)>���X̫�af�������3^P4�gL�r�6#<i������/�0�Q�܉�#>���;��j~3k��B3��b���5�R"��� �/ޱMR�ƚ����Q��+�[��ճ�8�EUm�z��2��( ��%�DM��a�Tw�1^�RN�Y�s3���i�U 8
����o{��tթ#����(�ˈ�W��άÞ�<f.l3Q�Ew�u��C4U�#��{�N���C��rƺ��0�Ȯw��߲N�wƐ��������(A�GO�@�GǵO{&�ކ����ɸ�T��ٮoН����:((�w�NB�������`�y����32����t �J!�k�3ٷ8��Υ9��i^�L�:CR�3���;xw��}}-J����@��d�m���h�m��z�޳����ႸH��	9�%�=6D�$!ArA7#��r,)��2\q�C��Ӗ����w�ӇD^�o��͚Y;"n��Ύ��M�kWx88�n2c޾�涎L��[���r���i�j�Dq@%%E��<+�SZkV�x�&]SX]�@1"
(�~C�ߟ�mL��ws1=�	pTX��`�Zs�@��%F��MǹY��и�_pC�5���+	�&��S�{my�/zFE}*b�G=�r= ܙ�
k�%�r�_0��3�٬���9�SU��|�*�ws�1mF�1>��W���������������|�5������dJ�y<�ߕYl۱(@>�*�/��ü2ħ9|�/ng��U]�κ�����0�ML�S%4Fx�ţ�nw�j&l�ة��W{�a^��^� ^�M�b
����xS�N�Hv��Q=>�vU��D�'�p��~����力�G���#���9�s�;)��"TL\|���l1�'�x��N�����: ���iD^	8�Ž�!J�oÞ��|�{���b�Q��UUVFB"С�8���>���.
���|Z�0�n`<����5-�6l�&HR a�F�
@!_�R�Q��� �PR((n�M%�"�$��1EX�*��"�`�(,��#X��*��X�7EDQ"1�DEQ��Db1�����#U
��DDb"(��J��-,�	H�B� *���R�,�,@��m� �B�%��*��	�a�A�`IXQB(Ф�D%�X��C�m��F�5�/� �.��H�� �!"���+Bn�ӻ<z�ݧM���쯪�����c�)�w���f7'�3���k�Қ3��*^�3���̆�g��)��SOJz*� �꞉}y���G���x�� -ʨ������r=2���j�jG�#Ah���c �{�b��r����AEŜv��ӂx�Zz|p���#S
dȘ(�z":��w�q�Q,b�V�IyY�����W�=\z!q�Xխ� �y����V5����Ϗ�4��-!b1`�$H�)H�H���D��DH�DH���"0F#�V �$Db�Q0QDDADE��b�F1X"#E����b���`��
)	-��0�)�a���LC"�B�_mC ����!���3� \\
�Z����"���"����2(�*2��"����1�g�{���r6r�e$���Q�d_�y�JQoу�E��Q:SU,��Z5�W~i���5d�ax5���e�C�Q��9]�%�ᇞRI��N����.�ׄ�؂��(��(4��F|��[io|wmH3(f�DR�_�s��tN������`��sCG��;`��,�#��T��p����*+P<0��<\t�Vっ�aV�hD}m�\��!�&�s�r�i�ю�wMC�\��C���r�נt����K��yL��Xӿ�?��<��'�*BG�B`G����K����g�j������v���e�(��D�H�:�j
.��� .��x�ٟ=����jQaкm�2.<\XP�
�U��0�s���M��o�&<�{���mL�`.��,��w�4쒔�)G����
	R�T�v�k,��� /��{eR��(�)��y���!�p@^�
�8�zfDx �w��d /-SR*5vm����sH�9�8����zy�!���Ql ���n��ܑN$:�� 