BZh91AY&SYG�B��_�pp���f� ����at�    � � � �� ��IB�T��#�    Q@�P �A�@                 P  Ѡ                 �   ��J���g|�����WN�uQ�.�St�n��ס������f�gӧ���F�e�  ��J�*!T"��5�Ы8�\�T�ٳ��*�m�'m��R��4�qʻ�Y�Rm��r�+JhU
�4���mJQ���4PUv� �R�T��S�Jt}p��XN0��w�R��j�WI�Εӻu���X��wi��T���U�&�F�ykg�Ӟ ��D�*�.;�Op�<�.oj�u��v��tdOm�T��:��w:��yj�z�U��{{�Yw�{���p9��s9p�[exZ�o]=���O83M�U�g=�^�/F�]me���Vj�Q�t�v�Um��  ��EP�� �z��аs4u)���6�j�/[ѣc��G/V�m�x��[V�u�g��&�݈;< `�J(�Z��^4��s)ѥ1�Y�����<v��.�K��3{ݻ�Iۖj�.[�m�X�X�� ��D���ތ�W.�jZGWt��v�����K���ui��Wm^�]�:�մ�Ǖr�[o �QH�&^���T��W�gj㪳wC�k��U�
���P�f�&n�-�:����Ү�ux ��T�PT�s�j�<r9v�V�&��eWF^Ǹҹw����/v��
�t��]�]���s����NU< P       "���L�)R� ɠ    O�J�M d  h  ��U)CP�0i�`&��2hD�*���H      ��FRT���1�D�@�L �!R���S�̣hi�#	�mO���UDQM�����z��?�_��݇��}�^�r�*��Ѽ�5QUWh�*�x(�����TUWH������QUX��(��� U{�����jEy������iQ5 ��S��T�8?�QO���D�OeG����{
��{�$�OdT�AOd��*��>��*���@}��U=�ȧ�
{ '��{ ���u"� � �"{ �aT�Oa�EOd�DOdT� `T�OeNB!�(>�)좞�)�U=��A=��=�C�'��{�� �
'$�UdA�PaT�� ���ȩ쪜�S�=��P}�S�P9�(��{'� �eT�PdT�Od�:��E=�G�7 ����'���"'�!�u�'��n�d=��C�N{�{!�'����a=��^G����'����Oa=��I쇰��{	�d=��S�e�����{	�e=��S�d9�!짰�	�Od=��� :�SR*{(���{(���{"���{���{���{��*{���{ '�"{��
{ ���{ ��"{"'��{*���{ ��
{ ��
{ ��
{�
{(���{ ���{*���{ ���{
'�&@!슞©�
���"��)쪞@��"��)죨U�Oe�QOe�EOeT�QOdD� Od�OdH�λ?�p��x6��[��@wHU(�;D��x\á�������/pJLL������m���(J��}]�1�DjB�:�pHw	���)��!BrR��(|����Dfm�<��^b�s.M7,��3�����'�ˤ3_w��od��ɪ2q=5mf@nRj��MH\��[�)�&�)JB��7!JR�Hd&JrB��MHP�]�|������+y$��Yk�]�e.X=�t�S�w����FBR�&N��4|3���>�uA�i��^4�=��={��%	JR'�y���ݖ�1�#"�:�ف�[�:#58h��捇1���\��d`8fb&��Z��(J��4m��Ƿg|��(M�ozÎ����ޣ���<H�p7�
��a����:5v�JR�sI�!����xh�ȓ#����:�~�ٮ���dpa9K�R�8	�Dpx�#�z�{�w��ޞ��^�Q���RDd��N1g�\�w�;��<p�b��G��kXD�7�߇��Z޸�z�v牎�0ٮ�$9	�NBPk}v�dF��wȬwA�14I)�GK�F��u���DR�;��熡(NJd��1�G]�Mu�~o��.�{ff�p��ozke1��
��(L��:�����f7Y�xh4�;��JR���<A�G��� �OM�B#�,8���M1�)J~u�HQ��N�DA5�bm��%	BP��}�k}y�w��誜H�aBR��	Hk=l� 9�E��Aq�r&p�I��9߬s�v�fb�ލ-����p���(�4Tf�m��f�8o|20�F��!Bn��a�n 슠Ħ�4�Dw��t�㠢5�D�Ѹ�OQ�d%bn:�%	�L��2p���)JB�w۲/zX���4��k|�A�X3A��L�������=� �H��c���>����z`h5 x�8�
\��K��u�12��C���ԐntTu�4��ƺ�a�C:�'7��=�ι��9.��j)���#a�uG������o4�C��o����#���²v"�tWlLu���ml�O����fL�ƴ��\�G�c�˃���y���s�����Y�txt%��:q�ٙ��<��K�J��(J|����,�l'XbY��F���;r�ֳhd%	BR��'�k]c��w�բ��^�&T�d�MD����i�\�IFm�l��F��[�[��1̍�Kd\��fp�G��d�2LL���0:�%)HR��:x�qr=`ѩǮ����}:�^��\�{�ѩ{rt��G��Ըw���Y��E��g�y%�G=<C����;��wr���]�^��\{i��Մ�����a�����)�;WO���2
A����|�;��Ƶ�)HP�!BR��s��{�M��Y�}h�~.�)JS���J��J�GY�Q��;�v�f���5��I�V:vӄ�	����r%)w�9�/%:�EU�0u�f�(��GV�A��NZ���q�NO\[Z�Fa�2����\�ǁ���V�V�|��+��wD��!)O!(�p�s�&5���`d�k 3:ѕ�7	Bu	�Hy���sg}�9��;;癇~z�!�6K�I���t�7��4�����y��:�;��C-���[v�`ՑVs���8�b�Rr��`i��[7�,���Z"#4����y)HP��P���'d=sܟ]�ON������}�X�yg�{�Xc�&��HP�F�a}N��&��f���R������\�NN�@��y� |�P��;�lul�<���b��,zyĩ�d[��ĵ��G7s^u.�=��)JC�:0���L�]G����7��Ӄ��W�R�K5�%G��}���%��a� �=S�I�P�G�@:B �t�Hb�%�"��B��zq��i-Z�F�c��bL'3�ăEI9!�!��1+^�;�x(�u] ���\������TB�Bm�����A�;~��� ˯u��t��h�Q����1:�ԅ	�!Ԟ50�2`���*��M�9"4'r�J��)
�	��g�LN�� xőVE��������28!�oh��<�5㽦�$0�ty�g7�qX<D:���_$�f���������pѾ�N�Q�N�6�XbU ��\ͩ�$1j,B �*G�׋�:�*.Z���\$��E&�7�=uh��w�c������y��h�$)��,'1�U�s���F�٧$���t��5!������e��uk7���Gfr8���@��rtE_m��D����$eg[��<��`tjp�ZH!0��)���_�;�>Q�p'�30U�y<����朔m]}�~���,uv�]�s�{��W�pT�O�����#��NBjM&��C"9�vz���쫝���[h9Ht�]tQua68x�������`e�T<��w�Ґ�)JB��)��,���X1ǌeh4FK5�ڔ�2CYa��!k322,c�+����ܻ��qٝˣX����Y4��#�F3f9�P������!`Y/A��`��d�����j,�C�jB��)
��+��3*�jB���d����J����f�7��<mX�BRr���Y��0��<���!�7�`�����U���:̵˜�8���7.����N���h�5.5o]�A����nu=��a�u��槃���.�1��"�#'��05d�D5C{	`��2��VJ
`!�*��8��S7!���	R勳7�Z��'PkJPdɩJrc�2�#�2N�1�*���Q��6Y�d�Ŋӑ�u�s�f�ћ^��A��zcy�a-��d\ݮ��o�Dawb�FA��Ԇe�h`bfe>Fjj�Nl��6t�u	�h��'G3~s;y���ӡh<%����٘d�gI>c�^����p뼐�:�Z1���Қ3��x�)HV��9���@f�&�Pt�BV��j4Z:��޳�lҰPTF��=V�=p*}�Z;*wQ�8��Dk��V!��7�j5%��3n�x��&�pUgT� ���]��x*�e�޺�f�,�M��;�Z�,�jz�1>�Ɍ��kfV<�F�6�@h�p=��3!ѨN�����0e�e�d�9.FX�Y&Dd�5��[��dRd�C����Se���W��.�HQDh���-	�'%)�7k��w:.[�bf<)���:h�ᑐA;�+X��$���"3:�ܧ���Om�dj^��xq���30P�gzU���gT��{�`���@d��c)2�����Q��r��i
��y�<�$ζak|:���#%�N����CD �cˏ�� 9�u�D2�^��וIAD�@�cǮ�њ��8�s�բ՚�삎�9������d����#0�Eը)����N@�l�Q�33����g��Ez��醣S�9�r�9η:�5��WV�[5̧����Q�.�Ј�7 =��,X8�c�۝�~(�q��'�R<|�er�
�%:૪6
wrا�6%*��ѫ.;�y�Xc8np���XZH::4�θYF`���=uʃ�@�*�B߬ ��Z��z��d0��y���Akf��d8wY��{���+]���a�s5a{di�:}#�,��I�%��gSY��((;�M.��uf�Fsq�U�����M�4��OY��5;�i¦,����"r3�77�R�L���6�p2q6nN�BntGO7�:���n���΄�(J�,!���y�<�������F�!�s�u��r��$�ˇ6>^O|�Oh���r"l�$�&BR�3h��%R%)HP�������R�9i5)Nd�i�!Hk0ș�
MA����'Ώ-��lد�BP0������姄�W�a�Ju9��C1�a��<d���\5V=l*�Xl�t/���>��{�nk�v��ݮ{��Jt�K�' �24C�!I��`oU�P`FK���n�rp�f�5k`j�F�D��6%8�:�f�8�V�,�af�bh,��NN�oTZ�����VG/4u���VXQ�kXyi���a�w{!Bjbz盷sۣ�C��)�����q��,��5���R���rОL"@�),#���'
594f&�x9:7��110�k�<�C���j�G]t5!ב�����z���;�r��ǎ��X%h ���Q��G	��)�)�hWB�`.#�bp;�<A�s������ˍɟ{��ǝ�=���c�*���h�B�٬ydZ͆���U���k^0��yݭ��]�&@O������߶�{�D��oI����A$�����I�����)��Ж��q��]�����G�A+l��0����<���fj�=y�vcՙ���ɾ+�Ӎ��~�'LU��w��=pn�����n�+��l�����jb�P�#��O��K�+�?�?������0
����G��?���Y�`�(̀��tx?�ɸcd�}��U�
`�w@ǯ��2i���K�Ʌ��E�����a-I"��������Ǖ��}�w�,���$G��uZ�f�������\Zu�K�-��E��N��V;vڨ�OWS����L��,(�`G=���b�5�כ�`��~]����`�6����K�b����H���qd�����N:P<���  �C���s�%�վD���ѡDj˯;��jI�k	Fdof����A����Ӻ){��`����ofC��������|���)�=ݢpA�;�%6�I"��bC�w���V��똟w��l�@��䶉*s��ky�o �:��5x���[H��GC���t:pˠCĀ����(�M��G|wfrc�k�\���)U�` y�Y٫|A�C�s�Q�G�+%"��$DO%�*.��Q�,�p^\�+�r�x�P=v��4֧�jꑺ�E�q*� +�;ϔjHa�$�� I�<�S�آ��j�C���t:t:� �C���t:�d��$����C���t?����t?����t:�C��輭t:�C���t:�C���t:�C���w���t:�C��-�I-�@�t:�C���t:�C���w0:�C��r�C���t:-��C�[D��-�@�t:�C��&��4H�E��C��$�4H��(�Kh�Kh�:�C�����t:�C���t:�l9�	�[D�[D���t:<dP$�C���t:�hv	���-�H�C���t:���C��ΗA���C���t:�C���t:�ht:�C���t:�C���`c%U-��LA��t:��/���|�C���t:�w]�C���t:�C���t:�C��� (�:�C�ѽ�2C���t:�N�$$���:g(t:�mImC���ܐ� p:�C���t:��$��$�C�F�Fղ����t:�C���C��2�uTZ�C���t:�C�Q��e�}�:�C���t=ݡ��t:�t:�C���t:�C�[D�[D���t:�C���wQ�춉$�����C�ۺ�K1$����t:�C���t:�t�%C���x#D�C���t:�C���t:�@�:%�C���t:�C���vKh�;�6��6��l�� t:�C���t:�C���w�~� ��:.��h[L���9C�۪�E���t:�C���t:�C��-�@�\$�Z;���i�� �;���8��t:�C���B����C�I`t:�h�:5�t:$��R�4:�t:�QyC���.��C!�@�bI��	q�z�����(o�\�w!X�<�*')��¸��'�kQht:+ �J�C��o�:�����|�o��W%0f�!�@� t:lɼ��[�:��Á�I �m�Ic�#��T6�V�-ݜ��v�J4���	�q%�칽l`��  t ��^��	�n���C���vKh�;%�H 5����uH������a%��&��'ͅ���	U���kw�ͅG��������<�l�q����
q��YM�hwޠ�s�U��'��w��5�5�0�C�p�Q�w@lJ�����S���~ѩ�A��jj�� ��bM( -\�`C2!��[�K'h��(Y��I�BT��%PHH�C��wP�I$�����=�qSL�΅E���t:�C���C�� ���(L�`�FM>0�aA����T�}�l�J�^�D���tk��t:5�$�Psw�V���y��9��I/74�[�D�3�
�V��a��{����C��o�`.ݾ>�zw'�bR-kΛᧁ&{��0V��DZq�v㫍{xV���NIT����HT8��o�nZ$�^��q�$�թ,�N*�n�^G��s�3J�P)`�%�G���ʸ�m��I�ww.گ�MS���o�h  ��k���t:� ���TZ�"��m��C6�m��n���n���(l:��r�rj�I����#՜�cz�)9Qh��;[h&�C���N�F��C��怍g�͹ĺ�HEu~�7|�Y }휈���i�$�C���m�m�C���t:I$�C��� P�t:�C���t:K|�Fl0�Aa��t:�C�wdJ
�pz��}M�-&��(�J�0�y�nhH��Ba��s7���=�:�]6$����06:��O��[�q!Z�d�HR�/#�������v۶����	��rtʴ����Fb?��Oz�����i�ّk���װ��i�$�*7^�]GD�mnH��s�ZJ�o^�'ۑTM��6�黾^Q��O]�}X��3/mK�ˬ�x`+2�7S#� ��l(*���;�xyI"-h��	�{8ý�$HFՀ0��˂�黳���.�$N�?9��c�3��C���s�ѝUh�u�k{����Bꓹ'ǒ���.�&�~��*k���Es��	���}M���=�4�=1-��$�(��q,������b�y?q��k0>Vjz���[�����
�p�v�[��$�}9�]仺� �)�H6%���[ +�&���L�,J���K[���IF���lHWD�	��m�It'0Sqq7׸�����v�Hs1$賻D݉��67��I}�̣�+_2󲀣o%G0@6�"�^��{R�-�1@��A0gLl�f������Mz󳆝{30�-�3���3Z���C�J6�tى���پ�-��x�z�2?%�l׃_0?/,*�^�z��un%,g.�xl�8��W�6��ei$�[�2���}+���F�&k]�}��!ٮx���=���I$�����m����Ö�Ј� ��l8/+]�3���vw�ܝ�j��IG�^����v�z���G�T��;�=���g�}�Fb�۩,���Mݩ�ݙ�F-D��Bn�w�vwV�r[Gz?A-�"gp����+čѤ��]Vz��Pe�9|���z>t�3&�q[d��C���t:�aa�[4I �A���I$\�m�q� G
 ��Ȑ� ���+����o,�]۞���3A�@d�J�t͑J�H�	{�Y�5����(No˪N$�2r 2�3;E�O���A�E3�j�UI �+�qo��D���RK�	� ,$n��T� ��w9�h��P��S�v&���3�]Ԓ\��=��<�+-�}��O��7$��� l877r���Z�g��u+�jH  �8�\�����TZI#�X�H�C���t:vK˸�-�C���t:�+����{��b�wwA!������G~W �
�Vۙ��� �ݺ=�d̰Á�]�KA�3��ɐ����p#����Ğo���u��71a������{�F+i{���m9�y�%��t��Ĩ�'1 i'��3w,F�4n;�J{A;�ߴ��y(���:W{��K����Zs���|{����R�K��X��Y@����h�p���y�f�ٺl̷=&R������o����v���H浀���#���o�	jI���_��W�z��}4��3��Я��}��  h���������=���gś��ڮ�2�"}����[�S���'�����>�G��$��fs��Cb�^���ۄ��� 9�C;`(iwx�f��J�Yx��s� ���Hq}b�gj f��>[���R��=��h`����r����x���5�2B�5A�Ks{I�4�=W��Ff�����[�ty����M+@�w�D�:1�T�ľ��b��@�a�3Q��K�:DZ���P�q��=$iP��2��&̹��ssu����*��}�ؠl੔��蓸��,H ;vZx�8 ���x�y�ϸ%�y��l�,,i�������)�a���G`��+|����j�0N�ww �;E��y4Kwm�"u��t:Ԓ��! ��j��b2��J4[4H%�BY��*f�Uz�����N�,�Ju>�����k�#��3L��X��0�z�[e�w}5��}��<k��2�$���[��ZI���I!�,��������sn�[z��o�h���#�>o����x��.��/i���h�l$����B�Ɇ}���'@��8�`�[��0g�Gܞ9`�8���s�H�*8R�Ss����"�����\�G���4'::�f��q#��#�ޗ�	=Y!J����I� sjE�/d��A�+��M뇉$b�$�H'�U�t�D�C!�@�t�k�NGB!�:w|�۰j��>�����=C��@LU����$p~�Mԕ�dV�Ƀ�IdK��A�M�Vl,:ō�f9�T�!�Kƒ���L���輆�1�����htX��a��t:�EV�$����t:<���	$S�ڗn܎��]�ͻ͏0��`�>|�a����_>)i`Rh���� N����A�����t: @
��丝�$�΅E���$�d0O��L�w�HZ3s]��{�HQvC
�s��w �@
�'��F��
�^��17@R���0�NKoN�E8��L\$�yBm=N�ز�r�C�U���� � �I�t*-�·C�w_)�|�)��/=Ь\������diA��_$�H��6�tn�@� �M���9&���Ӥ
�<��y�*k�F{�ȟ>G��n�b����ܯ��?�|���w��x����%9��i��1��Z|nD��՜伺��j�� t:.]Y�����)6:� y���ݩRF۠$/���� l�j�N�� �]n�ݖŤ���.@��Kڂ�\�f�d
�N�wKpH{���Λ�&�ʳ�g8f,P��7#�I�+uŠh^�sE�բ/}g��+%<������b�۸;�`�}����r3�|��^�zN�����Ik�q���e����n:�G�yJ��cu�p�p�^;�捻���SD5d紃(Z�y��EFC�yG "ogx�̩��wZ���wv�á��Gw�w����#F��X��5Իox+�6�/+<���3���ߏ�햨��bWwu�b�*,�I&�C��5 6�O����X�  8I�t�D�� �G�9qeLU�‒hM���d12J9�x�+eZ �i
��2uFm�$��q�x��C��������[�����T�+�����Á�y	45��4*�C��p��!�A��B+CZl�\�ؠp:�EP�Kh�:�V���U�|��`n��B3�Nn��u.y�ww@l8�B��aѥ��B���b5��GʅG�?����O�|I����]�B���F����;�O���]�B���t^E��*��P$�I&�`d�h}����t:�i�'��bI2��肙� Qԑ�b���w8�<��-,R�p "��X��fHK���S����$�^�n��S���Q�x8�ktOr�O���w���d��ȸ�֥�� ���-&����'=�Hti�q��y��N�Ԕ�@�t>�h�S]0E*BE��<Y4v�[4H&����a�����yI�*�qk�{w�&?�]��,��=�-�|7�e�k�5�^������d��B����=k�V$J�{45GPu�LO�-�>X	��笣��u,̨ʠ�ת�5�%w���f��(1eI� m�.��en���&TP[���C���t:��Þ|�Xo�=�E��$�$�(�0I��t��u'���0�L����w�����_|�v����t:�!�L��u�$5��5��@���Ԩt:jI��I�%����"4�EvH�(-�L�0F�Irx�t'�IXK.	C����ˁ��x�'!��c%�t��.֘�t��e��Ǉ5�.U{ \�q�š?C�Z���h]'(9`�'؂C���"�]�9����D�ҋu$�B��u��k�����zf9�ۚ�� Ġ�$�C���t:�C��K���{j���b�Ɲ$\�?%�sRH_��>|��e��ѻ��C��$���k�U��LI�$�՘��@�t:��"����>ݤQt:v�m�M	$J5$���lfNR:�ǹu��t:���a��r�@�t:�mV��$���������y�.�:�C���u�n�BI$�|u�7vn�v��|�Ux6�x�����sOBnV�A���w�0xj���ZH�{�;Ĉ$�}?r]�J��iq"1(t3׳���A��L���eL�|1��R�b|�`�{k��髉cT:Y������K��mlzN���mjv4�!�X������`7	l�ײ�@�)"��p�p�S|�q�<{�ͧ6���yw����&�DL��64ȠX@�ROw�  $|��6��^G�Q�^�	��C��uN%�m�C��C�����t?��O�|,��t:���kQٜ��C���t:�C��ͷg�>�kR�c�l:��a�� t:w�`>��5�$L�+�-I���W6v��B�e����C�����q,Ē�r��@������t:��E�����_w	{����r�Ɔ�����D�T�����v{��� ��'��_��b�#���ￜ �?EA8!�@����˯��lM~VG��� ���C�"'W��R��C�^�QzP@6`'�� �=TT����B+�m4t�,�UH�$�M M�=��S�@�#"�H H�%aY���U�Dt
v�! ����"�����LK�BL��N�<At"����0QM&�&��J�ڈ����Q7��}#�0:IB�j�P�T1���t+�'I*�^�C����QYO8I0�T�JA,I0�����A5D��D!�T=S�݅A(��b�Q�a�!8+�,9R�A�`8U��*&@e�:PN�|�JJ���	B�g3(&���>�QB�d�dI�$����Q�4L�IJHA#!.	������1a| �	؂� 	�X	e��� �T�(x @��|�O�ZM����/@�maP� 4!�TE�$�XG �M��P�t��� G�Q].���EEU�����?��������O�DUu���҄!BPH��IS ��@�BP�0
�f������j��w�i?���UU]�����z`��`jq�tr�j���,	���ú㌨[�
��BN�Y��Yr�j�Z��
�Au`���5uUS���*-T���^f2pq��kZh:U��;^�I:dq�Ӹʣ�AK*�����,���^�S��kc�4箣�kX����8ӕ�ܻyR�K���k����M���sQ�xxm�	���0�ʛ��:�{�G[�dͫ�NK����@pR��AΞ�a��8����c\���ֺ�eN{��3WZt�,�빂5�ݣۜ#�y�k��,��<�� ��+�7���[��&�L#��ʽ�m�L��غ��{�v狷M��nv|J���ڥ��'\�JD��h.�n��g�~�w�{����¾���b	�!�@����<�@������9��xY�u��͗l�at�9VC����1��g��S�f���Xy;�uɳ�j�Pi�K��ƣ�m�2��Fq��	����ws��9���Ti�(�YA"�����,/H3۷�[�$f�;����V���R��������z.@�/e2o�0��C2�x�N*Tҍ��.��[�ԏoU�jQ�.�{���FSn�H�u#�V$|�R'1��d�ra�m��Fa�,d"Fꪐ����M��hT�A p��Oj�<uI�;sӳ<[p��f���ٙ.�{18.�9=�x2�����<딫�g�c�ա)�%MT��7�=j������]�!�ǲ��������8�J$���R�9��~�9�JH�)���<8h��c2�.����JQ��8�N�7�L4I�Ӄ)��pq,�����nТk:=0܌�7-�i�H��A�L���B�6�}��7��L�����a)B��%P��s�1Q&��e0Il2�nC�+���ƒ��ˀ�j$����O{�2�6�}����IȢ�t���ȣ����vxI��Ί����uŀooU��<t܆{��w
�L��(ȄtT,D�x��ɿ?��μ�D��^�df��
��D����&�}��9܃)X��x UOם�D��{%~�َB�ӣ�FH&�q�!{]��k[� �r�Q�H߱�F0��� ������L��������8��y��u�-���18��3���A���D�u�e3���7l3**�
�E�w^7iR�k��3�m�w���:�g���<��6��I�t�S1�$�=]�)��D�{��L���D{
^�In��M#��D����w\X��${�Ձ�;Fi�xp8
��
@�̆�=]�:$�řL����G���O�	��S�B܆;kl��Mt��u��n3�cR�sv�.�玣[b:�՞ڷf����c窋1�9ٮ���9�;Nj���W@��\�xr�ڳ��S�1,nZ �����,�Z�rۥs�����8�n ZR��!�g�h'�5TK�8�x�F*�$���5	����Dы�
x(״�f.J�B�)�dH9%�M�}�	>�3)�y醉�� �"tU@Y�K�cND0�	���l�%{��)p��\X���8�ޫ�Ru*SS3d�LT+A�ڎ��V��{�Qւ�}����x�9%DѢUB�{�Uŀgl�����a���e������.��*U�$�rv�X�Qփ��hv�XGr�$J�YUiD�T�Š���OÀ�|v�Q�Yb6��T��2�Ã)����E��~��I�za�I���Dw
H�g#*O_%�D���3Sf�1m�v���Lm���ֵ����^��
��m�֚Ca��Ս�zq�Ty8��z{IHH�E������寎s��C��a���@��6��}�4��w g�`f�GZ#�w鞚����PT�Bz����s�{ �D�x��&�����4VF�M:�n	D���\���V{�������H���:�;A�-����P�D�Tɾ��v�]�H��>�AU(�H�Q�P���* �*Ka*� �m(L�������a�K���f��7w���Qփz{��n��S�Y��Qf�<�<[�^�):mn1tI���S$߽��7�A����%{ �G�1ꈘَS�UpD����g�vL�,1�g� !��8���2{��TI��H�0d���f�H��R'����7��I7��I�^�f�V,�F��)R�Ch;�Qր�ޫ {z�^7�M;@'� ۪�lА*�o=0�&�SI�9����Z����tqv��1�I���3����L��e
'3x���*�E!I��j�&#�q"�M�.��o��7�L4I���I�y�#��N4�URuEqI3`b�r���o���;j:�ø�&��B�h�:�o��(�o��_hE"H�	� ����j��&�&��
1�ؐԩAT��)��XEg}�,���粆�X�i\'.FyY�e	�QbZ)����f�zK<&��FV%O����C/=����U�أ.4�%NS���k��=���Qs�m:_�����y��e������٪���hI�s8n�p��%e>R��ƹO�<�Lɳ�T�"���iW/�1
�fJ��7���{(_N6^(�E#I��h- ��͡�,:Ew=�6Q�K���0ۉ��c2 �t��A&s�^�$p�Kek�"/����g�Tt�Һ��]������kS���M�]���C ���]rp\vb�F��SJ(���gkn�^ӓC<v{�v���ڑuy!�BQi��Q���r�8 >�a����g"�N�l����b�U�5y�� s8.M莞�mb�1��`���̮{b�̮{�y^y:��%.Yx�k����������9O�I�<[��=�|�_7���TM&�N�����s*��by�C:q��l�i6�M��]���1�n{z�ǹq7�-�D�Z��R ��9�3jd^nm�ü�3k�q�ȌD�8�r1Y��H)��G���ue�D1��yޮډ�$B6�nH��2r��e�1�=��x���P� ��и�ҩ��3��XBլN6�-�]�V�n&�<�j�<��)��������4����۬gw�'Y����1���\}��g!p�7�s��@Q'P��@�P�D"NH�pE��ø�w����XE��e�4��f��G��Y�e}�s���㺅�k���;��/P���{{��Ï���s��I�Lyn�Ii�&g�(�����m� �hw�ƑY��z}���b�D��8�8�RP����_'9��>26�y�J,a"��	n8�$r	�����cG���#�x���2Q|2P������2LEGM��}�/���S��T������i:N�G���=�U} 9�h ��^߫���s���:�db0d��#*<����ᅻO�ۗ�3�@�wq$���a�|��\���YG���>���L��M�n�t`���e["]�J�ٳʓ��=6�A:�]��6�.$o��#���=�1Y�cM�u���o|���J��z�dL�P�
	��6|��}̡~�0���P�՘SPG#Aġ��+;�D��<='��C��3y�p+���gd��R���P'�ٯ��̮p~�/�{����# A�`,�F:�&.�4D�dp-�4�i�z��4L$�:7�3~p� �2r �ŀ�mt������鉳Zw�w�n[㑈AQ͚l�����@6��'(g&��p�Ĝ�γ
��f,�Ԧ(D@�*|`q�{w�@��!RXP��\01	C��H���4htpv�҅�"�l�&#aaF���B*��мVJ������e��8J2Bp���ɬF����jL*���0-�X���8'R�������L>��{wy�~u�޳�^��iš���D@cfC�$'��5�;<1��O��n��WC6΀��1��˦6� $�*�L�Vq����2��Yr�2Ehb���W��)�D@D\DJ��H�,�9b"�"""��� �I���ļ;�ţ�7j䀥������� �m��Q�j�t��U�2�I �͆��۩ɥ'�d�;e���-[��Ȉ�j{q�q��k)r�Mʺ����K=����d���l���K��^���Y]!�z�E�0��i�����x�����8�&�y�5��J��N���3���s��\<Yr;���ˎn�n�L�SS�!'X��n�;�pG6x�O\�\���Cýa��v�"9�=��n����-�r��|j�]�ø�Y��N��f��3k.����z����,����unEM�q�?��\��� ���2F���2z��&����덮0�s��=pI��ڋ����%gf�=�v�82�]g���'4:u��P*kLv�7	�a��X��Z�Ċ�J�@K��fi��z���ծ\���T��:��\��T-��1δ;��t�$�d36�^�61#ni��,��֡��8ێ'�]��p���x��d{0�SgX�|}<��u�c�Q�~����G�S��B�)�EүH�wꈰ��� !��:��*)�!����"@~5�>���8	���g�9g����r4�P Ӓ*�Ԏ�<�G:����R�~}���y	�w�����)K��@q��V��q�B�R�q�t�u�d8=��8�ӊ�шױ���k�Z�����gƒER�����pΞ��c�����4��'P���ǿY���v��;q����핮/j��v�[�9	C�{�����߷�� i<��}�����/?k��Ҕ�~�����UF��0�	i�#�,�p��[�%(z��~��Jy����	���}揾��Or|լ����fo�k��͖�8�I�h���)N��{��2����I�)߿l��d�<�83A��J�Q��]�@Y�R�k߹�)J��G�buJ]��h#�1p�wfC�`�.5�b����SM�z�C<�Y��R�k5�AٮN4<�Ok�;]jf(�4�y�[�t����㓎�Uٔ��>y���bD�����i��:�28,�y��^Ͳq���Jۨ��U@fH�O'�ݸ��6N�u��m'׽����p�ߺ��}����yE��h���|޵���oYpJ�߽��`�	@^��Ǖ����<Ds3"R�3%�y q�D�N��݀s�޾{����8�yf�NI+����T,�Y6;ݙy*�X���)N��[��(��G�bu	Jw�����eܥ'�=����)�����l�( ܩ	�N�nP�g��_��O�)O>��qJR��>���@Ҟ/������f�R��x#�M�j��k��=޾�:���4{�R��{��`��~��������#�� tBdt�o|�W�З~���	�4�y���)O>Ǵ�<=�-{��g��0�(l)��BP��ז��ԥ�3�O_�k<���=������
*�!B��s^��<y�O87vMp#�x/����'��&=n35�p�Y�O�Ĕ�G����}����@Kc\��ӭ�m��g3N�^	v�����3���w�v{���6M�|Xh^�1����Y�e3�GN�w����|�{��}��*��{�PwNB#{�ou�4��}��:��.��}�)�JO��^���;�!.��_qL���0�eD_:xʂ 6(<�'��y���/䜁�������JS�����%'���߱:�R�^�}���c���:
*P�� p�;�{���8�~��4%>@d>{��}�ԥw�{�p3�=�����g�ܢ]�s�ԥP�{��	��=}��>��JS��ߵ�)JN����'R������m�RPUBJt"u�y�O��\@�<�����e�K� ����)q1�>��q�� ��������)�4��~��R�����f�'�Y�õ#.H�#�q��0�< k���WP<雯�߇{��.�Ͼ�:���5�؝HН���P4�y���)���3�ќ���7�z�2�|R����>��G��7|^	�O��_~�5#A�����R��~{��b���=��οoxkZ�ԝu�k{.��3��%)���pBP��}��#$5�ٯ��5)I��k߱l�y��j.6�N��ӆ(����{����R���������JN����'P4�����熦މu� 7�.QrRH<�$pQ�c�(p�At�d���(�)�M���U��K�eq'��Eo\{��{�r���kW�iMBP��{��,��G}�G�@�P$p�N�T-����uq=���6Z��1������^��ԥ)����%)I�ﱍ<G<���[@q��YL��w��7�f�u��ԥ)�{�o�L����4��R�~���)JRu��>��g�t�y��{"���M� 5��2R��s߾�u#B^{�}�5?(@D�ұ
&�TJ(X>΁{@��ps�����p��{As����:�SiƝ<�f�֭�8=JW��}�~�9	I�}����F���{o�L��B w����,��߁E: T��&�o��J��7��:��5�u՛�`�kVN�͓�J�ي(d0I�:�{�6���8	�f���)@�}���Rw{��ݜ:�7������ŋ����ӰM�٭�[޸JR�y��8�)I�ߘ}�'R���ﹿ�r��=�I�$w��B0)@�P�b���}��~���C%3�u���R�����`�	Jw�^��[��ʿ�[DG%#��T�;)W�8H�9�|�@�{ߺ���)O��_p�(JO|����A��S;rI@Up��z�	�4��pz��=�_o�`��'_}�ߤ��.�g]�٭�{,��ʇ[n��p�J�W=�\��-F����s��v�l��/jn/��76�a�'�M�0qQ��ѸrAix�v|a-����7d[�LvAh�܍㘬�����g��.*[b�Xy�<����~{�������8�yf��)�(Yદ�c�W�JS��׿b����f�\�kcۍ��tn��[�e�H5�S�H��0����\@�<�>��\�'��nc�<�'��腶���Q��q�~)�Z��m�5����P4�]����iO3�︦�h;��v}'R���k�:�
��%�,�).D��5F��Y�jN�����r��<��X�@ҝ�ֽ��'~��~��O��7�ٙ~����T j��%)��O8	�u��pY	J{���4~Aa2Oo=�߱:�� �b����x�[��g��\���7�p:��}�^��R��뿽��@ҝ���}�d'�S�u&y��� p�ﴙ�nC��SB�J\���x/<�j�8	 ]�)deɞ4��+j�U/sӲX���e�|^��_}�	JR}�����)M̓R��/w��8�<�X8~�|��nF㜎�Ҷ]
��u���2i	tY�9���,�CYR���� ���<��ں�bӷX[�ƣ3�T��v�y��Z:���~���<s�ܥN(�db1���
P4px��	�yk߰M@�}ߚ��N�iOs�w��_�$����~��N�)�����͛E�UCA���Dp9��mY���ܧ�h�߰MJRwy�~��R�����{��&�<���f����I��G5k�n���:��<��{���)I�ߘ{�'R�EHT�O�����	?}��Ԁ��y�{�l�( �T���g�O䣐��l�P���~��ئBRy����N�h ����x�з�I:�W,�f�[qZ�W�R�g�o>ޔ�*��oVh��k[r0���E�^�sR<[��F��W�#�ߴ}��	�߷���~{�ǩJ~<��Y�ќ�.�>���4�W��Pg��n�;���9uβ3\����t}��JS������'^y�ߡL���$p{vC��}��G�г�wN�7Ѽ��ԥ��������@:  �a����
�<��)?_����N�iO����Й)I�{��=��
º�}���-oZ�� ���Fӣt8	��i�!� ,�)Os�{��%"�BYQ�@G�}�~C�G<�9��˜���m��I�s��+[��'R4��	XP��G�߸~�A矵��N�)�־�Z�O� ��@�B�CAA�w}�~\G<��T_�5@� �DP�BP��o�:���O,z�7�4	�3l���{V1������qP� D�$�,@n<�����������`u)J}�}�i "87f�S�$�*x-�*3h7�p�ٹY3����{��w�1,� A���]oY�w)J^����	�JN����P4�}��
~� p2	=���8	����BRp5�f�\ݛ�KJP�{�{�W�BS��O��ٿ�BRy����$�#���jC�|@�߶��IƝr�s�f��Y�g�JS�{�߷�)JO{�G�bu!��`&#�K�s�pBRu���N�)�o}>��\����UÜ�7�2]�~�R{��ߴJR������)2���0���)O���<�O��G�g؎��"
�����w��o8=JR�y��8�_ǭ��3y�i�u-S�sj����r��gGw��9�ߐ@�<����~ބ�)=��{�A�%>{�7�l/���G]�5�q���z����u����6�(�s��H�}�Oǂ�hN��{��2�����buJw�{����Fh3��B�5h�����u)By�}�qO�jR��}���R���߷���2�^}����
xG G��L�N	( c1��8��)>��~�����5��&��R@Pw��o�=@Ҟ~����:�48�N9B�U0Փ�\y�O�)��5��	�JN����Kԥ)�y�o�L��tz���	�����%)P:�ݭw��Un��[���B��v�F�Q%���a�+�j�\�<�8��=��e7͖�k=<[Y���I8j�w-��x4dT[q�7��$uUڇ�Sv�m��Yqd��=���T�vKo@v	8�R�;d�ޙ��#ڑ4���#��{��3~���p���?r6�4 5*S��35��������(��XVu���>Q�2r�k��\I������[��y��Q@>y���ئ�)>���~�����=��jC�����fd
W,�����(Je� I6�k{��~$HI%^u���g9'r��O?f�~�	JR{�>��JS��}��#L�(@�+���Oǂ�$�I�4J�	�P������J���A��U"	�(���� �@�����8�)I���?Aԥ)�}k���# ���SD2,����B�(!�{Z>�e<Q6,I$��<�/}�}��ܥ&w�o��]a����'��ny��#��wp����z� ��k���k3yqNK�%P������F����d%�" (IrN��__�����~�:��;��w��JP�	)��	 ��<�����$pg�~�8�q:��a�儳��%)�}}��%��kw]e��vN�m͋�\��!L��k�Dӆ/����83��ߗ4%���߱MJP�ߚ>��Jo���3( ��9�_r�9��ׇ.ph���i�,�y�Gp鎶h���C�{���
�Cd�  �,��o���<K:j@�"L��%4�X;�[6�lN7k�l�\#��35�-��#>�Ak�)0'F��k|,ٳ���1l�[�I�hmИ�RJ���BJ�`L�h�@i4�H����W���ٮ��t���{������4+A3	��$s�t�w��tz��˥���>=�;�lvg9dq����6��͊P�ěG�TuA]T�"�6��Vىj���j]AV���V9�-[�K���-�X��iC#�&�3�<^�D��n�rmY�������I�uQ�Ӆ�]�����T6]�ԑ����6w\S��`��vz6�&��8��J���s��8�����:�j����Kwrn�e��`ؓ���L�) �t]�U�S��헬t�����'��q�5����2[9�T���cV��O9��&
`[u�Lv�cmi쁗fVPVr�!5F�Q��u=c8�gK��@�6�\4^:�5��^A�$��n 7.��lz�znZ��ۣz޵�f��4fj���𾪟����(#Ј�� �A�"��&��v-���H_ A@�w����k�qӅg�����7�����h#����7�W].����0���n�Ξ�b���	�N�!6A+��ս�/��2޸W�x�D+[����!
�o%��'���{�w{�|�7oy�)JO��?`uJw��w��r�Ry�5���e{��=�g�!������'"(Hk�@�*FUB^�JR�����)�S%)<����C�%)�~����JO��^������qFʒ�)*t���8��_~k�:��2Sϳ[�4%:��ʺ�����pY�#�>c�29�p�4��s���E� p����lbR��y��>��J�}���G��>Ϙ��'���M0�5�N�	��m��V��[l;q����⹷d�2�����ږW9����ߝI������1�L�sx�8����@�U���i�n@�L���_ ���� �b�+�R^����M��d�j�s`{v��=�"rML�]�*$����:���/y� �{���٭��-�:	�J��DF.���8�
��S0S�c�M#������"�"?���:�?s+��o��W~�g?�J��O8��#�����$N�U;Fʕr;��~���W����u"��� `�����S4��C~�}�E�P8�T�4�(�2� ?)#"I����~�Ey�߸r��7e��  |8��'��Dnoŧ�rR�s�FRY������.�A! ]�Q���.7�.�c3IB�S3D
��<܅��G��<�����9	H9E��T�2Q��Ē19$q�s���9�9�UT®��9�l���D������s�`ps�9�N~��
'~��?��IƝYf�B�ơ�$�kN�~��J�}�$57�� g�[�#�G.�0"�樐���w�<2��>�����7���_�"e0"�B%M���R(4 �AD� 4�ʃ��{ݨ/�d�߾tO�Ȍ��aWR�'f�J�� 8-�s��m����ϥ�|��h#����}H|�J��"[�F]M�fS�|�.�Qx��� m%C�����U���wt;@���Snl7�0�)��w,F��|q�!q�qB�B�aĜ*IJ['��6�7������B��r�'�3勒3቟�)�%R��Gw=3m>ps���[��=�j�K��6����pq���oȶbiەW�`���tI�����%��A��Ͼ�'�u��mFk�]�ȓ*���ʿ�D�]}�����+�����*��7��]�ݾt�~�[��\=�8����
�UgdE`�L�)f��{"6M�D��Ղ��х�F�,v_�=�d~Sr��㞌�u�Zܮs.��S��B=:'/s�wdф]6��79�;s�t�k��H-֫oOn6ozٛ޵�[5�d_���$�@�߿*�{�����R�K��TT�$�r���9�t	�QEG�(� � �[�S��<�Mfp�-w�ws�� �p8>���uug�:$�z�dn��~�bs�u�ۏ����U�aB$���I�{v��{���<�{� �e{�����r���h�2�W��[�%�'��h� � �dwW~~��:���l��+�~�y�X��pp�şE����AN$]s2C�$#ɜ�C=����Ѿ�u*jjK�W"A\��.��� .������6�u����s�!�DB3���=��������i�2�9�������.��;̥٬���N!@�p��2��ow5�${�m�z�si��n��P�.��s��=�pw�����McD=;��gC��qI#�tk��&5ห�k\8�C���g�K�N�\7�WQ87�Sl��<��Nͱh�:���ç]s���x;:�g��vߏ���OWuf�$�sg�_9�B?}�ﭝ#l�*�%N�:d��j� �Xϻ�y>sa���RWUS���7��Y'��6�&���g��  g?}?$��W��g�-��&���Sh���߿&�� �~_}r^��I��k�Q,�s�Gt�]�	@ʲN?��������6�v]�%N�Ũˍ@�4���i���337FqiͦA��ݶ{�ZCYq�Q�Y�ֺ P� ��k���~d������HA�M܇v���`�n�"���z!�ԵHݕUr;�{�4���|��pTu��mz��'33l_�s�!��z��P8ѪP�T�	�TO~����=̚h�� � C��W���9�}���i����f+���j�R��Kک܆���Hy�2�?|~��о����6��"����[����j�=�ͱd�돿��n��>�I�:�w��)BQQD��K�|A �s�ߏԃ_W�d���,7�PʹW2����FI����#;:�Y��4� <�;�~�� <�~��A�?Ar־�$��������]�Xy���������	RQ!�3��?�w����l���D8eB�d�䩳jF��=͚h���Y��p�<88��Dځ* ��H~��h�}rw}��6�'�WJ�̭ky�Z��*b���H��9��G �  �����p��}?$�dݶ�,j���:~	8������;I皨�F��f%$	LAƑ�-A�vk�z��κ��o���D`D AbU>��D��R ��f�$wF��"��E����lhҬ�����5����D� HR)
QD7�g2�J�?��2��@����b�M䇟Tm#y�5�)��JT�n���帶�� �����
000J�s/��~6I�oߝA{ٵw� �9�< �^|~g�#iAE�e��
�O�>�������{���ͺ��i	Ô�+M�VeZ��0"?}o���@���0/3�߹����J�A�������,��@6��V�bNҩ��Z��d��QMP)pi���0]fk�Hꮱ/Q���@�t�R��o.ɶ[��b���vCBͤ�eW��$�:R���M[Sa�/F9����V�Dʮl�l��|~3V�7o7��_�C��Z��Ӿu�_�;�h8�I#TM�$����DӪ�ai]v2�ص�s�g=:�
 @�
���n�A��ݖI=՛L�N�pk!C-�uu��mD�`�����NP �RGvI���$�6���뇑��7��D���)IM� �*kԏrei��p%��|蓙�_Z'��m}� 8��s~bG�7�s�L�� 7���ݮy!�[��:��v��5r���i�#FR �y� ֍܆wu� �]�l3_)h�L]K��U���`�D�8Yi��+ʓ$�;��W��)�533PT�ԩ��m�hɻ��v�~gH�l2(�RUG^� ��B<�$u�ߙW���6�5��5�l�5���:�n�2���'�e�d��۟O'���j�b�X�������m�KJ];a֩Xv�;�x8�48P�R�n�|��6�wuC�w�`���y��nĉ�����Y���=Y�k��πC�jE���gR��
�N.�l��`�j�(p���6�*�����t�]I�-m��r�|37��b�]������1��������=Y�i�88@��Ͼ�'��i�Q��7���D��,�d����e^ߚԍ��n�%�$"a�����);�n�)-��͸OW�m#�xbkYܹT.�-����H�"jA\�I�*8�u`����n�7�����Lx�m����'PSQ�S��>��n�@8I�����kY�1��XB`��͢'�C�w����2��~Ͼ�D��6U� !�~Ϗɥ��)��tn�f��}h<�y���"���}�[�����jFRfU�V۰d.X�_��	 �dG<���~�+��l�̯<���F���M��e\��B���*��U,�<�Հ�*WH��ġ(�HM�$B�M��K�y�7s?û����8y�8�k���:�Wԉ���e�����O	_:�/Q��a�n��6"��$�'}�6�:���y�~�\� $�v��D|>0(U��˒�T��u�G�y�y y�;i��P�Iĕ	Z��s!SI\����}U���떌��c��nXV! �;�# Ș�7��PUD2#�`\"cd�ye1IEQH�&�2i�9HK1�C$�#E��Z�a�S
�U�j��ƇA9�`�f��F��~�19�?���Hm77�= ��kC��=�B�k瘇��G�s�<��u�s��tf$dtH���E��cJ>MS�{qc����TOY�#��V�
�b�ȅ��Q ��TH��f`fd&�ne\lƖF�e�&�""#��vP-����%R �0DC�"5�3�D� DG1\�$DG]�˥�S#n��B�m��$͗�(����Okk�I����*�:�V�y�so=v������p͠��d۵1�J-j��NN�����=.i�P�&�%8�,��[�K���47`���C�Qʜ����\���E�Ղ�us=����g�#��wl�.f�NwH�✸0
p9�ը�!o7V�9���CHfzj��x���b݃-���$s�c��#s�A˱ZLP�8�{���9��c;�FK��@^��i1��Ƹ�T�I%���Fx593J�F-�I�&��9E�v����lLDB�� ���$ԢS�Y��O�aۖ4r�䋙�rLn�ش�8���,ۋ*,�0��;+5u�\;v�G�b��ʉs C�MX�na�Vf��T���{6ʒ�,�q p��NɌO'gt��av�M!ۗ*�p�>�<C�wA��E8��-�#�C���j��R$3�1���3WJ6t���	��q�rc�Q0;M���P7������UzP@8��E�DٰP�C�Es��>Y N�E����W���Ъ|(y�;��u�uiݦ}��N&�e��R:�M}�߿-n��A��ـg��;���?Zռ�wy��1��JJ��"jSi^{v��c��q���s��e���\DH��B�Q�
	���}�ukw^�$���D����w%Zb�f�4�ڮ�-�����wh��??�Zs��ǽl�=�P����$7~���7�'�D̪�&�)��P��ɼ�<�;��ky�+ӭ;����n���T�'2eT�U�K09>s`o�7��%�;��{kM�4����q7I8�u�� w�7n�>ܚh�uw�0U. ���+ ,�4��3�1i�	���~@o�*{�W��י�]�a#�
e��Kmڙ#(�/Z�Ll/W=1�eL��<ێ�k��#�n-u��V�砻�U�ۊ����9}��[q��;��8���N�vuu=iz�%M�F�t<m˸Y.�l��uqa���?~�8�3ދv��N�tk!H�HRGvI��ڶ�-�b�H8�N[F�bGn��8�BIj�U�~{������\������D���)I�R���w�R�M9,9\<���$VG��!7b.�Ͼ��Ϫ���o$=ܚh���X���bY�i7V�j�|�w�$=��0-i�'�/�4XI�JJ!&�ED��em�ux��""�v���я�4*)3y9T�eB�ϟc,�ɼ�<�w$~�Ƿ۷d��$b&[���N9I��c�~!�׿0�8C��s�rR�GM��'8� �܆E �gs�'=췈5i��8\�d�n�d�t�sx@�G��|��q�M$�	��ļ�a���+�у�Z��nykPخP�nzWncFV?��;���s�l9KcQ�Y��A�h�۽��������n��$Hmsn�d�&o �1uf+���o���'��ͶOu��ヂ� �}��d��j�(p�*�
��5D�=3l�p~�g�P�O�ٯ�D��[@ �xo5���*��8
�!�<;A��{z�~H�o$�jR"��QDh�1)<jݩ�e$}ɵ`{��䇵��{�5$)���j˪�9.�Ÿ��'ԅ�`�p�\.�"��[h��q����#2L�+?~��� ޖ;A��ǈ���s&�?7v�|r"�	,��Pj9r4܅8�{������ͦI��w$Dd y��)-�NT��fs��f�}u]���9�(�`Y������!����*� 1 ��Up�/3�Ͼ�N�Ŵ��ͻ���������H�����U7a���� �t�>������!���rw���r�e3*��J��x>�g&����g�l��d�k:�-��G��FJI�CT"�Ź�Wd��������jR���t��Y�h��(�0�������?R&�6��'�ɦ����F�*��H�E��!��$	� J#��R5ޓէ6�����uq�V�<���IP��v�M�J�<�[��n��<�Ny���s��l:~��c!�i�v����h�f��"s�ݻs���88� w�O��'3�v�щ�EG�+���M��>�߈�kv�����<���9i���9��$�NM]e,�
�3�y�����X&�pY��/:2ٜ�@S��@Qm@���pg��|���Z���"7��J���qS%lx.��ݹ���u�r�}�=�d���M�L߸8��@#�s��g��D��!h���b;��T�Ud9hs������5=o#2>���<9ČߛA��$��L:D��}�`Ln�ݖ�@�n�؝ �B��K*Ĺ#�?.� G8��}_$��~��qx��0 EUH�!��qډ������쥪����&�3Z��7l�W�ݸܗ	��
rX���.Z�����K����tt�"�`�n�s�t&��rsE�u>Kdk=r�C��[�;Bt��c��R<�qU�͸�Nc+:'u������{߾ 3w~�g�ē�܆&i�@���${��h��v�4"'15�9�͌5�@4������|#���Z'����'�Nm0o�����wWl��D�YRD!2$ED܎F[wd��vQ'�ɛl�ܚ~���I�3����e�����I�U*��=�S�(�5`g�� ��C����Ó�6��˽E3��Si�����9}�6۳�$k�p����$�u0�R��8���? �ٟ}VI՟|�ou<����7as��������8eѲO}�m"j
T�I��)#{H���q뮇���nw�Ԫ���y q�̀n�d�riTLME:{�rT�v��&�ND[M������T ����n"5�W >���ͮ��{����ތu��x:pKvs�lZ˄�/njz9;�ۃ]��gC���.�����`��`�[��s�l=wȏ�������W�`yi��#=�ـ{��|�r����ɤ>�F۩T]���;�_� {z]���޷�k�X{<3Ap8��wlѹQ���8�����ͶOW�m3�s����o�dߑ?)���,�4)�h=ϭ�He�F+�P��A�nSh�;�:v�U�jk�/��O����H�.ўc�Ө�ʠ�6�\9���ouR���%*�J�0)v�e�gl������>~����Y�(�Lʎ�i�.\���}�z��8�4ЕD#���h/��3�/>�g|���7m�չ�W�{ﾇ�)�mv�ݻ��Tf���jR�>y���-o� t���<�-%%%8�J�=��m�{g�W!��m`A�t�����.�����=Zsi��Z�@�����yM����N����5E_�e� kr�y��r_��+��*|^#8,�޼�ASH� ��HC\7r����m3�t�Ĕ��e�Ғ�['�����#����_���sY)G�r�HQ��I)�J3%"{���D�shQ�x�a<�����3�z�$s��S>Ӛ�IR���.�*i,�<��r�o$=׺����l��Ǽ��EQN8b�j�=��5�,����!�S8�!ڸ�M�Z��o=9��{��s��j_O}b|�,'|�]R�/�௱�}����%̗i��-�QTUV�N`i�����Njn#�p�O}�}��7>l|K&�3�*&V=�y!���C۵�`n�w����#�,��}��Ue��vO�ߨQ$�R5�e�o��`s䔺STR���U��\��O�`�
B���~�[ ����GR��l�88 ����c���FS.�6�ed�T���"6:�$�Be�\m����ڢ�W��W��[Q2�iܭ>{H+������5^:�:����(R�@�x���N�
/A˩��'dy����U���s\��hs
U�:w>xL�[k�@q�y{Nh�wۈ=�'��*�w�I��m2.ᲂI�$&�5o 5������x��f�1��"���	*� !��~�<�o�,��<D7�&I@��+�%���j��nL^��u�k�����nl=��Hy�j�5�`�b6ܷr&��'�N�|89�8$��T�%T%]ן{��, �U��z�#�6�h��U���+[���ʯ>�߹�W�{����VPBQ�!=�߿u�^g�~�+���h�H���wFEv���d��ߺ�+����j�	( ��!�̃~�E���@Ā�M$�*	�&��l�� �|�B��Ka�������]����ꎞ��?���}G�|�� ;�]���h����3�눛�0�	X`�Ō0�%,(�	��� �!�$��N�1*oF�(�!�
JZJ4��	1G;v] ����HC�� ����]�v���y]����aw^�=�7�QNa�&6"a�������]����
�ԙn���h��[+��T*�+���WU4�Cj�*:�-E[#�n;W[��Nq��kqԬ�ힱQ��%k<(Q<�QH`疭P�S�ەc9�vs��F8o!�&�ԱPq�y��6Hi+W]V�K��`N�ذnx9�u������.�IWf����v���DspD�����n�F9�M��P�h�.#��P-�Ӳ�C]�r�̬���u�M��]��$�@v�N���θ�^��b���r8�	ɂʆqJ]�H��jݜ�]�ɮ)H#v���<p7:��j�|J�l�VPm�.c��a��m:�P�JH�i��I��\���3��q�@��"b�"=��p�(�<@�P6>#��A-�]}�v��zƋ=;�JT9L+̷�ml]t=Q]�+�s�ŷ%qXi恻��b"]�x(�x�=��H��9`<�zsjT��s�dDC�E�4�08}�o_�]����m���7� �x<d����d�>M!�6�H�"���&��3m�{��D��m�{��+���p�w�ߋP��w,MT�W��O����Hyw9���l��j�8��RZt\t���s��/ߧ�￿� �_��!����@{yՆn��Ȝ�+�ۻJ�U%�K��B�"8{=򓝌��v ��bS��52ML)�P�O>�f�v��A~�ͶG�fȢ�9RTb���["q&��M��\�R����7קZ�=�P�>��Lws>��r�Z*��ݚR��ՒO}�* �8x@��/� Fg�TŒ9��*@) C��-�T4E	�L����B�Ȟx(t���ve���~�U��6�872��HxbКJJI��$%`{�\�C�[�>XO�~�!��>�x{9��"
ꤦ$1AvI���Q#�zkX��܆{y�ԏ�p	\��&h��.�9����7(ը�1) H��bQ����s��"f��3���}6wS�"Cˎw'p��S�����Cc��ƕg���
�T�SD�*�W�y�C����M�����~VH��kDT�
�QS2+��ky���7�Q������CV�7�s��U38]fV]�4�`yq��3��ߵ��A��L 	��� �S��<�9��{�;��D����ÏyR��F�p��tO��,��Y$��禎}���4� w2��7�!n��2�K�ʦ�>^�tI
S#���T�E���qù(�Jd[���q�������s����7��0��R���}�w�F�7�܎,;��۠�����j'���؀�άn�4�s��I>�ͦ|;�	����0�Bn��uC� �j�Z������Q�#�.���Jj���J���=��Ӏ{���{���G���V�j'�)UHK��N�mՓK��g�6����{vA=̃i  e�zBmH
qD�ʡq�ŝ�����W-$9��3g.�l�ds�L��Mŧ�'M�er7OW���lv�ط;�g��x�Ι!{v�=cqɧj������ġ�6{N��5��8�t��j!�`ȢLm6�8M�Z.pM�|7j��=��RR�R��r:$�f�&ĭ�髊8'���6��L�E��Q6S�8���/��u���5�'��I�oسJL���*�pppJ�v�
)��ڷ �H��=��w�w�f�{ ��hh��f n�w!�y���z��EJ	�34I����9���y?�C���`�n��M��bn�d��f�J+0<��`wo[��'h�Y�bͬ�j��8l��J���J�ߢg�\�C����j�;&u��'G���I�J�ٔ$��I��d�TA�s�QEk�jS��B��))"59�1��{����m��ji�Fӧ%; g9������{�O/*�sv͖�=�Ö5`ݼ]����=�]��6��^7�;wi�+�MI��r{DG�۵o5�V��f�����B���<���ep[PF�	�Z(HА)B����Œqn-�M�o�p1{������J����Y2��H� �\����曹l�������������b��������`7�6�Kb�G�DaL1M�T1���s��6�'��i��8��oݲF�[�@��)GN"��'�zwm�L]�Cb2��%
A8�0!J%P����H�R�fi�N{ӞHj|������K	����T�H"�\/S�v{]Ej�w������v�Sy!�t��j�#`��%IE�"
�y��j_7�� ގ�H��V{��y!���+{�V���.g/"�Tf���J=��#.�6>�x�Ԉp	\�ԫ
�D�z������{�N�PmՆp��Q�vܰ]�'#�'��m"v@*p��g���K*fz:b�8�(�BH̱}��Y'�qm"{���]%�+؊��F����8Ĵj�(�����A�6CFA�O~ݯ����~�m`��r>��sB�݄��f�D��;��_� 2#��߮C�����w���ӓ��2*�hB���z�g9]����+��ߵ�B��$I�8��R3�c8�A��EdJ�F� �Z��~�O����v�߾��G3H[��]�Wq9,�Ux曹y�<��V��#ۭ�%�T��-�4���v�Ws��p��D�j:�꽎��.B�E�ْ� ���?}L�} j�sa���I�sX#/�m]�6��g��Sukw��~Ϫd��k <�є�B�쳟�O蜆F)S(�TIn�;�6�������� ps����D�����'��v���Q.�SR��u�5���]�l7��YԢ�FTD���ퟹ�߾�����.t$P��]@�)��6�o$��� �shM�a1���;�������۞��m֑Zܼ�����U-U���;bҦ�Dp��'��;��ƻn`���N�fA{LL���F��OS�fыW-5σk=Z��]w��6H杝�ٴAn��m���5Ӻ8B0�.]��b���]:�-�s�ǃi�Ɔ���۔�4j�'�ۮ�;w\Q5`�QD�����E�
��^n:;tS��~{��� �9��~_uf����۲{�c\�l_�>��n�t����ct�ISRQV��j��ά{���ps����_Ԏ���
AԊ�8�-�eY'3 ������r�l���uo�Ή=��ݶ}�����q۠��Ow��~޸x��Ts�ͺ���ne�J�n�	t7d�8ۯ�D���vI��6�9�M�g���"��RRAJ1#(��zh�d��s�_h�}e%��$d��WV�yN1�([J~����D����Ow �Gك4�	QK�t�
����0�0�E1�lt��R��ocۢC
.^W���mt>�q�f6�[��fD�c��Ε�586���v��@�GN^ب�zm�,���#�`mՁ�us�u˴v�X�ˇK���I%�*:D�zn�� ��?������ouC�k��!Қ���We��S��T;A�u���X�L�da�z�B�7)�r�� ;�Sk }��>�t�MB���5��r����n�U5ud�fA��uT�F����N٬5A�mz���I)�S{���2������:bЋRQt��DD-�
q�h���p:0!(7P��&m�O��i��� i��ωĨX���M���|�wk@��|��E����I��6�;�M�|�<��`J�iQ-�$�7�P�N�o'w!ۼ� 7\�G�Û
QӶ�X�Q�r]������lw���!�F�ԱO�?F�.�����E�)�fH��m�EʶB�]�\�2P�j�O�]�M�r_���JT*�|��T7��	��Ox���TE����LP�Ɍ�p����!��Y�P�ՒO��e2s��y>s`g���497*&R��l���T���|�0}P���<��j��;�B�&�ԱqI,�PK�������/ �{��A$�(E�I��B{٣4
�i��cX��4E�J��f͚8#BᩂI5����y%aF`���KA2������8!a:�w�J&������,0m���	�0���N!�u���)�'`٢�Y9�z٤���։���'�F��)
R���!�����0(#*2��VI�����ɬ�DSP�H"Y^N�Z�X�e	���]�ܖ�.���3z��4�A(AE"�B�ԫ!,�%T�r���2 ��qb
C���8��[U�AM-$LYDK)�a�QK@R`aX#ŉ^�E�&� �F�� &���}��[�]yf��,��	et��f�
]9��K��[�9�� �=�[f��3� �I2Sa�m��6�*�̼�322Z UO@Q��U�.d��(L$J�[�T���.̫<�ʳ\�p�E���Ȇ*�/i��XJw4f�qnT��.{-&-�ʐd�ʻ��W]TS�ûE�#4��"�,MJ�%P���5����	�j{�X�Ƞ�Q\H�I��^�r;j�vn��y�#�Ny��Å��imqqb�n�.Z�|j,u�\4����(x��Y99���!�n��pl"d�L`�vUvٺlL�x�
��4�\gdMy�\�̫r{]+ٌ�/V�[m�6v�[��n�b8�t��t�<Lq;��:s�Du֎��V������;r������1�	z�h:��X���NWv9�L�ˉ=�Om�c��ۦdԓ�VF�ʀiQt(ς��Z�n�V�5���l�G�3�)\�����+��ƞ!<uֱ�=Xݳs��`5�(n5!X�=E!�U/{	��W��B���2��Km:����q�÷xm����%<d��@("W��D��m8:�cEeW��<eKpZ�C^��Z؜7�������֥�;c��������9�K�Ƨ��qW�G�%�@	���(�i�88.ΐ$�PH�C� 	P�TW�k~���{�.��~�/�ɟb����vd�j�ɢb�}��'97r�<�?F�T;F� :I��j���t»'��Uab�E$PD�M��s���k��c"7l�fQUQ*��l7�ڛ���w�`7�)t5���O�Gi�tmA�L�RSTT��\5��������I%yn�9��=�&���JN�-L�{���~���#��d��0��ިM���\R�
jˤ%iM�����y�n�qg���ަ}����_Z7w�C�EH�We�����V�܆oW5�ou2��s�g{D��(�j8#,�$j8�Wnݨ����T����\��V�pvv��/	���8]�8�ket���=�7��T�7�q�;v��xؚ�f�n-N�26��-��v�� ��h.�vx<A�5�.�z��e8�����8/�}��l��b��2H��J�G���=�vI��)?d1H����<b��T.�L��*W���}�2{�}l��nТ}��)R+j]�Q�D�H�H0�&F	��n�ո��1�� �ܝ����`y��Q1U��m�	�w������  �����N���|�֝ܙ��fh9��V`n�q`?mG<���3����v�����"��NJ��B\$�?����G��[�����ο��y y����q̕AR�
��S3� �&�C��w���W�dvol��x�-�K�6h�")��Ͼ�'ٓMs��v��58I�U�sØG9�� ,x��=%������@bEIp�P�ܯN�"��8<��sŰ�UԳ�7AT�^x��/h�zpKvP���5�v��ƾ��S��]��]n͸oqkzȶkv������!`YM�N	e}�ل �K���g�舏 �u�a�G|D�5D�K"�rJFI���rs�� y��A��y1�~��8x��?oȴ�!JTUL�D�G�d��ܝ������6��)�\�X)��.��f�oS,}\�k����jS���2I�~��ߵ�F�[�%�(���$�zn�&���+�v�7<����D�!�����r'^�f�$�vn�&ֿ�g��cZ�AZN���6�E��p&b%H�`���$e���'�_*����Uw�>�"�	Nr�߾�vOډD��bT�)Q4Z櫯����?
���D�]�}��o�X���$<��؍�qH�A3�o2�-T�����L�ﶶ��9�  �8��M�����9�R�Y3b�rT����s�y y�V�n�`nҖ��3�'��M lW}��\3�r����vK�e�JNH�F#a@�3�A ������1�r�����Q2�Փ6�(P�`��i�I��E����g�����v�o?�#�5|?��7��s��� S6)ʃ0kuq {�7��s���{i���C	��ʰB��
�O��l��͔ss��
��� ��C�y�!s���]uT�`TG����?�O.S��$ku`y�7�n���*j����3d�@����&�;��]�8{E�f`zT��e�Xb!�8��n�$�lͶN/f�'ۺ��bb8l���RB����q�1��K�)(�+��f��1�� �|�×�qo$a�.&�����)M�\��o0��`w���V󛔷ڹCD���^\Na4f��܇���0s�v��y'�G&�I�GE�J�G�O�]�a��d�f����}����?*;Q	A)�J�B5H E2��{�s��k�5Vn��+ �J�UdL�CF��LN���v�wn{��'��rS8m2��L��Z���^�:��u�D"]��4�����=7���FN	dηn�zL��ӹ�Ȝ$��g#��4��썧L�&
���f��t�7Ճ �LR+jXHP�h��|����aWh"	F)��N��˺p7�72�.��v9�ys�{��`{SL����������0|�v�+@�عS5
f|�~���$6���:7��~��|��s���n�)\aT]�sr����H��,ݦ��E&��e%��&B{�ͱd��2/�W�7r@ߟ�a��*�*k	�"̩��0k�h=��0Is�h�Cy'�Ƞ�6$�*���}�M�d�ʤ��cus\9yn���]�ZI�����(�Y��r�瑀y��hߏ�}�����\����!1,�R8R�a���HNT`!}�F�[���=cE�+¥C��+�:�g�\]Vm�lNe�'N�s�x�X�27�D������y����v@��m~v����5Bp�Ր�HUT�$���֠�n�y��@��v�Ϲ�h�D����]�ԩ�RXv����r�X�M��Y��Y���ϋ.�JʥE�HKI��>,}\�~�����?�B7����8$��)��t������ݲO�}���7���rg~})̨X���)T&�$��6�2P��.6�e�HܑNO���%�k��Q?o�������7\�N�p	]T�we�XKt�ۣn��a��*&�܃�o# =�.�{�����,7�l)DAnөb�JR�Ouf����"����� w.w!�m6���j��1HP��J3A%Z��{3m��u7r��F�˴=��Љ��U5�*�JY���Ł�����s��{vN%�,��7*�u�P���n�ߐ������-eݓ��M��@�H�-���POg�V�Nw+���n���D� �����"�7ۺƫ���~�~���CyS�s�x���ŀ����F�p��*�����ܑB�n�����r��ݶOu��s�`��B��Bj]�uQ&�Գ�>�Osٶ,��  �s���bĄ� �Z��. 8Tr��L����ROI�2���ڋ��DX_\<@y��A��� ��l�}��=�)ҸU]:%�vK���a���U# P�p�LPS��E�Y!��m�C�'���͞���:�}�#�Cy8��P�����N���!
n���S2f����y�q`=}l�k�})n�#aeDnS�\��Wd��l��ď���ȐߝGփ��95*J���V�+�������m`������s�}�(�՘`�LRGq:����ՒO}�i��l��͔L��F�mA�A�:T#nck�(�Z��,6ƭjg;r]�u���E���y8��Q�&lkץ�8���#�1�bJ�N�;t��F�j��KW76�:�;J'Uͫ�`�k�\��gxk�Fؙ9��$Q�6ÎO���m��,LHIP:LG"�M��ݒP�%��\���V����v�UQ13PD�%O�6��sX��(�ẒZ�������Q$\�8�(G�@�Wd�7hQ'7�Zl�}�i4��M�mw4�48�ԪaP�����N��C���c|� ���L�̕MN%X��ʕ!x��V�i���uC����!�55%
�UIJn���o$<���=�ӞI�u0�k�d:����˺��%�`��������{�rk��g[f�16a�1�	�+7��ZI=��D���6�;��!�"c������W�� .�/�Y�Ug��6_�|0,r�M!2H�ִ��fA��P�`X��ܰ�b��%�&�r7�\G�LI`�u���C7�ʋ0��4h�(W0��X�	��bF ca����G�ј�K��c��a��@%	A�w�6��`��
�IÂJX4Ћ��	��X�C��M���d�C(�(���H2P���
$��#�:����"*YH���������*j�(����Btac*mm6��▌� s���Y�yG��~0�o#��B�`D����B�+M���\l�"9�i�P�
����^�!��-�g�J҃D�WPAA�֪�:�m�n���������cn`���zX�v��#��ŵ�ՎJ^�vʫ�s<�$�n�"���l��P�r�]ѦN�����X�Tv:�cv��<�ɸ	�����@c�T�����,�P]�X\g���r�� ����kD	�P��s7F��p=�5�vstJ�`�p�#p��۴�9����5M��u����a�y��q�[�����q�λ(mQ�:��mK�p]k�dɞ�f��B��oW;y���N�2=���0v�r�bwA�v̬mu�rn�Y��C���IB�q��}�w{���;�U��
&��T:���ߞ�_o��ΰ)�ٖܽ&�� ��-GVN�g�L��^v����nWr�V�v^̊+V��#��y�snc��\CO�������w����~m����v�su]u�����)0<�n����=�M��	p���&ȦI7T�0�+,Ef�T;�B{�0�u`k�mg��P����P�VM �����)����S,��r�sn��Br�%9j-\)��Z7r��� ��h1뷈�s�P�mT���P�+^�k ��#!j7b1���k�/8��pI�� �$$��囬���݂NfM4Ozs6� �.7c��s�'Q��8���D`%�/:��H�N�Ϧ�׵�$5h�ߣ�~�A�<����_'�2�E 4�f*D��kn��>c�9�8��m�$�a�Iά�ؓ�jG4*D�%%�Ԕ*����zcz�5n���\�F��I%M]U*i�%Q=^�tA=���'�6�����1���u�,��Y��K�Ud�Q;���w�v�4�&����DR�D4���-������--����~�v9�4�&���2;�x -�*��*0��6�<�71�\���>\��䆭9܇���ڎ�ls�:!F5�R���Y��ۛw���;�2�';��d�q'��q�r��I�*D�Xݫ��yL��8<8����6J�$��Mm��T�TTV,������������'�g���z�R�g�p-߶��cZ�'UT����2s�L�d�n����F�3t�չ�$$���7QH\�s7F�{�7i�O��������)�A� ��n9)H��$�e�\7d�^;����;����-v�x��r��5Su �u	�ܡ_ 9�'|�i���o�q��M��0G�)#�V"#�9�v�w!�|��~���2��L��:�
�UT��"q$�{����Ŵ��ܡD��.���&݄#6�N+uΑZ�U�gq+cJ��W\��;-;����������D��u)� ���M �G�I�kXd}�pX���w#�kuh�ܖ� ��Z���v09�Bd�j6iG�0�q�s���@[�k��Yc��������w{�߯�~��#c��ŭ�ժ���N��{v�s�p:$\�[��i6d"�Е͙ȥ���rU��n�j<�[�!���0`8������'=�#�����W#� �����ˆ�C������oy6������1��7
*��;A1{q�T���o$;���3�ܛ�GL��Y4������{z߼Z7r\7a���a�}��F�$QEu%�ųdݞ�6���>��v�X|��o�4���CDG"i�M*$�XݦMi��Ż�����Am]�!4=�*D�LT�_�ǩ� �o0Z��wy�ѿ�����uu�����p )b	!��$����e��P�h�A�f��e�)�
I��� �e�&g%�J��YI!�P�RJXV!�&�&`�	P�`���I���	�j
��*jq|�7�y�F�k7fluۈ��g�,<�8n�ݹ' .�.S�=Ham:u���lǰ�;R7)<��np"�l�rlӷ��Kkx`*'j&��&֮Q�խ��Z�n��c�^'��6�����$�n��Owr�;�,b%2QNP7"�;���Ի�Y`f�j�7�z�����^ߑ��a8E�"�'0ﾛi�G<�����&�����N*&f�l�(��*R� �7���V{]�F-�l��qH�A3X�e�b��R;�6��:4��f%$	D�0�M�"�RHDL��	�9$��=���dk����#��r�
�R]*�	�hIc�q��Q�v�?!�6� �ӝ�y����]V\5#p�v�U�qP���M5y��N�&�(�	`b	灂.�#�`�M��!����%��<D>�̟���w\�{���5s�Q2�j��I���Q'V�d���)|9�^��}���������(H�&��%9W�)y���on�e�Y�ڰ�{��ِԦ��#J:d�=3m��*�<Q�]{��f���1sh($����u� �t��'��H�N�B��i5Da`ƒ�"j"l#�[�#-�'�s]��I��&��3���[h��Llq�%3��+6[V�ޯb�\�C��v��j]RUQTa�s�P*�=�P�����k�؋J� ? �D!IJ3("(A
�U�t�f$*��e��[TT���9�s�����~��D�a��"	�*�M�!Vퟸ�/�d��l�щ_�ݩ=�V��ԨT�W91�U��f/��_!{�)��)�2@���ź[�'lH�G[��������۾�H��f���i���f�j��q�Us�n��t�uk;�<���;g�n��~�ߣ���A��|X|��?��H�]���*�I�f��� C����:���D��)I[�k�A��UN*�'y��l��N��?�>�>��v�G��R(�����/0{f�$��̦I�� �z r�Ԅ,*R��ԓ,��]�K�Rfz(x�d��:==���K��{)�mi63�B����T=���]�����/n;g�͆S7c{J�n7Z��c����ܾ�'��w<�ep��H�y�5
؆�IV6k����{�if�<��BIH��]+����k����6�~��s��4�r\�2��(S��O���7����̙���<�D�su�$Qے�a�[�Cл\u6��6U�0�y~|�h=�L�7��`�L�@���N�D��*��W*�HUp@��y ��v���Uo��h���N�$R5j��ųa�g��3�_������Ke����Yd1$B�iF)�Ez��i���2�3��`���s�覄B����������D���?�	E$�MQ'7C��<�y��iЧ߳>��	n��L���i�H�yc(ɒ���ޭ��m4�4��r�!	9;H���i�9\��]T�VҜ`�@�=S�Ph�j��64�ð�8`��aѫ�P���e֑d�����  ʠx�P2؍��,�D��������_<��7qg%�Me�_O����.� �U�Y(�'0[�ߦeC��^ޛ<�I�.I�E)����D�QR��g�2������:���;��᠟��b�2n�*����r��`����ôFGA�8��3I8]G2�7ݙ��t,_�8�6���ƞ�M��X�$Ȣ��	&Q3����ok��3v���13�n�U�Tː&�
I ��ڄ�7M�b����4A=^>�d��̦M�n��|�CA�ܪr�)����ϵ��;�R�XX������,s��?v�(��o���}�3i����5%	��̚��0wT;A�m7����c]��=�QWSj��R*����y�v�5�C�}��[��ÿ�/��aG-۪�Q�c6�?�������\���v0��+<� �f@���$lH#.N����Nw&$�~����Ğ����NO��:1�ek��-m�Z׎��)6~���֬ܻ�$=��d���,3y�uIUEV*��XLц ��v�;[�vxe���_߿~J��d��*�"�h���}��{�i >9�ø8b$���z,�c�b�0HL c	�.&�8���i�x�"P�٠��2i�W������j�f��4=� a�̑@4!�S1!���5�ܰI�A��W| �p���:�/(��y�׽f{�j����x���P�D�/��%���]G���$�/\�9T-�"�vK�K�7Hi��N�����,��� D[bb �)q�K0f�#�2EhI�""�C�����H�D�Df
yD�����|�HlW DnJVK�I[=����#S�c�^�� J�2LRs���Cm���5{ ����HF��ܭ��[93iUy�3�Y�3I���7hĝfؚ�N�˔A�ٻ`ΕM����ח��m���u�89[��r���s:��8�j9�.���Ӽ���r����N�֜�^�2;�룃bC���ڪ�&n4I�綆tܼ6��+v��A�0�	*��Ga�[��n'���͇Ǩ ����\#�5qY�:B�붚�C���.�mO9ዝ���i��2ӕz�Y��/�G��^8n.�>�2�Ӟ�F��Q^j�MԒ��5\�t��Q:�}=�tm�D��n"f݊�x�-��Fޝ����;�����#c<W�t�ۦhM:���m�����IT\$����3H \�Eք�Ŏj�+
c�!ͱu�'����lh:���t�n�pEEϰh�ۡ�k��j�{U������dq�WA��"�%c�v��-��]ۗ3va�g��c{���Tݛg59�ٽ�n�{�{=G�P��D{����#��!LQ}@N�O�C�NHT.k�6���2o��?-���Ί)Y791xU��f�w�c��g�{[��[L8�tc�LH�T��٦�5P�p�{C�����Vg�O 8��NG$NA��i�H��ͶOu��GA�9��ګ�9O����!-����(��$�؁@����/��O^�y�C�wن�O{bQʢ��*�bnb��a�ky�=�;A��,ݮ,=jE�Ma�*�Y����H=�ܬܻ�Cݵ�$��9(��������EE�':7rgze�Hn�<��������a�=�R鮍j%��ڕ^��Fs�(.wWe�*���,��fڀ���e�BMfH%�ri�ɓ�d��Od�e�G�uala!�&�sU���]/���y�u��ut��%�N�ӣ����eb,8v�.٦C#��&g9�p�� ?R7��j8�vܺ
�&�r���ɦ�?����a4Y/jx;u����*@
&�f���	=��}�Zs�9|�;<���_5wò�Q~l����I��C")�4���L�d�m
$�ݦI���c���[��RQ���W�~��ϫ����h3���2:wu�CD(�TLSiS'�}��'����y ����z��Ve ��
�=�U4�܃��x��y�3 �D��,LF�2SfBjᔉ�����������񫔧>�]>��4 �L$H�4a!9w�su���[H��̔O{��Oad;q�o��@' �������U��e���P�r��vOj1����ٶ�V��J��[�ף�ך�l\n�9�����qJp���uq��7tvN��]���{��������^w���)%B���`r�s`���v�12tA�N����h�y�Mo=Z�r� �cw#�7H"Ubɴ\�b��0mՀ�i��{��V�6ut`8�F@����q�����7m��<Ձ���f�GZ�5#�B�˺��1Ev	=Zwi�R K��p��*F�I��ᶸZ�/a���{US>�iڀ�ޫ�k�I�˜J�&f���`�b,��trOq���M�8��=�Ds�2�'�������#r�����~��i$NY&U�W�{�g���RG�Wչ{���]U�iͦOu��| �z -�E*�H(�u?�C_S,�mX��V�( �y��vh6n���4�H����D����E+�w{d��l=ndtܧP��TI��N���R�V����O�V�=j�����-���� �S,:7��)*��}�����U�뭻�%3*�j*&h��7[�wi��է?��s���~�D�iA`�Dtd�l (*D��7o�s� v�����':��"O{�+@�5����TM]*�R.��$����r���Ϲ��@O��Av���<ݔI����g<��i����J�G�s��-��ƢG�����}=7m�� ^}�p���3�ڻ����O��i�G��/#[m+��%�Њ �b0S�H{���I���D����ؽ��GT@h��pR�xLH�Q���7����d����X�Q֏G8Q(;M�̲U�=[��� G�1m"N�X�s�k�55RBT\�ݕRO骰<�7r�uX�M䆭9܋|޴�2>�5Q6��$�v���d��U�}���x��D��(&��%a��!�hG�����a�u�$�LF��nLi����M�Nz�MJ�Ý��@�DZ��]f�\N�y.�<��`�������+���ۀHE�����x�P.nrٌ�]�-��P��;�2˖#	����Je�X��\�r\T��U� ����=�X��FU0YJ�T'=��d��*D����)����0�.܄����^jԓm�`?L>��3��.���K��j����༻�躸-��뚦�U(�(F`yh��f�3��,{3m�ӻ�2�!E�TlSiS'�쨰9n�����۸�{��!
�𜄊������0Z7r��TH��bb4Y���TȅE���d�iͦOw�B�_s�=y�i��)�!�T�0+d��ТJjQRے��\EAv�ݤ̵rH�r'y���D�t�)��{v샸q0t8
�J���r��ڤ�b�C�v�I���u����g`�V%�g&M�sKjv���Y��;����`(�ކ �;�����.x�g���q�Q/uƉ�a�Ϟb�QU+$=��Vn�|��)9�ż���E�iA�#6,��1m"w;��۸�<���J��:g�U
n��E�Ԓ��7��^ գw!������D�tbgdP&�]X��Q]�X��T��z��座�C���F�.pI$��*�m(�|��Cit �]��d��wr;��U�Q.Ѫ�T�S�1�!��� գw&v���bH��бj�$�m��9 F$B*f�\݂�Ya��e���Hjg?��>�6�31耶`�����{��y�_<�G���u�;��(��`�D��<�k�bE�ȅ�*06n����%���~���1��!�f�M������*������a�I�}�����m�X=�7�MX�2&o!���=Y�iN���E�$&p�d�s͵qzz�������,u�n�y!�[���H�@�c����N<��U���2�/U˛��Q6��r��y�q����4n�ϡ���dS0�i��{�$��M��}H��zn�>���"��pʃ{��9WY����uߛ=�|(EJ�JG9w��s@�뙷d���g�;�&�cr�Ud�EBȼ ��W n�s�6�,?s�,�ϕ��4uA$�t�lRj�����K�E\.�Ce!J&�AW�����:�nz�~??�ۤ���e2o��)���F%��b�:r��'Wj9�I������9܇�k� ����{��$��j9��i�"ÎQ'�~�D�]Ŕ�۴�Hr�sa�nEU*����2����`{z�����>�I���`.}l�z:���e!A��@D�'�zf�'����Ty���Yډ���YXg(���I%C��y������Q[�r�(iX���j���
�R$��F��7Q�n����578����-�J:r�������8q9�]kWC�F���L�BF���1���M�/3��vh'=�� ��.���*< ������{�0�L9�[����vN/�v���.2b6�%�T6�Y�F�ӫ�m��7d���|�Tu�~�oB�9RD���7o�6�u��K�H�.I��I\��ŀ{�z���0wT;Fs'�aW�e�E�	f�nn�ms��n�1o9�D{yZ��D�V���ͅ�~�o[�{k�Iu{.��A=�����+�Os v��&�C���a��!�]}�s�>��2�A#Tɵ��D���z�j��z���49�A8�D��W�!*�3��sA��o�ՖVq���XRҖ��/�x<�l	�>=�a�.l6Z�`�hLR�Z��z(i�dZG!�� �"LX�#3@ڡ(`���1LMoh̳�g1,�
##3	H2%�&kL4�`�Bda�c�a�Ibe�of��)
D�̇F§2+-	��BZYff����@�@�ж$���4894�E�i8�;JZ6=�Dۡ�/Bh2YJZ%�!�E�p�0պ������.��\���~������p�n�rGn5���Z�l�%IZ��-H��@���]PR
U�Hhꪫ�L����S���3��5P�6��ŋ`r���4Pn[�8��=���f��+�q r��8ۄ�a��ˣˡ�pV�W6g�6[=���K ���INx����]t��ݮ�E3H��K�2���$/#�2p��Gg��Tu���nx6Wv�v��hM�<�]��#��#�6��ݵK!���%�z]�"��xXvY�]b,WHh^�ǲd,V�s;����$ӷ-�M6�N��!JO,Ӌ����8�(��N6{]sʻ.9��e�ؖ�C�9���-�YyY��1���]�_Ƃ�8�ou����� �x򀆍)���Ҝ@C��+� �T6
 G,��g��5��z3V��d0��eЋ�!�+N�)�ggq]-�51̮��:Ӯ槙�zÎ������R8p�����w�{�^�����Ӎ(�gZ�6�*&�W��5��Cۼ� �uC�yo:�A��t�RT���(�y�w=M܇�>�=�u*�r��*S9Ww��7
����Xv�`�r��n�ĳA�ܢ�M�t�7սr{����@z��3�ĸ�U2V�e�U�{z�`B��?�.�����5<�ݸy�d(8��.U�T��?��n�ouń{v{�ˮ�L~r���Ϸe���ȳT�U��j
��z��ϩ��^��s��I��g�bA��T����	I�n��~�F�S�����y��_gɰ��b�]S�.7H�f�
 �-���JKw���&�L�Mff+WS�4�05��{[� z��~��ÿS#�
�D#���b �~ﶶ�=�w����H����-��^pQc]GX��Y��_����=�޹�~t�e*�Yp�z���0rmr.6zLkR�0���� �&�@�[�!�m�����(��THA�M�;�ɾ�a`?k���.������꒦ee�Ҧ�RŒNn����ͷ���p���@�e  ��	T1T�-@��%-	JR�P�JR%	D�"�0�!P�1X)��]�`�����W�g��W���W%QSPX�q�Q�ae�{[Y���z�V���+���4�@ĸ�6��wd�b״����5e�÷���n���v㲙 N�x�4R�mǀ;�z�}�\����j��l}�~�~H���t��%=לSEUF {V�����;ͼ���ý�T�T�ef(XJ����2�~�o$;]CW!��qa
�U���J���%'���ަXn�Q$�,�f�=�SD��"-T-GvI���D�Xw)�}�H�\�ாw�$�$�!Z�&Y]��G�R�T��T���"GB;<�uOSf�g �N�[���ql˒xu��p���q���9�s�:��] �Vz'l�;
�θ������9�c]ʬ��fwFە���p]�:�8�\>w32ݟ{���{~�����֤PIpQ���M��B����z�$u��N(����uٶ{d93�68�����~�t�oz� ��dXg�=C�+y������{\\��Fx�]V+��)��R[����N��krZL}�D{yZ�T��V���ͅ�~Ӟ`f��� n�X{��
eđ9wU���,�>�Xy����T�曹~�}l�L�R���	T�#�K��mGZ��l�w&w�r9B&�� ����}���ENFJ�b|��꓎�g<GƣQ�E(U1T�=�� ��2�3w�ô���];����m�|=5[y����'e��`.S��8J��ͫt���j����Vz�\:�e���� ��uc���}uGn�����3�*���|9�>��n.�k��u�g�ɴ�}a��y ַ6�>��FW�o:����S?H�n�T!�
2��9�7k�D}�;� ��Vۮ�GJ���J�&f�����UH��3w��3˺�3���)9��D�x-"��f�n�V��-g���Aۼ� �Շߣ��:�E�#{�����n�2����vI�p��I߱�n�{�����Md�Ԃ���&J�߾ kn�;����$8���V��(�p�l��$�� �'��uf-�O��:$���)��Ͷwڛc��:�FU4��M��eo �pp�r�D���"}�ͻ$�r4N{��.]ݨ��qV`mՁ���O߿%�m}h��V��,��5�S���O��ͶNy�7j:��n�w��Xo?�PFR��If��]�}�ύs�Uݐ�8 ��9�v�ơA�^`�1(�J����|�����3��y0xѰ�|J>[Ǜ�������o'J�T���.@׮�{j:�=��)g��{Ã4�m�n�v��F��'ٕ�oo<�<��`�z���ҸU�*�6)0�o�7m��1m,�p�85���E?l4����|0{A[$+*k'Wb���Ձ��h=�Qփ����;�u��P��7#�`q�$���S'�D/��,"S-&̑�*�E00��e�n �))�o���&��l�Ǉi��Rq@����s����^��QB��g��\�i��>u�`s�o"C�a���FP{���#�a8�Ie]Z$&��Z���b�{��X�n���rg�[�J�b��E*�Uf �xw�����k�;yТL�z�z��ҤpI)T[�d�T?�p ��Zh�{��'��ͶY���d��Vl�%�۶��h�S�3&�0�F;Z-�r��\�Q�6�DLv�tTݴ�8�:d3�h�7&#7��&ݝ9���ո"v-�ݸ�ڥҜ�n�A��q78�8�+����3�FF�ж!�8:883�6P�oB��jM����Er�iݒ{�6�.�QF�2�L-��ew�ո���zҤN{���Zv����j�0�)*QU_sT�dXj-��p5UJ����<���$�s���n�u��ܥ2�H��g(K"�f{[������r�o0�S��]��H��U6����oU���� �َw&o�r9B&b�Wb�0wT;A�t�Hy�e�g.듼l
�0D�� �S�:�o��vI��`�.���a �����k������ʦ�K��m��ր�����L�Q��Uhx
�۪G���"�BnzΕ
/��X�aNtκcOF�6�J�4�Lp�.ݳ7[�7��I�v�Dt81�s���7U���f7^����}�v�c�DM�Gb{�C$F6�ZC^�
���d�D����D�rf�#=�[P��-4�iԖ���@����sy�=�q��o��J�,�y*adQ�e�~��+m4��f�&��u!�G�ٌ�MR�l!�W<���3���=˺�~Ԅ�N��ʺə���f�w ?�_��9R�Z��/f۫D�H�B��H˂W��is��;�ͻ'}�2v8qө�qGe������u�Fӥ�~���Q@^������gOh�d7J&J�.�B��U�O�n����� �Sy ��� �9v��:	GQ�n�ԑjb����0Ļe��{]C��\Q;�a:b�AnK!2-ډ]����}�@���6�]�!����5�Jb����t���B�qt��%�D����H�&�@���4�����f�Mf�Kh>y�v�Ѿ�����N�����~�rwOg��.�4�I5BSs�k[�,��<��K���2Y>��XT2h�B��UD�r���w/�@��zёѬN��DvjS��ݒy��D߲���0�;ڍ���ц!$���덭�[�p�L"��a�d���2�{	���G �&�ZD��L]��O�T�=�kBrb�)i�N ����T�1��e̷��84��fvZ����=�w�;���=���O�ؽȁ���PXLY��8�s�)C;���� � �~��+
 h��FS" 8�TLt��ohFݐӳ�D�-�Uq�CK�NGc@u��֌��EG]!͔x�#�y���8����!���-�t&�OX�69�N1�ñ�@���h�:�O�Q](�8\,5���Y.Gs؝��=�Só�M���qQ�����+A��9����l�l��̫33*������@$B�H�%�(hK��$DE��E�� DL��7feY������DAրH�35)���&�f���{��Vvx�i�x�]	�9�j�WS�s��d�i�2�<c���l��fB�qv����l��GQ@3u� �Ce�(��.�#���C#�F�3�zN�`$�v��cgi��q�g��n݀��t&B��^�{@�O7+]��w,\$S4�z��c��0R�X`�붣'�;��;vq�4��&�tU�f`j�S�Y���e� Gl�{]���p��v1��E+G;��M�K��ln`	�q��\Nu�=����ۑ�qLgq��S�3-��0�n�;4�=GdQ�{F	�f��J�*Д	�-�N٣d��r�]O"z����K"V/gN�Nm;#�iVA�N�7mV:�zKt��#\':�=+�LR�jK�y&M��ud�ұ��[)�M�ƴB�'SAӀ�ԛ��v��YP+�Yg����OYi�Jt���Dy�k��-ܤ���6n�&��hJ���XGl͓u�L,ru�)ݺ���<5�u�G��n�x6��L����������u�D�x���=D�"�� �lT���v9��9� ืrN�$��ѷ�tӍƣM���H�隣�1㢒>�uX��A�S,���ؕR�^��(�eYi]�sm2C4��HRrDTbM��ڞͶ:��F�
s�7�7-�<�:������G���[�bם���mMB	)TTՠoy���w!�uu�;����G�AM��vj][5P���;쌰9y��yw\�>�x��Ú���J��$��7݃)o2�N�n��cw&��fy��yy��g-R��y-n���us��L��1ޜ�J�+����y7o����k�צ�we�#�Zwl�	�ێ6��W��"�e�Ƀ*�W]u�l�R��\kAE�1s����q�v��ϜsY*��B��p-�u�7��4��9�2Ǟ7%ۖ����l�]�B��;�' ����8��n����q�d��I��*d����D�*˸�.�d����ˎ�����Nbj&�&���c��v�7�:����+C!�)��wˢ	T�f���8�12PHH�EJ��ߦ�!�u;@gvO��}�}l�����HJ��D�N�����l�]�!���H{z�a���K�0�&k%D�
�{�2�׭��c6�6�唈��:��"��a�cz�d�}L�9{���o~���A�q5�Um�P��{�h�(>���n�9G���GN�G:�@܄6bL��'/s�q���D��fݒ=���rJ4� �A��H*���C�=;�@�U��g�Ɔ���-�ٓH7)���U�YG�l>݀.��rfE������G��0��ͭ{{�����K����"��6!HF�.t�康��^�)�u7�~���7_�^��>Ue�U&2�V����y!�:�h3]2�3zz(&)�ݨ&�%���<��Kj�ź��r���=Ԅ�rELeMܥ
�`�L�5x�r��6{i�g٥3��!�Ѧm*mS&�f�$���~"�a���\��>�� $iEr@��GwsN�}�E�p<皰��!ĵ(���2�Z)B� ����>��x�c�����N-=o0�}�w�A-;�<������Nr�8��}��n�> 8� p1�H��n�'�醉7�j�����ITd�b�d⤳vy���| KW�m"}�}��>9��)ʠ�L�MI
���]�b�����MZ��6�V��9/�)[���t��٦�v��a���;l�����:�s�2NIn%��n�'�y��7�㔎{�{fFMRq���E*�b�8"�Zm��j��'�g�]��n���Lk���+��bu1S���Ⱛ*��1��1�q`VovFrf۵�;�7�6n6"à��<��Q�w�{��\��b ���*�fu�`��,5���U*���̊X$���l�n�=���=��O���W�+�	�QSU�"�EM�i���z�����xȱd-����E$�-�l�M{|7u�KwhQ$�y�#ޏn��q�]�R��I$�q�Q4�RD��B�n�
$͘�^7���o0#�Қ��SR]U䆙7�uWÜ $}�uQ'�}��w�n�7�Ǳ���MX�C�����x�u���ڇ���GJ��*2���2��n��=���7���9Z|E(d��� ��A ���Ī8!�#�/������4
�BQn9/�aL6�9栮o�>�~��Xks�ޚ��H��ثnk��Y��d� $5�qr�Z���շNR�v��i�J�&�tu�f��\N����;�$�3��3��C9��u�b�쵳�Z�fk�TW߿����W~x��B$�v�v�V7vOu��d�����S�r���s�t��2D(�J��*�Y��4uo\����G|50tHJ���) &A�1"b#m$p5!��I�}�&׏u�gsy�{f9ܙ��H��U��%y,��Ձ�i���n��{k�,;ML�"���t�
��a�� o�Ő��;A�uu��CR:T��g	�wJ����]?�����\�t�.����31�Ȝ��>RA*��~�}�e/������ɓ�w�������N��7_�������D�he�s0o,#!��s�T�>�Y[%�7�evU�-]��0񵓆�E��Ѥ��Z�ϑ�,pX��WA���)I����R�.�}[��㻽��o{����0㞌�	F $ ��5
��t�|����jZ��������J&*&ɻP]E#�7 ަ�a)���w��X{z��#��SSy+2js]��Yin�����\X�M�ؤ�.dtU�T�TO��)�|~��>�6�|���Թ�w'oA����p�˚ʎ*�I�ehRH�k�����]ۇ�լpֻg�A-��J���{!������a�A0��J�}9~*2І�]v��rU�)U���o$<�s`bcqr��D?w!5J��ɚ EͪK0�n�x�R��P�G�_{��*��̔I��n�;�N�J�U#Q4P�=�X]�:�o�Sy!�����oTn8�\7q@����s�^Ϩ}H��f sM܇n���=0���QsA��Ow�v�? 89��d4�+���m�����%�o=nz�pA3H�����T��L�5n��dzN�#
;�VlZ2��i#.D ��fMB��WeU�yw9�11���uG{$�y��*J�Q36�K�bn&�ݮ,<��C�[����Y��JbZRл�Qf��ཚ�o�7w�G8�iҀ��@�]s:��$<�saА���E�u3%�TR�@���@6�U���������n���6c��*�Q���9�i��\�`.ˮn��V��h�Pݻ�#|(&�!.��3'���7�7m�����t�أ��/��q5rĔl�	$M�ԂS'�{���mC�_[�kuaܺg�\���˺˙�Sr+����o<�;z��zc]\CمSQ�$�Ԇ6�tI�ɻl�-9܁���3�Qև�N\ �SY9J�I������;v��[�r_���-�����X樴�Q3E�������f��ta��3���v���ʇ�:�.J'�S�e�aG=e��u�������
:�ָ�dV&:�ۉ��*:��՗WCtq�A.y�a�] 1�ƙ�ՠ��uZ�%ҽ��[v��u' X]� S��m�v6����9��'��� �����*�t�0\	H�ޯm2V݋e�`f4���(��:8�+���i���kr���o$������FL"a_~�#�&��"\��7f7]��l�UUA$�ިv����@v�Vn�u�OF(R¢�m](B���o���o�-�4�$��2�&��+��ps�/�Gɟ���ݗVػ��$��禍o۲��mq`=}o�$��E*���B
�j��^��I9�L��3n��s����ŇwG߾�U�K�����=���[)�\�>�;c�鴚��%�mS��i��O�$�����'dd��<�����5j�v��C������?�1�UEUs������?�
�*�C���5]�p���!B�!DT�E�����P�@7� H��" �� "kX��u��D�PD�B�G���]o-  	��� ����B"�� u��
�2��(�2�����{��L�޿����B�EUJ����Y�o�~����{�������������]���g?��8?��?G��7�_�����������TUW����A��o�����
����QUX����_�G������=���C�����B**���?��?��:�y����A]G�?��������lr�?�'����� T�(R
D��J�
A �@)�J�
�)! �� ��J��B�
J
B� �"J��
H� ��$��
B� �ʉ
Bʉ+ ����ʉ*$�
@�
L����$����� �+*$ 
B+ ���$�$�����0
B � ��*$�*�(�) �B�� $�$**BJ		$�
���@�(B�	��		"��!��(H��H@))
�	 $���B�	
�)��$�	 BJ�H@��CBHD	 BJ�(BB�B(BJ �"$��� �� @������$�	!2���) @�!
$!(�!*H! B2�!(H�� �!(H�! �H���!! K@@�BH KA P��� J0���,!,(����) H H�B2",��J��0 @���$(�) J�,��B�����
�
H3	�a!��0)� �#!J0+Ƞ #��@�# �BB0B0���!BH0���!� �@��!ʄ#0��2����J0�$0�B1���S[O����� Uh�/�?�?���У�!��?���y���*�����������x����������TUW�O��C�O��������� UU�z**��i��?�o�������5�
���������FӠ���a�k��f��C�ت*�uw�A�W����*����h����g�o�8u�O�2��#���*���g�o���UU����������t�z�����]���?������~}�����t*����G�g�#�M�_��O8�o��������_���"�������O�z⠨�����������������]���_���b��L��<�}Z�J� � ������!������Q�C���4�Z���>     ��   K�U�7���:�A}�/ x9�Wl�r:i�եM�gU�ݼwl��ZhJځ�:�� 4N�U�3���RK�x �z�`�K֪�&[2�,�;p=��w�N��2@.��j����g9��)$�5�@��ӏ/�x��Uq}�s5�>� �：ٹR��+��s:��|���}�/M��scvS�+����]i%i�hsu�
P@ �@DUO�R�I��ѓ 2 4�� 4�	%ISL�40&4�F�D�*��)�14 �A�0(Д�CC@�Ѡ�ё��4�%$#I)�i�z����<���@ ��BM4&�T��h���d���i�By�	z{>�w�V  �����/�U���({ޅ���U�O�W�����ޢ����������?������+=�_������?�����~�^���3���ϟ>]N6��Ϩ��R��zv��`5�z<���6��!��z�ajHw��<�x��K�x�b#� ���f	"��?f����_�o�?�	�}�=���I�$[!l��V�-�6Il)��h�ڐڄ��l%�(�)�E�I��d��F�M�RM��HlR؉��� H
�	�8[�Rt}m��<���C�΍�T���n����V����uz��3��"���ܻ��.,��z�?��MSV�H�W�J!Av�©n�q��l��qNQ�6�t�TH�*K(�j6eb��"d���u�e�P1p���QE�("��ZA��-�u���D::�"I
-�z�g\����SLH@� +D��*����KKa]��U9x��_<X(�ld����P*
���x�T��NYo4�ܞށ	�8L�W!7:�c���Azq�۽Ѡ��4���Hd@�ꭝs�L�ǧ�Y\4j5g�ӛ�\�1��g���m	�q��H4e��T�f���YD�`A����F]���G	+���h�2F��A��A��=b�n�^�S�1Ûɢp��	4Ņ�(�!`��eV�E��gE�)��_^��@��G�z�``���,Z��I��B�Ü�(J5�o���Lb�.��������n�p��4cl��zR�%5B^BYlp������ `J9Q�%Ʋb��Dz����G�	X7�)�7�zN��I���$�ӗe���c3ZA�Z��X��U�d�N:��^�����e_	g��
b^`*�I� PD��ixa���jh�P�J%�%p8V3��1�T�GF͐�������d�)�ǹ��� �	׎��
��� �	̹wف����j��5Nx�x�.�*َ�y�/]L۞����!ԃr�+�tf�ƛi�5q�Ȥ
BB��c1$���OR���)`L PA�F1��!EF�3����t���%�M�l �5ˬl�/&I[�r�B)E<�D�22ejY���D��26 "����"��׮��1��a�9YM�x7��t7`�e��âU��*텴J+A�}=Ntp`��n D$B\�&�i�y������.پ᣼(����>k�!Emu���l�ۣO�+�$Լh��0±��ǉ�H:�8^=s�����vE�#�=��@�����[a=h0����у�k�:ƶ\*��``�t�(e����k'.�l�իj鶜��H6$LD)"l�����7V�m i9l�n�uH<���!D!��E�؀Xͮ��Mh�X�˜���IPr�Z3��P!Kx�g0IZ�]�DPJB��A�:���բm?#|�6���5�k�i�>�P?o��j��G�i���nN~X^<(�oi�.g0߻���>��,�{HOq�gx޳�o'��@�q��zbU���]]�$�Y�L@6@�|bk������&��t��e,�&�_>[����h�!�x�r��eE��r��tˊ�j]��	C���t:�Gws���t:�C��-�I-�@�t$��	����t:�C���t:��$��':#��t6�nI$�O��:�C���t:�C���t:�C���t:�C���t:�C���t:��$�mC���t:�C���t:�C���t:�C���t:�C���t:�C��-�I-�7Ͷ�C���t:�C���t:�p�b��$�� tr\�A��t:l0�t:�C�����@�t:�C���t:�C���t:�C���t:�d��$�����t:�C���t:�C���t:�C���t:���a��t:�C���8I!��t:��|g�|/���C���t:$�� � =S�X!��6�^�03��k��^�(�%��4C&�C
"Ģ@�t:�a��$���v�I
�vBIG�a1 =ʋ���BzH$}����=F���t�:2�,s����vKl�Vl���3��%�l��'5���wb�|/�����E�+�.�W����l�$�C��ߠ,����,&h�P�)��;��d��&
&�N�a����~� ��Դ�vw�a�}o�z>w��\���ݧmu���t:+~�ҽ���y�֮nޔ>��?;�q�$����!w�\[AV5D�,dʵk���Jl�f�/ݘ��M���7ӻd\����X����r�[ز�`��������R�!>a>PD$���鞾����t��3�0�,�O �t�m���	$�U�{� +wR�v��}z�:�$����%���5�kxe0H'+RԒw�
a|�h��3tf㙽&�n�޺�#��������Gf��@Nm}��8���+M��g���6�Yt�9f���F�V���u�O0q��=c��!.�]����;Ǡ���S���XФ�3
�r[Ow��t/��FM����Ja�C��ݹ���.mco$1t��_�� �{�nw�Q�Uی���w��� H�I�ovr��:$u�5�n�a#�C��& ������Gt�J~Oŋ�kK�V$���z�r��!�zVWP�^�t�����A�p/'Nl<9��;���:��]⧮�/|O$`6�n����6��ozx�]NY�{�q��8������FN��C5��O�{��'wtȎ�:��nbp���on-�&��������"�ɿ%����n�I�$G�UM�jwY�1֖��4'/r�bD�w2%pn���>���  ��t:�$��#���"��K��/�r�D�`��7$S�@��9�f��Iͨ(l������B�I˷pqz��!ht�t��7��jn��e4�&�����-�C{f� �ۗ��V��dIgK�u�{�'�;���b<P�(d�HF<=��륩���~�o����-sz���=��^�PS�3wzo)
��b�|z�,�N��N�=-f��8ٌ^l(�v�62�`���2|o=���!���Ҹ�I��4���c�v��(ʠ 6�C����-��Imd�����t:4ȠP����t*-�C�l0�t;��X��(t:�|���t6��O�V� v�Qhtv���b�Rӌ�a�x6� ܲh�귻�Qht5�t����F�5�vz���שu�*���d8i�_�XR��,��rU�� y*�.��S�Ը+�=��H���*zĂ���
�2����]�P���%寲�3/f�{9�g��0�b��"f$�1�]LCA�N+���j�@zk�{4�{�6�����S|��ޱ	�zH�5�֭��w��-�Sq�7�׾��Y�qq��浛�Ř�c��B-��st{�Ӵ�V*���<J.�ԯW���}�Wy�ܪ����������PUW��p`E>�2�����u��������!� S��#���~���_�������/�l�i�}�Pt":R�ċ�xD�;����Tv!ái��xc�$bd2ץ��K�"�K@�"DRi�#(�*E:ȇAhp�)�ֆ��@1�"p(Aoh	�2�r��+%�pt�S�Zq�X^΃�x0�"���Ev�Y6F��"��w��U	C(Ț˴Cj������!ҏ�7�u^��u8X�;$ �U0 H�S�ۅL"�*�Q�d�Ma:3��8��±P�x�"��tpH�2(<4Xtt��{��Iֵ�m�t���b� �'���U�P�똬�*VLo�@SN$cL���Hb�UYF���mU+�@s6��X�+&�P��ڳN����Ҝ����M�.��
��x6Q���S����e���Y�x�Vfvrkq�I%���d�Ln'�Y�,qil�p�Ĭd��s2�m� х�p��Bd�l��0+�&��r�Ϋ��럃��خ0�γv)��m��}��\#d0�F��k�$��?���������9�6�#c��3V���z#HY���z����2�%H����wذMi�M��}~��y�_��uT
]ﻉ�5����F��n�mvB���ԗy���Ғ��3v�q�E�b�v����~�$��vf}>�	�PuU^����s���X�<�����(��j6Rx�u޲֔M�Co6m�d'U����Xk6gݗ��+��{� �xbV�mH} ���.��7����v�.(�fJ�	�K�H���,,޻�3����:~4��F���lA�i<3�;Ϲ3o����\�������]Ȼ�M�]^i"�7R{:E�7}���2�R�	�:Y�N��rVܩPN
��J14ܹ��#N�'�~f}�3۸��~��	��"���y�Z�6���̹�� �!T$ݽ����c�"��h�$��A�#�k{~Ƶ2f�Ff�W��Ƿ/�p�t���ȑq��x�f��-C%[�ݻ�=��37`�٪�
&�y��kHgOH��ZG���,"�mBT�@����n��B+M
B 7� �о�X��&*�,���qkukH�	��w��ʡ�k���n�ڐ6�h)�>�j���r]�Kh�!�p��Rh��x�U�Cúi#͔�M~�!��/.��l6�-�@�CMa�ߐ1�0֑f��-m�CMY@��Ļɸ�Pq����Z���mH8����v�6��!T�X������]p)�0�C-�#@�F谽������I$.Yh��Q���fb�Q��B��b�_"YD6k5#��|�hx�P��Gh{~ՈZ�c/�}�XAB`;�G�L�lamjq�ݍ5i��>�[�bΛ�UN�$�0��q?)�1��������UB4�5���7@�=�chȂm)4D�4��f�BKE2��5������61 ��/��#�H��O�W�u�CQ��g*��q�M<OOw�p��R���:j0�dX�ƋB�IZ�}Q�����5���,�	��`B����4Bb�Ĥ� (+&�@j0���B �)��d��rT��)���2�D�3�b�l�}�(n��]b�����""" �����D�R[�_>�"".d�""�9؅��v��.�d+@�Gf8+�q����{r7`٦���g������6��bv �5���� g��'u�VIZ�>�뗭OZ��C�j���*8��=לM��A������h|��>�N��\ՓZݍ#��X�$�}A���J |��R�6�ÈU�Sj��=��B�����9��[���4����>�?�u�{� �'��r"��Y�q���f4l�I�%��CO��3��"�Gr֑f��^�K����5-���x�@�@�C���Bڎ5.H�����
�X�N}X��9 �����V���������lLx�7�T��jCs�2><Fm��F�e�Rho!���5���e�\E�����{��q�P�hi�s��+��
��a������U *O���)+�Cs@y}�����U��+�NZ��uߟ���
}F��뢯�H�F�����
M�����;��{������7�����@q!�q�>���Wr�#H�_}���w��~�U���hJm�^�"��^q�X��,�eH���X{�q_m��)�8����h�z�wD�gn�a��|��3��m-Xǈ$�!�8��o��|#�3�/�}$E8؉30x���5�P`�d����*�8�ߎ�r�j�5�7�;���;�ǩ��hI �]*#�8�܏�f?P 
>";���	���E�G�x4�p��'��?R���"��i��r�F��0�Kk���0׍lY@b����D<i���C�?\����8�o�p4���e����?�na�q��h.��Q-�[��Ny��.�����>�fF������~��a�P7�ڈ�������i@�kia�x�#��_62��ɸ�!�7��`����v��I�}B�C���`Y�1T8�D}C��}?%v<k���FR)OY �;�ݾ�݇j�L�����p������N��w~^�q9>S�U��,�"��Q�����^?�!���#��r��w!ը#�a�ߵ�yn�����j%<� ���:�V�bI[���*��뉈:�L.L��hq�������B����ܡ�pV�S�"�d�����%��O%u�u~/�V�S����w�2��`��v���ִ1uu�"�/�n4�� ��! =۬#ƻ����c!"�E߀�����^��k>`C�g����N�u~��KG����ƿ2*��3D E��1���FZ��MC��'g�آ*����~mi�E#�(��gP�G�����ErM�Ix8�"�W�~;������ʲ�����LqZڣư�lo�]h	��Σ�a���TB
0�G�����R�Ϥ6��sk�`�s���H�J�Xa'1�Z(�̊�\*�|v�b۴���6��ah���2����rl
M@	!�8�5��T<���r�9W�fz���e4���J�߽��F���w�b���X�Ы�n���08��v��C���4y��ͷ��`�"�~7Ghux���z���y�i`�=��FB�ȁꐆ�uǪу"N��Z$$�SW�XQP�~Sݫs�i����2�͍[TQ#h�` �	M�0;�0��[%02BF�. \/8���R٠�T��#ABL��%!`���M7�Ÿ�0E5"p�ےImUU�f5r�h�A�Wk��+�v��`��,\gb��l����+v�k�2�Ph��K���Yt�ݵ�Vݧ�\��+��lV�H��M��m&�)8BP(O���z��	�oa(4��p'p��JN~"���H$���n���V퍋B�؅K���+��������w��������Ѻ/@z�� �ʝ㞨�G�@~\C���)v�󄒱!�?2'���b<�`~����[Ʀ�n�H�0���Q�t"@],�c��4���5H� $��� ����[d	�h�#��H�>�#! F��I���$�sX\^%fT���x��R�
A$M���	��$D�J�H�9BT�]�ԓ.�f\�H���;�IQ:z3qw��ba���2b�z�D��K�6�2捓�9�mNN�\�F1c*�_\�ˬU!56<�̛]x�4l��a�!*&9Cq	�R�-�ݘ�߬�YMA$ؤR,@�@J'2s&��x�Y6O<�m�`@�"�D�A${��o����$H�.�"$$�~[q���J �O]P�) b%E$r���k��bn��q��1���Q	�r�F��jm���SPu� kt������8��	"rD_��R��I|��$�uT$�c���FMD���M�BH$����@'|�!���qB:1��L�آ��f�4M�2u�Y=��m.�*)!����jbĐ| �����&ɷ�ɴ�2la�1ٛ�����	|�)"�KJ,�d�:�H%�)"&��\HH,d�A��I#ˠDD���!�I�R	"u7ED$ME*/nڼIsx�0�H&�I�3�K�H&ꄐIQ**2<�=���n��$���\A:�RG�
���M�!"�﫮d�MX��BM�jr	Q	q*)"�=�{������K�i8�bUP��|�ۣu��z5�lj*�\��x,���b�4���o����W[�V��6��H��Q	�ߙ��_{(��E�С���)"&f�\A;�) �5�0pfg7
����MA$nP�	"bjY6M�uU�e�M����HuY-j���b) o�� �J�빓d�y˚6O<��m^���D�ߗ��f)"�RE$D�$�I��$D��K�H�����q.Ԩ�H��PI��$�H=n���(�I �3��d�K�PI�i$���n�%�� �F"�!�P�)"n%A$w��9Y5b���p|���BvM�@��n�+�v�k��q/E��}{�n�"u�K�H$��TD�P�$�N��߾��J�&���BA9T�"&"TRD7E	"����$�;�V�&1ް��H;�Q	��J�u��%���	9��ްf%����3��P�	"u�K�H&ꄑD�J�H���X\e�\ $HH. "$L�o��[`p��c.�PI�.A$�J��o}I�Q3&u*QUF�����MЕ�:�PI�T�	 �t7��k���Z��7�A���j�BA$M͐.	 �U	�b �}و=��k!�$�Br!PIY�����r�Pn) u��=����K�Y�$D�(n!"��RD$MĨ��������|9����#H�#��B@�����4�𘫺��S�^�3BA!�R�&� \RC�\�Y\Oe�2����2!p[O:s&�ێ&��z���emb	"�U	 ��Ჲj&"TA<���G��f�M]jly޸�"A;J�H$��5��{񬭓6JB��'Sp.	"��BGZ�r<O!�-�4��O9sF�����\�ļW�ΰ�O�VƆCS�ۉ�6<i̛'��A �&�h���%/U�c*f	 � �! r~~C<�v�Uw�d&�o:9����'Y6O<�H��1�u���._:A"D�3���	�(I�5�K9CW���]�I����B#|�C��E��(��?9��Ǒ�@kLj��㒿�	�X��@I-Ƀr%�ݲK��S�W�����.'��5Ѹ*�]�W=�� H�'�3z��j�u���%�!�:kH��D�3S��
ݎ�ZGu ��-��E� "8��`P�����Z=F�γ��~���=��,#��@�u܇��"`�#F*��j�ix�`�����$��pI����'͂��7}ξI�����#P����c�>c�U{0;��/�I^4�a�#߭��������/�>��Ռup"�_}<�YD.T�w ��B8�("U]�#���,��d����`�B�4�C$��c]c��i}�@��<��uG�~�zz��OY�x�V������G�Ǽ��v
��W��x��8`��E�dKP	���0������|%i!�*�f����!�RC ������ef��Jٻ�*B�iTÌӻ�f�M9]id���r2���D��c�����vb�LPOEBɎ��d�����"""0�DJ���DD@%�U���z{Ur <�SV���>�g��Gd��g��lUg�]�'��5[[tǶ��m��$�m����5�A�ϭ���>��vl9�/\y�t�u��l�]qͨ�n���^�OZ"5�E�hDMAn6M��*��#e�ۡm��������4؈� �݇�쮁�4�]�0Dt�)9�+�9�{N��^�5�G����_���J)~M�!� ��F�o�ĂIB?>N�α�{������v��#Hk�9i}���y#�f��~&:��1�
�k�@+������L�f�{el���^f3#)�ub�c���,uF�T���HHEakP��~Q `L2a�Y�GƳ#\8�[m� d��d"Z���꣄�Z}'Õ�����x��J21���\ �_}��ۻ� ��jL1�A=���=�Y�*�_����*�7k���=L�P�U�� ��g|L��<@b��!=��G� ����7B����q7�d}��@b�5�����t���	�$1�.z+QP�Q[��	X�f^F�D@��`i�VG�k	\�����Z4��M6�%��ǦtG ?v�QH8��׍��g���L��:@w�b���41����ߛ�N&���a��]h�?���i�E��:�?fn��UF!�ԶC�}$j��@
�B����=| <k1�#�5==[��|����'�P��v��h�D�k�A�2���9\C f�g��"ؤ�4�GHi@����s�b<Q:�.��Sk.zAz��g=Vn %��]��̑���c��j$�M�H<����]����6����8Α�1�]nV̐�1��>��r�G���� �m�YQ�Xk�i}�Y˻�Y@�A���<�!�Q�zƥ,W�ߑ�~I�������U�p �uv�����Dde8Ll�\H	|㳵f�*�,Տ�nk4��i�?o�4\hNUf����	�%⸆��?8ľʾ��"�����H�{6*>Cc��1f�UY�5����wc�
` 
@���G�,��*V�#P�?޳���<0Z#��ip�~W�0Z�-�|�L�qH���ʲ��q���q��m��!��	���C�Q��G�����f"�% .�Da�B��a�"�W��|��k|Po�&�E2�g����C"[�R$��pi���La}�� ��4՞��K�hij��t:>��8�IzĀ���5�P���2պ�nn��s��W%����-�mfl(~\C��߾����(�O@���C�7�ߕ���L)[� H��XG�~�����\@���9wcMC�/Phd������α�:��n�mT!�k��0��'V�>ب��c����Ȳ���p.Ã�cMɳ��2P���L1T6����ۈ�dƵU�UU�V��ڪWf��H͆VѻiX0��jim�N�������{rlnP�>�V�b�-�޵=n[U��+���s�: �V�lZz����GQ��[w��8���� �	 ��1ӷ\
G\iD�V4ZNݑk�+���w���1�p�A�߂k����Q5D��x�	Ԃ=GK�.����QG��vy��m���C���H��5)>ʆ����de�a_��w��Y@�C<����R�87�(��0�	(G3j�l4,�ýwG��i�j�W�8`�kMd\x����#w!�t�u�Y�U8�>0�h.�#nx�5�U��H�%bM�%i@��a�)�W�(��\F���aM�0���{dX�FBG�#��7Z��������oގ�1�p�6��W�X�hi��|(
�wtIe�s-�Ƭ�i�͚��ZB5dz���i:@�A��"������t*������n*�l��n�eXP֩N�c�yk��c�m�ՆY� ����2c�G��ӨQ`�*�[̃h��ʣ� �� ���� 1y��U5nV����Z�+э!�CH��wf��*���`��H�(ק�����}�jG\��<!0��XԒ�tI*T �u��U�B�� B8��A"� �4����'߃�#�Y��,�����@X�4�CRDf��4��(�}�5�m��^_'�XE0�`��Y<�j܍$fALi����pZ
�i�wTP@�Hi�F??"5kHz���4�i��^8mzA����m��,E�"����I�-���C��Oz��c1����#����-1��W �Y�h��*�%�����N6x�#�畴x�#Q��[]�6-�A�w�C6Zh8������!W�-��6��a�������!���1t�Z��h�:C���go����q��iP�+�m�j8�%�#/m-�fa�Sg�3�g��Hi��H�X�����w����L5�����&�P�����j�b�T5U����:@|A%cߔ~��5Y�B=q��vlR�0�#Gy���B 1���M�:�#�.����$�I�V��DeU5pĘL��!�'����s��J��=���a�i����.�� ibkH����5kM_�)0]a�x�>�BT�#�<���QH���q!���$ٰ�J
mV���$U��@�4�eș�#Uv�H��S�<Eo!�=�F��A�|��	��hYs6*8�LzaL#$����L�4:��6�đ�z�;m�b#��Bd���W�_g ]�Zg#@D5ڨ�h��R	�=͍X6B$2�!�,E0��Z�җaNU�$P$���,.J �]���v�*�e^!
!E@���m��U�]���ZX(�	�Bl0M����n�nS.0�S��6�"""" ����-$]9��"" ����U"6�kt��HI�U�z�j�0�E�\���kŵ��v��ki��òάCnخ\����&{(���f��s�l�px�g�d����qSi��a;tu�p�\"�6��&�inx�Q-�ٙq��6.S�i�ϟ�H�y.��.��ƽF�{�싦���iK8��;;2(��::��kU�����Ȳ)D��/*=�f�W���m�u3)��qD��-��!�ec�\���@Dg��Ǧ����P篅��G#�෨bnK"d�v^F���J�����p�c/g̴L9R��jے�W��1��%�0�'����r4%����V��\f��Ƴ�VG{�dD�uS#M���Ӭm����;T`b���֥�F�`&�-K���I |I	��x*�d9��+s�ѻ[<EPt
#��Иi`����1b�~� �?��<D{F����jm���Z܇;�<F؝��a��tG"d������x��L��e�"u��G����� �ы ��At4��w>��@��{ڛ�r�����=���-�8/�� �*������.�JCN5� ��}�{�$#���q���f��v�[$��j�/zTs��"vMuj�v�S�뭪㮄ؘ�f��wUC
l��Ef�0���ڬ"��0CY��֚�ɉ��"��@����k�WlJ
۶� H
P��p��S�$l��" KPȁ@R�����H^�h�li�w�"E#��Ha�4�`�ځ�� F����ܩ��
�-m�	Df������� l��!��
��}E0K0�LN��5�gR�Һ4�
��U-�(�(�=hv4���'?ē0�մ@�����O�����yp�������ԓ�dS��=��%�C�$,���0Z}@��V�dy��2 3P��(��i�d0��Vh<�i#��l��a�j��#�vz(4�5�ArG��7�
M5{�ҋCuU���[^e[k|��������R�ݐFch��9��}���66�^E%�Wk��E�Ø�%*�@���CoU{ZZF Lq^u�����1���$l���8�,+�e5i�(3b�CB7��f��5Ɓ���Ѵv��c��S�C��N"O�ib���<��	��G��iZ��J.V{s�S���(�+0ŵywb�O����Q��U^�G�o2iU�����C�b#�C��X�<�*�3��д�Y�B<�����4֑�+�l���i���J�f/Zo�:�I��2q�x\di�*�Hk@D��SP� Vp�)���P��H���mM���t���.��k2KN;�m-8�n7�6�#�a�� L���	TB�G��7U�~{����@j��2(�V�UYF�5r�mU��l�&��M��	]�nwnby:ۇ#���\f�кr�1�k�w8�����<�͚���093�c�*�Pۂ
�U��j�Đp @�P�"lզ̦)�ޱ�kF�]�����қY��"���2��ٮ� R"��mAu�Y�w�	r���B�~����V�����=�C\hz�D>r"�]��d7�eLP���ΐ�9���V
�tr��Yfa۶/��������4CVE�>��Y�Cdi��׆ݠ�j�4<@%kl{�-���Pu�C_1C�H#�m>/7v��)4�pQ�3UYB��Pv�MJ���t�`c��Ǘ��6�\@�������MR+���J�)6���g��AD����t�j��*/��L���� �C�x�g���N��c���&!�k'���������:Ф�f)��
��4�Z}<�Q�iN��R�KRl��׻���}�,�ܥY�~D�>B8�a�'��3C/6Ż2�($����H��{>�ZF�١��������K	�ZB��C5p�#�^Ϛ�˶,o*�M4RC��l�'A^�,�lP"Si@�B@Qq�-�zv�s��qk���|��O*�q�"�P��p���hf���
�3�C#�	����2D>r:D"�!	垉֑�����R	#R��̚
d��������h/7 �
PIT��<nrz��t�n%��q<�m��tl��ߟ���>�wB�[~k;5����2Cn4�1ߓ�GBjq ��۰�r��͓/��4���M����߉�i3{~�&Ew��sw�<<7��ъ����o)�hK,�߀ }���1�ߞ'_��1�ɗ�s�\�ϻ�����~0,��Yl��J�v������.�N���L����-3t(*]�Pf�%y�����/q�����L�p������of]��dK��͖��`�|�����	S���Fn[�v!E�V0#�p�WcNx�q�\H�.Ȇw�g��"�r�>�o؁�ϥ�k��6n��y��h��4�M��6�MM�Y�7-w���OD�	 �C�,���#�����ۅ���oՙ�9�({;�q|�@���{��-]T�m��>�ٿ?�ikVl���frk���d��P4�1h�$�9�,/BY�h{dd�s�'q���bֺ�Ƶ뮝�m�۷�&�v�b�DPD�� 	�""" �����!�U�����""&H""]��E&ݗ+ ��Nmqu��k��m�U/6��]��p���E�Gg��_Y�=l���z2v�ʆ�رmƺ��lr�r�i:��he�\ ���\FsQ
ci��5u�ݨλ!ά:p:�	8.)#��]\Ok���H���hۑ,��W)���:擀�!I�	�\+e皮��;�s�rv���< ~�~Ih1b�+<_�������ٻ�6^8{�Ʀ�]��9�ھ��ͽ>^�ͧ����k�"v��Bع�G[��ȒX%#�:Eۚ8>��;%�Tߨw���lȑm�5/{�%$�:2m��_�ћ�7���둶['��?M��u��{9f�n���vd��۽:�B6��$]��-�B�v�N�:1�A�{�ߟ����iy7{|~�*5|w��	#f��͇y^�r|E�<�.����{{G��縳5(�Yc77��~���O��xAs:'��\z���d��xG�}��h=5��0�2��A:�hM.wS0-�$���՛�����}�Ⱦ�w8H�����ֈ� B}~�,~ ��ΕW�|8gC��Z?4��
fr{������%�#س~�^��������س�Ж-��^Ȣɼ�@�( �@��	 �*�@aBr��7�w�L�\�j�[z^�wS"rv+m�G&us j��lc�!��Kv�͑�����&ԁ6����Y�4H`��͓nw���vnݾ�����g�!����*�/�ှ�_&�mD�f"��;76�N�4�'�6͓��љs�gD0s�
	S�7f��w/A�vo�y�5�&m�jd�gWۣ�=�w�����|�n�쉤����n��6��e ݷ���6k��f����os~h�֍>�FR��
�4�L�˽D"�M�����'���M�/�lk7T��*H�"@"�ؽ3<�ў�:y��hÍ��<��%G�;Vx�m�L��)�w]����83f��~�Y���\���C�@bD"� �۷������~:�
L���y�.���s2�B�G-�w-b&3#2Q�#�;2Z�7}ȶ�D/�h�����ot���A0�nM��w�}����=<z���L���ɢ�O�Ʈ������D��"p$S��v�&|���Q�DK�+�U���akڒ$3۰��9CI�I*��Y4�l����7:j��f���Y��b&2�]����ѩĪ�U�UV17T�[UJ�խ؝n�������a:1����]7k���7k�n�E�ُs=������|�����P��&FV�B����J��/v�v�{�F�D��`����@{=zB'���@c��+nȘ�!mv���d�C]Y����hyￏ���+l$���}��>X�=����snm�<^������{�ܺ�I ��dIⷞ��-�I��>�w���l7�����{��݊�9΁��/<�z��_���/���_�RM�}ka�˅�-槷��Ĭy��׉��~����d�@&D@$P�h�ɩc1e����v�㸳m��7F��m�sF��?"��g����a3AӬܛ��=̇ߦ���]�kc͵��ۛ����1�x�I��b%��ۨ��*���H��q��50➃p���9���۷rM�#�1JL*qͷ���O��߃۰H������Z�}��?~G���${�����V��ɖ�k��mg�M�zÊ�d�	E&Zq�!k�&�S�I��ʈڷ�������O8K0���=�(����pgy� �^�=\��轥XC��>�ь�Ҙe�췛ono���@�uZN߽�����Uo^{�|��3s��:���T���&�1Dh����y�(B���Rf�������}�oڢ�DH]�ɿ[,�ۻ�Xpn�y���	#e���{���&8D�[y��>�Ml{�}�z��Sw��nG�[�up���|\R;��pE�[�LcN�9�e�XzEFאmx����f�c��x��:e�Z�mμ5/�"Y6k�޳���^nެ��n$k�r��Huf��<�Ǻ{Ο�!H��&k��'p�,�rH�p��!�%V���Ó�����n�v{�$L��Q��iUK�����Ϋݿ�/=�Ox?&KnHӨ���D��N$nF�^����$v� ��*n	�/��ؘͩ�w'.���|\��2z��{�hK�vf����7&-��ڌ9�:��2(PU<Σ���0��e��:��QʕP�db�2$�8^ �K�����N]Hń��rƮ���驄���;N��H�:v�E�b�Sy��cVb!1!�0~z�⛪TRP�MKvX�5 $DDDm	ɴDD@2t�9��k�� ;gnU�H�4�1��n{oF����q�[Jj�\�6�V�z�tWh�L�uݭۭK��!�T��\EE�lc;q;e���Oa*�+s���b{Q�������L���+@@��sѪ�z^{;�{=VhUZ�r������@(�#��u��.�A5�"R6l�'�]�a��7�����I}����$
H"J �,ݛzTA�I�����sw\[�[mf͗o��ѷ����U'�<)�e��I�v�=��sb$��Wi5'iڠg�k��YED2��kB�4�xs��r��~�|�f�~�EDF��y�v��vD��`�3o�&��\/��*�{_�zQKͤ[����� ��Ϳ|#��}y��{:RѮqQ%"F����%���v}�.)��/�������`�=�mݛ��$bj(
Bc�fe�B�m�:����^r3��U@^���Mg6O�L��g����������xv{=���3���oi�� d#9������2�!͓�xʇ@��^���&�ߪ�>���}�.��eah��|s�h��	����v��{[%�z^͞e0�������^�&�q�rFm�Q�Fx�ی�Ӛ1�G�]��S@dB"̒&*�P t�-���>I���eE)����m�R0��H��a�3e��g�����6���}��S>���oˀc��!�i�-뽵�UQ�v~v�����j�.l���nXq"��@�,�Y~j�{m���s��L��3��d{p�;����E�ȿ$w��C��##m�E��/Q%&��SkdͿ/	�������UV%��3�G���_~��N9�zwo}�����������\�3��x�Ѭ��a[s5f��߬A7f��{p���W� p(J����ӯcL���<�n�]�M"��#�~�9��`�O-˚�]��+F�l��>���z�����a�ٛ�,
	�� 2HB@����PtY�F�E��趖ztX��˶����n�͠�-v쮹�-��`).�$w��ɰ�nH�b2�f�E��������f�\/1��6��*�K�o��x�F|v� ���W	�P��8Q�QD�r�U����|~_�~��>��!.g6�l�m�q�T�n���B�y�>��⢧�Ȏ+�m�"���Ɗ1�k�ل�&*GQͅC2�Oɗ����mix�Y]��kD�v��U�T�Q'61UŚ�%�߉R;s9(���jH�e��	�R��@v��iF�%�(Y�n9#4q��E��9�*Wl �H�n!�q�41�V,�k5N�����}z�Q;���Sj����B�D!C�:�+����5�3�V����҇��K��9��17�����xng����N�:}�l�}6|J5�?yG�>ܜ���ڨêh����n�F>
*�Cӱ��f��2o�(��?�����~=g��}�jM�?̃yv���O��RP����HG�W&����o��^��|��������p�P��P�;����k�"��y��:��'ԋ�z�#|����v�n���ߩ���4�G���~��5��/������8�^���X���\��Į!���T���2�5G�9ٌ����|���o��e�F0�K5����_�ޅAS>�Blf�5��(�E� � nTd����[6�fTثh[�f�d6VѴ
m*ڑ��ݩ9�ګav�K�,��j��L��0M)��U#*�U�iV�4LTe��ʌ�ThiQ�ʍ#*4�U�*4��0�UTʌUKJ��U��ʣ#*0b�&TjeF��2�FM*4j�UZ��*���iQ�2�b�QZ��L����*�Q@�^-���k^D��7b�d�K���L�c��z�|����}O���!T=M摝S�:}��� o���?#'c�W�����@�ZW��?>{?��_�Y	���z��@|z�C�����a��?��56|V�?��&D3I��a:��!�tZϒ�$?�y���}?�͘���{����udʟ$����1&�?/��c������<�|�����	��=~,=dO���������>��ڟ��������M:>@���6@P�ck�{����Y?��v~ߦ�=�ޟ-��n~����z�3�ɝ{�8~HG�\|w��O��;_}�ל�����]�CY<?gcHѰ��G��?���"�����@�5$ @��Se��v���5�Q�r��>���^�����tMQ���1RH�L�BT�(��U;��q��1�-��y�FP�5��f�C$>�Rv?y�Q
/Q!��<�}���tKG�V����D=��}?����;z������y�E��#�������^�����P����O�M����|�)��~��F)��C��ϗ���������*{�Y;�����<?��#g��(��y�lY��z?�On��l�[��\����,~3����
��Ր�>s6~�W���_���Py��hO��{�Њ���7˺��n}��3�(�>y��c��U�\:!�ϳ���J������������h�v��zD���~>A�M��s^��y,��M��Z#0�Tp��!�}<�Ӓ�����,�v�O>2�!�	�����ɰ��zG���ԟ��/���<�:2(G��}u���0����	�c_������yhA@CПY�;���t
����V�7@k,7�9�=��>>�*f�>���!���R&����7��ܑN$*8�@