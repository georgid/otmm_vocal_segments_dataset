BZh91AY&SY���_�߀`p����� ����a���      }�XIB
 �(!=5.���P��*P�HD��R�%  �PP � 4            �                        p     �)UI\��+հ5A�V��Z:�C�u�(=0��k�j����mc� 7} JUUEDp�;m�U����W4�U�^�n�*�G�5����L�+J����JR�Z�+�(V�;٬�v�:m��l��h���ݧ�����p�ސ(!N#<��1�t�9Y��:����f����"��ז�=ڋ9NPt4��w�]4�+6�ip �AE*T)S�z�hq�Qp�z�םg�]��E�ݷ���vU�%��"�����ͷIu��{z�m^��������+�� �z	I)p-N�*um������ԬuYK����< ��[���z[W��!�7�<ɝ�ymn�R��x�(� ��qt��uVh�Sgj�K���e�ޖ��yU�{U:{<��U��Zw͏lD�cu�KO  މ(M���hy9zq��U�/{�eHgL��ݼ�t5���eOr�ݣԫm�Қ��=���W�>�RT))���/�Ҝ���z�8t�޵#����ݨ�z��]�9���kӪ��/c�u��=�x oy�%N6�zl]y�קK�=M�x�=;+r����\G�o`i�0ruF�@x ,y
��R H\q����Q4�3�z@�t�y�ѽ�ֻz��G�l%C�+�3T��          �!�%)��h4 �dhm@O�J�SL    �#��UD��C `    Ob�HR��44  � ����*�       �!R�§��B4bd� z��O���I �~����\���W��=�xŻw�"���������#�QU0EU���dW@�����?��-��^"��"����ޔDU_�� ��B��?�������H��*��p��(�����(� ����{ ��`�@�y	� '� �@"y ��
'��@�d��'� �Jy)�*'�����y ��('� j A<�D�P�O!A:���DO 5�(�@"y 	�'� �Hy*�� '���@���@�@O!<�� '�����������P�����!���X��!�C�C�C�C��^G������%$%$!y�BH�<�<�<��@�W�z��W�P�'�������W��H�<�<�<�<�<�<�<��$�<�<�<�<�<�<�<��|�2 ���@�@�D���<�2P�@� � �@�W�_ � �<�<�<�<�<���P�C�
P��@�P�@�P�@� �@�JG�C�C����C�C��J_%!!$% !$%� ��W�����_$!2 $ O%|�<�;�<�<�<�P�������'R����S��C�C���C�C�C�u�!�	���R������$O !!|�:�<�<��@�]�yy y yr���@��H�
y+䁸�C�C��C�I�	��!�C�_ $% Ny�@�@�<�<�<�<�<�<��O% M@�@@�H�+�!�RJ�+���C��C��_ �G�C$! O$ O!$ {��C$%$%$!$%<�
 ���W�C�C�C���V�<�<�<��D�@�@�@��
W���C����C�Cȥ|�<�<�<�<�<�<�<�<���P� ��@�D���@�)�C�S������O$)����W�G�z�<�_$�DC�!T<�P�@� N�A<��C��?�_���r���������E�1����>S�Ii=C�vP��
y��O�9��������]���q�a��ׯ�	�g̘���?lao�{:�~ma�%_P��
����yT�gs}Y\73�c�cۓ<���t2DY9�Pv��1g;܇��O��w/��U�e�/��֮�>�$*eyW�w�ϝ�ͮ�^O�w8AA�K��d�׻4��99���t��]��)�{[u��3d�k�zA����1�
0Ӑ�bA��Ǯ��8^>*�=�=g�J��B�h{ ����B�teOb���u��a
�M��:*<��k~��kf6����֓s��a�u�3]�15a��Ø2��r�
�"$`U��]�M�w��ΰ�MZ�� �r6y����'�+4�0��!2�r��[2�g23�dIE:�(�LU�N��Y���[䄕PU��1`�͸�@�9�a�K�r �D�@A�xvr��~�e[E��H|d8�E�4�}�1	�:OE^AHyDz;��ֵ�\#rMx��|,Jx�4^{�!X@�x�.9Ӂ
��:��V�4�5�8s�/����͉C��;�F�AX��/=x����ժ\�e�gw��3Avhݠ2Ó�ܥ!%9��XkMZbzDQ�yH��" )ĺ��Z�d�N�ѩJѡ�a�ԘQ�i3�F����X�rp�F�;#[݁=f�N�M�ְ�A��10�$��vV��9�C�d�	X�P�!���9�%)
�2B����)�JR��)J��5�GA��zz-��ȓ!�Y'5gfnݭ���9��%�m� @Z=_�����<g�ah_Gx�#��O���f������9E����q�������Ƌ'EF�Aө#��`�`�,Xkҽ����~BV�z�q�5��ڗ��C�u�&䪇 8d���n�;m&]zoFO�a.9�2���IN���x��"��(d�H���<��3N/!3vT&��9	����	BdE�d�FK�]�P��)z,��3,b���d&	��)`�A���=F�ǥXS�
4G �$�8�dC܇���#D+� �;ʷ%~�W���x��!9_]�@A������%� ZE�s�v��'#��� �`dj|tކZ3�Aw�2�F蹾�{s�q�Eo�^p�[�v���0���c��>����y=��'�ߜ��`��$:�Q�c����夓1029ֻ�]�߇��Hիn�e��G�e1���Rp�a���u�3Q���h�˝�����D����p���2�G0�A=�e*&׆Z/`W�����j���,|T�X�<�	+��m��T/ȱ��\��j�䫺
�����/�����<�@P+�$�\�#��Y��S���E�0D�1,�Wk�*���B��)��"�Q��D����J�E�<|x(���{Mu����2�<��VV�&��Y�μ����� B��o����:���0�|�o.X�PN}���3�s�|�B�zE�X�P*����_pgz�t��1y��~L�3ـa�N_I�����S�7Dv��P�A��<o�����	�oF޻��.	w�|'&�)
LL�!�$�#'N���1JB�.s��ӆ�μ�g,�ь��j��U��׹��Y����B5A�;�=6�gQ��#lt�N`e����C;Fy��=|�Şn��ʛ�� &�1�P躝�
<D���).��n-�k���2 ���uC�~,_-�Hj-ŀC��)�+n;u1A�hv�u�w�<J&'l�;�ǿ,�o�Z�x��`A��GP������ ,�@X�	1���8�q1�hw�a���m"y�a8!|7H�|�Ѿ���4�\r4A��4�\��"�\�Ĝ��Pa
�D&'.��Z�7��;^p1�5�GF���:�=�2R�bfӇ\7g<4xl�NF�2ԆFC��2�=#�aLcՓS4d=^��o׆��TZ��|5]�����vv���Q�\�RC�ד=�����ꂇ�v��x�B!�s�D��X�2:�!���c�-��Q�z`}�p��>aK࢏8S�;!<d7q��e0�<a����\#ɢ%qXW��2�G�������W0�-�ݰ.�@���\b��d\dK3:Wn�b��:H�����{�J����0T�I��1s�*�ܪw��7tN`@X��+��3�k�c#O��0#AJR�v�X�:��'D����ִ1T�P���JB܆ud7�ǒ���	�JC����K����g�!2S��Ԧ�3����M!Bw(�"7��!�E	��P�RBl�m��Ӓ��٪篡�W�QS��ܦ��v]�\���Ԙ�A��uxvl�Lp##g-�g�/���'u��ȃ��h�M�\��
�
�n�5==���:3p���理�~=���o5Y���t��FՎ��ĹV��>�K��O�w�yw��{�;����Ώ\���ޏL���P�5%X�x:���&���<;��`6x�H'��<6l	�b�$�'IQ�s��_
��|�-�|�,�m�]�T�08և�׆&�{�
�98JM��bKbs�Ƞ�J��`I���G� �Iu1�A���Ӫ�Zδqw	A�k|7��L��F����z�9j�m�:k]h[����#�z����(u90-f6�y��0�#	2�l��'!��ѱ�!)5�o����پ�M�KK�2r
p�k��<ӧp��ɻRuw��n��9�ww�G
�ﳓ���p�F�B�LY&d��2�1y�4x�s�QDT�w%�H)�A`l��[y���5�M������q��T(U ��2�g��qPg����`A�Q��ܚ�7Ȓ��m�.8BPr�u��Q�٘�7��V&FF.bj�������&G���,8��|��*�!>@1(ӈ���_E�:��H�\\.�d�j�@�������M��;�gx�����8�:�'�ujMɓ�� �ZfTt<��A��r5��f�� �@uA�B��������q,���D��WF�U�(x,�Z	hr��rA�� 4��is�!g��@��  l[���9:y�I�����zM�bd�F�����u�a�����r��F��F��nq�o�܇nw�q��F��Os�z7u{��r=��T�s�u���*c�]��d�5l8zF�t�>nñ�ޫ���e�<ݫ���!�h�;�y�4:�Q��본xu̞C��;4A��:�-;�G\�i2M�q�k!�.A��<l�U�5� ���2�[cPs��!� D*�3��P,D�N]fM���\�r6N���i�`I����&�F�z@dg��"��"���Y��٦﮺]N��'��Q�d�=3Ԯ�����A��ö�@�"��$H[�E��a⏐�qԄ[N{��5��h��C��rM��;�:�te�)g��Ք@�Wqr�WD�[�qpGN��hٹ����p.�ղ���C�dh;7w��:��MF^o��6�^��袏=0���0��w:�tf�(���F�A�A�UI<�F�O�,;�ͻ\�&8��L�r�	������'�]� ��FKA��[�g$�N��_�$�Es��%xxz6n�#v�AkC���]��z����m�|�ǐq�s��֌jq���8\��v�N}!�vY\=�E.�Kg���p>�Πe����O��n�^���٢z����<kWRi�{ːx������g	0��wK9C��,�<��&�o�\lB8g�0O��8p�'f�:k��gN�	�	�y��ʓ	Ȥ�α�ѐb�d%)@r�H��r\���9&f����y��\��k��	I��(�.�4�7��PFHU.� �V���&C��Y�Z�Hr]9F�A�V@k#2�N�cޣY&����%&S��N�F���gy��	�Nu�ݸ4TӸr�.�'�� �PT���=r�G�G�w4nUbw:�a�X��9�<�������`d0:*�\�)���w+�e�Ud�-@$L���tRN��&L�D�+�	�ALJ�h��t���uq�|��<�0�n]6XOn�)05h���;�ᎃn��'!�}�#F����G]���gMD0��&���n���$2L�޽�8ws(0r��^�jIe��QeT4vL	1 X!��w�bi���uv�Aއ�4k�o�KG�A������RaFF�N�㴷�.��q��g0��ӣ�C �uf8�F�W|�5z��1q	�D�B.B9f��+�w]��!���j���:.�7��G��מ����Q�r,��sX�gY�8ɐ�^���-��w�t=��G�0I��"�ǎأVu�Q��̴bF����I�&�0����Y�7'ݒ��4;����pc�����մ��0�JB�&�,pr\ra�,�'N�������N��"j.@��"�@&E� 6�����kh,ۦ�뮼�8��!�u����\�.,e�:�ߗ6�;���%7;�zs6ܴ�8f��v��d3'(�4��:�n3ސì�.��f�̠�2ՏE���4N�Xy�{��]p;�#8��<���I990:�ȵ���fsz�F�ݞ;8�ε�Ƅ�G��X:����uc��I9cA�����:h����{�r-��Af�2u��,�d�1������$�=���0��1ӬȂ2t��`	�<nIfk�j�o|+�lN���5������	JR�Ky��1d���N4;ڀ�a�m��D�Ճ-F�sa�X@d����$��K�P���(��h{Ƭ��j���Χ�c>#qy	�@P6'�ٜ����ng(=7.���{aN?ٙ�{|����N���.�Jl�w%��IM�fk�"����󋏸g�_j�m�!5_�jz��N�=�Nw��L���� K�ׯ�0v��
M˾θ3{\Fد�DD}/��w�W���w=}B��
S�����Vg�WG�&:��+���II����_���GA{�E���������d)�3,�{���H}�=!K6�kl�`X���kW�|,�"Y�����t:�t:�C���w2Kh5&��:�]K1�P;�!mY�H�%ؒ( ��@h�!e��<�ZZ�$p:$2&d�C���t:�I�P����B��ox��׬hP�j�۪^̳T٠�d�6�n�n�7�c��z�orS��bI#�A�@`���i:2�X~����wD��.���*�`�Lw�sm<������3����I
���t:�C���t:�C���t:�C���t:��$�m��/�۴O��:f��?�a�@�t:$2$�C���t:�!�@�t:�C�$��C����@R�k�6h���a%���� ȗ��wv�w]B�'u΂)	���	$��H�H��$��AD�(��\��� p:�C����۳�VzCRh�o�;�4l".��I�ݬQ[�<���&wn$�+� 7u����0��/Z���P���6�ַ_(��6�5)�X�Wq�`|�TU��Ɇ�J�r�x�t�V��-�����н+f� ��L��8N��
����|cH��Я+�;�Q)b=��r���k�o�����eZ��˗��>RK�W8��f" ����R��a{kn�3ɐ����Y>���=f�
��P���ɚc����nj@�{����z�n"B&K�Y��=耹�16e��G��$L��_0N\mb�7�ѱ�\����O�9`�⥣l��v��y;��'�#�Ixw*}.��j-Ԧ���I�M9��Q+��	ֺiB�y:�t:	>m���)ǁ�׎c�����Su�h� �ݥJ�Q�>�A,S�[�f#���w�ŧ����8�t:g(t<�2[L�_Z$�4 �r����.�|j�[D�Yp�I2CT��F���D��R�4:�t:�Qyok��A ]<I$�Gwp~�Jh��Z$S�:��}q��ts��h�C��=C��-4�����t�%��t��t:PwL�	���������3C��]=C����8ꐙ5u��5(�t�G8]�Y���F<��$2�m�)�;���TOP�f�L�A�C��Α�΍W]�)�k�.	p;�h��Y��H�:��:�S8:2Z�_Z$�0:S��`XI"@�$�`�R��݊ 8&��Q?Cc�m��o^�6�KV�FF�#�SĠ �C)��� ���g|8_  }�G��7ݖCQ],�0h�Vn�`�}��Y9Ҁ���]�H%���$t�a�y�K�,�at�`�:�8��]K�� Q�� �r�٢��LNhKwP/MJ1}]>ɽ��.��w83F���v�:�[8}�~�՘�a�b>!F��@���l.����ԉ�����C�]�k������v�~��� �݊�:�U����y��Ɠ�����zE&��I�e�j��i`$��2%�lquI�I`iHM֟Q{��4��.����F[�M����	p�`9���R�N~�J�BA@��ў�s����>��[NkK��g"��Q>C���ٰ�#���f�n^���
�[ےܲ�`��xb��� lۇ�x��%�c����Z�<��f�X�5��C�2s*x4���M�.�-K��b*��Yb�&�z�Z#>��݄͌)����?&�On�1y�fxnL�طV�R]��� [��RR:A�-���{5׾ս߀H�uw��_|-�I�K�����T�ZJb���<�< �ޙ4Ơ���[D��d�I=�����ۊ�4�*�� G�̧��N7كp[xm��A�3${w]
��g��o_k��_���J�[$��}��9����a�ɂ#�7w�-:j���5Ϲ;+�p�q��ˁoxm��3"5�7%a�k�Iѽ�[�����ɯ���~�x�s$s�S��㊜����y��ޜȷM��uڥ^/��ɽ��<B��+�r��&Q����g��![�?_[�r{3�;R]}^un�����Á�37�~���j�:��j�^\�v��K�滫n�{_%Z����v�}�-K0Z��Y;���5�=?n�ދ�� 36����9�ه��+Jy�$�a]��Q�{_�
����H:vK$xS�o/�j��v]9+Ƌ;����{�}�v�G����BI= b��xF$��\�E���T7�d�o��@�{�zn�q7GT-�^	j���H^����p$ǄN' A�_�Y}Q*l��c$���땑h��>�&��ne#�x�C��K=���#�\7���U���kj*U$ƽՖ�˨ۤ��C���&k����sm��7����Ɗ���`Ufzq�`��w�<k�粽���Q��z�^��T�������;�/�y�Q z#�����ɇ?m�����4�6�����>�Cq�"�=�j�c0���xD� /S�;v��N41��8�x-�8]�N�~�u�s{~�t�%n����$�	$y`�
�C��I��/.�k��B���?�)` UגbP�w�P��H��9�DT+5$���=HΎE*^�{+<��'}ti#\7��8̉+�>��f�Te�ww��pf�Sḿ�k ��	á��t:�C���t:L�+"q:X4H�}%�ڕO7L��k�x0؇l���9�,�dº�=^�iz&��c���N�\��g�ۜ�7�70wb�S,i�D����j�9@�p:�:�C��A �t:��^t*%���vKm�\�q��م��n���|p�WG���`�EN��f{	��ކ�'�ձ�F�y��cIyc�����  P8� m�l��zi���b�H{B��(w]�<���������d�����T�`m�IP�p:�ǹUh|�ᬤ�d�<�����t:�d��$�]��ɅCo��-�$�C��j6��CZ�AP�t6����w}ń���"�0��Q�g�(1ww�َ���S+�	ȉ2WM%�p�c���'wB�U<]?V���ۿm�9���p�`�55@`�:4Ƞ��t�!� R�@��h��u<H$�C��l��6�I�@6�'��t.�T�7�f��$�����1�[���~��$u��=$��3uZ�;����C��$�Z�d��sSL��[B�ɴ:�C����8� ��{����-�Ѭ�(��{���V1��)�z�sZs���0�t: }�\s�����R�h����N%�y{b�r[��h���N��Ƀ�Q�"�X�q>�?_;퉽���4��{Q����'�4n��A�a��=�{5WsƗ�!KQ�w:;���0I�{����{5����ڔ��� ?�� ��4�����x^Ν�sI��������\�۩�Eibէ�Os�<;�ɼ/�HEj�UF	;�A�=<����f��H��c1���t���o���'7��oKC���P�^�v8g�pݓ�VK;|,���޻�s:�b�{˽� X @�y�2j��y-�Y�Q	�o1�� .��z�F;kJ�Ż��c��Y�҆���1���T-ݛ�Xy8'�	��":�~@�^ݻ���vgw�\XJ�k��������h��DH�#{=�){��{ws9Rmqv�ܩt��Q/���wq'�̆**�r3	�� ;<�t
�e>���k�ٝ| �^��4͇��3��םû������яcU�@BRg6nU�$YwOQ`=��=nbS���ݦѯ����9����y�I� +�7���G�8��
�C������C�9@�p:�C���t:.�D���t:�C�H<�(CSTI΅E���t:�C��L� B�-�@�t:�C���C���t:��r�@���C�?��6�?  }���wgC������ٺ��f6$��j8!m![���u�:=#DM���_��-
��1$ �:< U3�
���:dP(	jI�<w̆I;�$C��1DG<�%;�� 7f��򀌻09�D�c��F�c�����<$,%�e���NI)��ovN�:�c�	��A����E��|�!Gkz_�,��F{}N� ��aذ{�o���}�a�@��\��Gvn^����gpI��Q.���<�&�:{���� 1��c�{���n�p:_n�m�hQ$���0�sw�ZO�d�m��ܗ|�I�� t:���7��ڗ,t;�(�����I$��Li<�<�0�>$�D�̙�L�;�r���ݑ�����t;�N�w�!>��=����@��� C��Qy`��1��H��:�C� #��L�ܢ>�UH� �����"vHLD>� "�n�LH�ہ�����K����g��d3ua�T�cD�2�'B����n�`J��{���f�	�C�����|��I� �HEf�BT��%nogi$� ��M5*%��O�t 3h��Q�H����z�F	d�B����r�r|�Ic�;�.��5�<��p�p�{�ȁ�{�XF9�{:0^��hb��L` �I!���5�D��cB!���t`V�
�EümKZ^Iq���6�i"/{w{�g�ۋ�)�^Jx2���K�J�9�B���e-���7�� ��mg��F�=�aV(�:_\��P �f���Pw��ܧ�B��%�w��8���n�u�j���<�̯RY�u	�C��ٵ���5lp��r�$�K��>��,�-I&;��:/)]�����u�k�@�_qSy#��С�w��tPU_i� t;��� �>{�%�r��G�T#�]�2Ia�\�s ��@`��	o�lH�H�-$�3�rgw#ԓ�g�#ܻ�B�ڤA�I$�^FN�.�;�Hl:�����t}�b��K$�}P�h~� �@1���q�:�'�U��Rlr\�B��	��_{�M�>2)H��z]�;��$�\0 8Mť��
K�G(�:�E�^�6�$�����j��ͅB�\�Z��w���t:D�P �r�@���֫L]�Xԥ�2�Iwh�BI�Ֆt�@����z��F�u��Fɣp'��7�-�m��a�@�>yծ�8���@��C�U�$%�I���t:7 ���%������*6�<;7b��S:&sR�5�|��wor�9f%TyL�j���x������v@���)�%$�"��잢 f���GH��X�8$2Ԣ�{����f >Q��p:�^6��C��G��	�����=��=�;�(䳙�I/74ȼ�qڶ(���JH���nͪ�=n�&�l��&�2Ξb��b���s�	4:i���6�C��·D��d\64�+�  ae�����t:�36@`����A  ��m�����i=©�VHs��0H��}r��ӛ�]���
�CܣL()��(����^s�����n��P�J�Ib0�t����<�3\4�'
�fqLw	ڸ��:JPJMPΐ*�A t;�C��`�(RXMU�-�A�輽�L�s��..�B�@V'�&��O����}Gbi�b틊���t:�n�;�z�P[�/+]@fg�a<�|7w��~`��oi: n�N�B�;���vn\��9.�ӥ-3F�Z��6 v )�t�7�}(T4�J��$�%F��M��V�iV���t0�a��2(y�ID�@�<�@�:7u��CZ��wwG�%�J-�'I����$�9���שOk��"7kHf$-��]����B[�.Y ty�}��=&"&��6�d���[D���t:�C���t<$�I,ww:�|�d��`�8.\�\���q�ɪ� �i˲j��wA t��ڒ�yP�&kQQh|�6[4Zg���Z\#n�h�@�t:�D�C�U�C���tXa.�γ�F�C�R�ca��E�#CA�-�I-�@�t:�C���dQG�`�5%� �5�0J$�C�.��$��x����0	������<�y�l�IH�4Ha��i��0�A���$���!Ã2���3{��ws���
�h�C���vKh�Kh�:ԗ���Ӎ�׺�֪oH�2{��BI$(��I ��t:�:wht:�͏�wj�'��_@Kz����d �'p�j��d���?�ze�/`��@��de���Bqv�̪��H(�	#�K�.T���{8-�>p��|����9xP��6�G�ew��`I�u�X�:����P�q޼�At�f�-��=#j��ʗ ���p%,��o7�s�� `s�`���|����$�m�טq�S�L�=4Լ�{�o�����w�4	9�6�m�U�f��= |�ټ���rJ�ð�$�x觐=j��Pz��C���$��r�D�K��Fbם��}�s����	'�{�>�\aQ[�ܭ�z�Ƃ�GDC�
�<���C�	̑�\�-��0I  A s��Mұ{ϐ��E����`�:�C��p�ЍR(�O$���4 �p$�we�`	h��L�גѶ�k�MݍM�[mz���^��,�Y%�^E��L��1���$�B�m��{��\<����
����t7R�8���QK���~~�� ppp��� (���s�?��T �$@?��X������޺�C�x�Fӯ�� �(F9�u�GV���Up�M����k/M(w��|�!�y���W�x���{��N�D�F*�jx] m@�3J�h�� z�i8!�|�@ɍ��
�#�N�z볿M�K�N���K� pڈ��� �C��|h������@�NpW�C:}TCL��:/m���Aѱ@�-�mg���(�z��`)y���{A�"F�Nx
�^����C^�؀�u���^����i;8�	���O��p�S�Cy�pW]h
�Wo�A��_QP��]B�<N������b�@kã�=4�C�v!���F�bbZ&b(<;�Ch�'G�IL�X��3�Qک�v
|I/D�be(1[1��x���=�l�"�@@�$ )���E3�G{SA�<�C��)���Sb<�ﮄ�֎r�t�H�I�D�T7�!�C�R:�	���(l8����9�8�6�����ok���QN����1$I��� &�;�D<A9qeS�TM����]����E�a�u��m^�#kB���UN ����S���[�@�y�*����N�M <�:�PEU��o��?����������������~���J~�Y�?���7(�
�P��"HHH2L�$J4"�0'��LL�%I�B�S3ELDP�M�@P2CBЁJҲd-	HP� �P�PT��\�)F-	I 4����@�u :�J�eNJ��1��oXr�_G�o��U����Vw)ݛF����%�E&\��W���55k�!�ݲ�ֆ��N��qa�sV�+!/V�˷\T�t[��ip�TPt�{#4S�v�����T�1`�E��\3d+@�^.-�7ٔ���b���+�)���5;O)]߳���_���u���W�p���٫��GZFY�`���P�J��;}}�o����N�pn7dh�3�3`ήr�.�S:S	Ո댛I��p���@U6�#�ڗ�%�xً��zi�5�K�	�磄�gc���.�GUGu��.iR�q9�3`e��q�p2*[ѧ�^�D�9ny�K�^�I���Kcrp�c�qԴ\��6^�4�����Ü"<g�ȶZ��h���Jn%s]Y��9~{�1E��GI�^
|���I�Pvz��
�b��A_1�)� pW9�;���#.�]4z�]�7� �I��f##�x�[L�7je�9�5�����D玶=O[]��#���`9�9r��� cF�L�k=��yz�)�G-�u�9�F�u��h���onv���%�m��A�ͿA�yD�1"���̍
�}��>���̓�>~:o��cI9�4h0r�J#1r��M#���{3j�Nx���4�{3���r:<�c����� ��~Yi��$j��J�T/�1a�i)##W�wA�E�=�rd�[(k�K�E�}��Ç1Q�y9���%�3�{�O����.M�.�Uw4p� ��{�:Y&�2�֌q*��E�jE\�P�g40G��s/4�p9����OB]���fP�@��ۀ���%���]��o8������y���NiWntcmزz��{2�z��o =���p��M0�e����s(�Zj��!NB�q��'>=LƞS����m���߯��_rN]��?x�>ȌL�fHI)�[�Ckd�NP���K�Ýa�߿�����]r�߭��T>�^�M�e�Ld���W�R��̫'�hwHŢ'$t� �)\��g3;�LA��9��r�*��xy�һ�P���l�����
�����-������A�=g^�xM��~D�������'�Ma��O6��b��Z簄��Ǳ��f
�Y��l�yi���J3Go�뮮m�{��l��)�I߿{8v��?F�'=\�v��^�o�觴�e#*�QJ�FJ
��0���(w�c����*�59 ��!����fP��A��a���=;�1�M]ԢI�Cx��5r��,�[8���o̾�/�nܪd��d�J�S+Uv�I���:�Z�`b�VЀ΀�Pn�Q:7I�l�q�r�������8 �zV�h�g*b.�r����'m<��1�v�ġ��n�n���i0e@��N���t�E���l�0������v���m���HaO�7q>V�&�c�|���9�<,��cR]�H��0��3�ٳ���(f{$Vw��(p�}1�v}ӫP���"��%�I�F��{��9�eu,X|E��y/"�E�$�I�ܞC��g�A���r���U�d�ĕRAO0pd��?X����-�{<�Ktw�)�o3��|��(^w0CF��Cۅ`�ӊ��N(E��:�6t�\wi"�I� l��f,0��"��FdPB�d�	�^��������A�⏟�Q�#˫�E�jFٌ��[<p�&�o����9�o<K=Nv��DQAό�Iym�PT�.�ڒ���z."y�y�f�3�ܒ[I�R�$�#�[*D��d��o�h��Vfv�WX�'=�&�bTuHҌ�%��/� �f�w�1[K{�[���za�ReE���������P�W3���[hHX�QFڦhw�c��ey����NY�W��̑����z>�~����G]����K[�j2Hق0��s�����g=}��p��G�*s�TID\EÅ>\j!�d��,A%���,b��9���[׻C53[Rn�n�����f�|�Y� �$�D����=��v.!�\����;�{+���=�Z�q�*����5%a�'+32���b��w��,�-6f4��=�n���8�W�O���zq�#b*)�)��T�}�n]H�l��M�������ܴ��-Ba@���yv���{r�O|8\���8��S�qɘ��V1�FBJ�fd�����s5���tn���NEN�$�
�ufo9�͡�͜}�Ξ�����Z)% ${ٔ3�f$��s�~���'O{���爐���i���y�!~�N]�y^fW/��ce��e�Ԑ@3�Y�/�| c�Ƕ�nD�����0`q@�"�P�|��*�{,g��*�l6̩4݂��wN(R�A��R �P#$��ǧ���B��f�i;�品{$i��H�Q��*�2��n=�w��r�{�o�b)��I	#N����������)�:7��������̃�<�������X{C���<�&��a
8Q����*����;vu��\����ӞT�j����*�=z��&q�u9Ҏ�	�<�è��&�ۦ�{]��E��y�r�ѳr��	5�p�0���Z7�G]Y#qs�ݒ��5\� s�y��G����N
�� "������c�*i-��]��\���k��̞e�&�???���fc]�+�y�.I N	#����pS��z����|��\��#���s�{���;��g\����Z���)�?[tw
L��&`�eS7�ǎ�����1���/M8�IU�Cy���sXG�����a�pp��=�e�E��nM�+��Р�Pd�C�O���@�OI�ҕ�s$D��������_r�X�9�7��y��~����dMj螋\QNIŨ����8�'6���|͹�zeCM24S����m�r�n��
�'Gmϡ�;Zޝ�,��2�F�6���S�l�.�`���#�$�&穰����˯�<r9ݞ�Z}1��u����wzh�.`z���h�8<�m;C��䊵�X{�����TD1���cH�ﲷ���=C��9��/H�E�$�	Q.�g^��3q�:� �G�جn�)iQĨ�T[&�*���.hʨ�Vn�sr�<����g='����$3w�/�c�^�2�N=��(���nK���1�|݂�n�ѷ��77;ގ[��gQ�M��޻۸)hӔ|�^G��Wfeb�\�����/c.)-�"�������/�s�@<r=�^]�@����F��� �C�燝��!���{3ha�Ԝ��)��F2�#3�UF�7�!�a㞹N�8���ps��=���n�'�z7n��*���z]��4i�}���D6=�n8{-ܵ�� � T,�$;��:f���>̀_��cb2�,4�q˾�)E~�F_r�X�>����Tr���MPT;ҽ��}��Ü�|�3�m�������rB��9�mI!h�5�a=���aZe�,p|c!�y�Rw�@YI�-�|�Ճa,Y���&�8�h�Cya��I��֞c6�k�Z�[�3K:�Ɍ�A�8m�{�5��V��t�#3�[M�S��bn(���9�6ui���9���d��0�"hѥѥ,��h�^LK�����1(�bl�$ ���Z�;��G9!m�<�6b�S�e �����ӆp��O;<��'Ͼ���,Y���9���(�z�8���f�4bӗ�2�<����B��/�ܶ8(ڙ�{#�y�A`ւ��8����!׆�3�x���p��n���5���\Dt���@lE�:bh ���DF�y��ٵp�b@�������]hM���mWbG���h�ٸ(,mI���dV���)9�5���� �+��nnH��%��%';t�5M��\1��[W�'Z����\�(:�s��
�8��3�p����kZ��W��CVT����Nĳ��!:5k#��ɸ�ᮌ�^��mҪ�6��<"[ѾW���Q�a���QZN8�T�r�a^5����hy���_5t(7`n���Df���k<vݵ׈\M�B��<���b�N0m���'T�U���WB��cU=��a^讞.��:^:գ;���q���Z(�Y�3Lp $\�ny0���e�"t�tlr��E�X�Kml���Us[+����ժLŇ(N`��֛T�&K��*"���0�u�e�·5���.��/����n�Kc��l�:�F�0�6�B���a�*�)���*APY���-��HT��lB���[I��+s��ۚdJ�r��;�g� ���=���g￾��q� ���� �4�o4��� ��(m\׿z(`�> �f��t ��T�Wz9ځ�u�S�����@�s�\��k��r�pp�@�w6�:y�O���M�� eM湼�o�P}.I��o�NJR�]����)I�~k߰z��{�ݛ�����Zu�h�x*՞ �Ѫ����$pwr�p"	P9E(ӎD��W:�8LS9�څ��F^]���h���aԥ$���ﵡ)J�1��
<�$��g26�������m]4<�mX���n
5��P���߷��HО����`���A���0?�������_~愮y��ȦT�g��شM�D����8{�K��R�<�o��)߾ow��y.�i3�t}�R~!����ֹ��� ��d�� p�f?����^������=��������M5�x���r�a
T��rG�[Zh�x�e�y�O^3���u)Jw��>�9!	���Hx�'�w����=����3��S.�,���|�Hg�<��f��b��inNKu%Y�p�q���9������ϭ,d� (�5�//�x]ع;V��Cv�Zq�@�k���s�mWD6�5΋����wV�kq`҈%�^��7k,7�of��\P�}�7�.I����8���I)Sr� p�=��b�8	 ������I���yX,�H2���� �=��l�]u�,�޿p{�������3���~o�O}���c����5�Z���mx?�(�}��`��'�q︜��:�^{��T����Dp#�w����$��wT6\8��ٽa[��	�JO��/��P�|�޸)I��h���)O<ѯ~����qP���.�����	߾��w	�|�G�`y�!��P:�{Ay�Oz�(�y���x�pW T�J�:��#�@G�=h\= Й��7�&@�}�}}'%)O=��!�O ���iG�,�U[	]�-ȸ�Y/��O}ѭ���R���]�=���!�`�C.��7\{"`f70@�]�}�9�<�'��I�!ԥ'�~��\�u)O��񯷻Z�p���������"z�%�E�I	G<��T�m���ѯF�����v`�I(n¥�FF�k�����)���֏i;m�,.�K']f��{����|>��m/�xn�p�	�S��g8	<:D���.��{��N��^��˨�6��� �h�m6 lW,���p��R������x�����������������:���;�zE�9D ��br(�t 2T�%(�*������؝Jo1O�Ͼ�)�$��7�%�#u�k�LR���-J8�<ಘ7��<�&��ﶄ�%):�>���/py�}渥���nE���8	�I��*��գ[�n�)�JN��_C�_�_���?S����������%�Zh�	'@�=��� q$��@Y� G��,�p�0�(��Q�,�Yf˧j�Q�$D-$�mBD�B�-�Y�s����%�:��}�'P4'�}��b��Zt�Q�=�e��#@�:IT2�%'~}�Ϡ�?l���k �J�w��O�ѯޘ&�h:���^MJu����\1�|��m1
t��vi�G�S����Q�~����hJOn��C�us�����!����G�ޏ5pY�<չ�9jP�Yg9�5q~�%�(��}�r?o���~k�Bd�'���g�u\����R�2�jp�(S� 7F�]�Γ�qL�O}�\�R� ?�������{@��:*"b
!��e����o�!��|�=��o���	I��︜�����rM����"��p[)�0�1.(OD'
�A�s�!%A#F�s�}��J��~��b�)I���_�/P�������2C�����7���Mk}kY�Z����;��s�vo���g��JR{��?�rR�����qA<G�_c�
<���Է`�l�@	Q�QS�J��|p�\x����)�����&104���ZSR>��`�
x��z;� ��y��ת��՛�!h�)ΰ�]fsY���"�����BRw����'R�&Jy�7�`�'�!2=�_���?{��oZ�f��s\ޢ�|4\��q��{�'d%��y~���Ol��ƞ��B4Vf�Yk{�͚��?����O�SR��^¾���)u�k�qMH~��梙R��
�c��8 pu��I2Z�2�ĚQ�8]���D��J��y)J{���ÊR�����`rR��=�7� ~�XHRd�v�#O8H��[�"H[�9�[���z�G�r?����  	 �d��7�㇩�y�H��?�g��'��c�S��H��@XRV!d��=��ߛ�0d4,�Q�J��LP�y��7���j�����`��Xd`"�=���1�!)=�?|�(�~>��A#�9J�*n�r_�
J��;��߸=A�(�؉Hp'��Wq�#�G W�/-_������y���hۍ�m#�Q	�i��Spt�6I��T�����\9Q�F]`<���m��|�4���r��<Ԕ%�؊�KA�n.M�uv<��]��A����<c�n9ӝX�H7U�rdz���7����=�~� ��Q�0�,8�E5��í�.��u=�d��ѯ~�5)�ςR��.��]k�|�%�㑴��>��b��ҥ)y����'~y���JSx���e�( ��� u}��L�>!!i�5e��[�{��;��{ᙾ	@�{�}�������SP4y��>�:8	�8<�MK���h%艹(Y�{�\���Z�רJS�>���K�ew	I������`4'�tk���]��t{凂� ��F�ăpP@Nݻ$o���R��{�~����Ϸ��l��؎���7������~�4xه5�NP����ݺ@�%g�B����4'^���9)@rz��n��O��'�����>�?E�!n %�܍Fk���3��}�Y�8	 ��+��I$+���(��{wF��5�<)w& �;������08O8	����C�G<���M��������Z֍��é5�>�WQ2�n���7��6K��H�aD\�>}D��Vpa�knn��W�a�Z�=�sv�){v�ܛc��ZM�;����\9��w]P-�B\����r�=h�r��^,����g��2k��	�}k����ӯ}����R���w��ǒ	�1'^}��y�G�<���[���7"�@q�Jw�����P)O�ѯ��5)I�ߘzA�J��=��t��C_�,�3z�P���0l��h<�$pQﶦ�8R��{��{���P2�B�/y�5Aמh���)�>�ﵬ���	k\ݣ[�32���H��w�������:��n��;�$��ϱ:����S�� `;�&t+� Qt�n�]k�ԥy�������{���_Kbu�<Yqt^�ƞ6��c��V[ѽ�t��}��~��R�S�����{>��������F��k}������Ňu'�N�W�"��:��y�8%)I߾����J�����JN��G�>f"JO#������ �8��IDU<)���-�p��@y��>g��:��?���)�/5�prR�������u)I����P��V� jPG#U"!P�$�c����R��z��hJ��e�ܷ��(�y��a�y��Ǽ,�%��Q�n\�h�R9D\�����s�;��~��ԥ)ߚ׿kO��'��ԟ�~���������Z7���7�泛ֵ���%'��Oq�}w���m��߭��n8B��|W`��%��-��C���٩y�I���%(:	}ּ�\R�����44��g��aqr���y#"bI)�n7%�D�j��,�#�����r��}��^JR�{��x�d��8	��լ�17 %Mf��淖o�R��]�����$(�ߞ�k��%'����A���O.��j\�A�<��z��Fg�@�Xou���'R�����z����4}�'P{߀�]�D��>@��3h28	����<��y��S�������!)�Ď@�p �wX���R���~�	ݓ����c����,.w��Й!���~�޳E�x)իfHJ��,���}�b��O�q��(����-@�b9�9��4�tq���}���Ǚ ����?~��R��<׿oN��A<�?ڇ,�#�
��I@
T�7�|�:X�z;�������{9ֲֺ�Sp������9Bw���	�HPw��}����JSm����H�y��QC�G�LR�SR�ZˏQJR�~�����M�Pk�~��:��<����	JRww}��B?/��8!�|v��A#�8~"ĵ-����H�^����*�Dpz�f1��ЃA����<��;���g�s��9B������\@�#�d�{�^����R��}�ג��מk~�d'}Y� �C\p�		 ��&�#���o{��屶%9�v[�v���+Uv�����F��$��6B�Y�{Djs�CpA9�(������1]��*֭�I{>��b�f��Ӻ��Y���:����x�ω赁A�Ȋ���T�7�ww���w{���������
<�'����.O �-g9���)JN��=��n 3\�Yu��a6��dݙ�3r�o7�efQ����F����_�b����ϵ��'P4'~h��)����>ݼnJ�����␸�L�GY������V	u��[�[�X��R���~����JO����w��%)�4}��J��&�);��}/ h��^$�@	NT'$̠�p3�x6��Ϡ��Ȅ,��������)<����ߺ5縧���(\� r� ϩo͹$nP���ͫ�&�J��vk��&�-bw�?{�ԇ�C%;�=�ք�)?y�_�`�	O���{!n�	@�F�j�� ��q���;��}nN@Пg���CQ�;������J��=�����BW �h�E1�"�3(��3�Dp�k��� �Uj���!	dĚ�<)��ջn����'*�>����:I�c6Y=Xo&a]^��&������]�^��*��݋|�#G�yk�`h0(#K}ۙg/,��N�m�0Q�|a_;$L�Z�ÈY�޹�C3儳:�s3$�9k�x�l3@�[���z�NP5\Fjp�>Q��%pz�� *�M��F+���4�k�#[-�7�a�[@�!�[7޹��vs,�Qk[�D�.�9���`�"������@��N0Nc�Gy�4XZl����D�������s,֌�z�N>ͦ�I�搝�4@4����^kŹ�s��v� L:�i�:�se��ٜ:�=�		]f������^�n;ԛ�F;���0ޣ�-7h�}4vfyy$����aV܎3��stR�<Un�m1 &�g�V�uA���ɷba�P�����*�	�kj��_o�n�7H T��,��
	�ݪN=[4���V�^ydݷ�;��Y�(�c�qu���y܆0s�	�.r��.3k��鞏!��)�aʪ�If�LP���HN]+�Ed����i<��n�ύ`�6x�P묅.w9*����HH��\^�����nZ`6�`*����[Y�Ō�]�P���g�t�8� �����ݣظu\aD�����	����.�bD��Ԙ��v��/�N��=��iݰ�A�=;Um5�sjv��L���0S�'�v��vי������(K��w}��ow��N��8kGt8�h稽��PUҨ��<U6k}T9����7'j�t)�@(�w��^��h?_�n�؎� p�ch���Z=Q���g�,S���C�+�.���T��cl8?�z_��	+�a,E6�V��P���j~���{���{� n����!\/��{u�����㘥P�4��s�F}NRlfz��싀O�H���Y��-J%AK��H�&`Uۼ�?���2u;[0��3i��{>��5�D�J@U\�:1Jd->�d����ٻl���������v���\�s��[�q�U/}�(��쭴Os6���|��i��q	$f�8C�����G���d����7�~X7n ;q��Ta"rW�1 ��QG689�~TI8|wi��~9^k�p���h�u"(@l�M��mE�#@�o��R4�:�	�`n� �ziT�7�dT���Ͷh�j�dK뫫aIL�$�w��a `8s��#$����)4�!��6s9��h���1ca�`��n���` �o�7��FW����j����##y��8/9��H�TB��h7TO�`l�j�2��#��3�v���mO��y���Sp��5UN6�r������nx���hQ'W}��4�9�ܞ9H��Z�
�ZUm:-X7d��5Q$N:�����GX��Q[���Bap0aa�Q��w|��r�M��ۿ ��KECpԨ#��I��B!�1X�������������O�O}wI�r/7�����8�fȒo������\�tB�F��B{f�� ���6�=��Tb]Zs}{C�-�h둦���i��i����$n��Z�?u��,@<����~� v�@!� �!a D��pp�v�j�'7J';����.��u��9�f��[��hO䀌�{�_$�Y���~.�3c|��88�c���`�EU:!K��'| ���܇���k�c;x��Ŏ����<p�y+o���{�}�ͥ�&�����{��իۭȚ�ڪ��w�mB
j.0و�����]�i���}�~�N�f�{�k����\�'�|�7��R�"�Q�+���m�s��'��m2z�5�&��e|-p 8=��nD���.ЀӨP�'|�T�O�qfN��G�W�ɾ޽�${���e�(T���dRb4eZ_ G9��E��M��RJk��޳Vj<_�6�(�u�,��踹�r-���7#{qVF���5����{X[�8k��۴����AY8��۳�T���+�)�x�s�&'��	u���}!�8Ӳp��,E����J^{�Iҵ�VB1b$�r��8�[�s��p�����o�fi#a��-]�R�Â�=����?�8!VA.7h�P@��Gh@�9먴񧛝�����67Ȟ��᤭�a�}�mi�I#�~��1�{y�vSv���1��Eu���m�'��uQi�ť�s��>ǘ�;��[L���W�o��L��G͋��88 �+�s�\@�D�ok�_ �9�B�H[QRU)7"Q���ƙ$�]Wr�/wo*�>��2O{�����30�#UQ�pp�pך��{���=���9�K/�]Wm�p�t��p���K��emm��]�G�xDU��n�:�������uȷl�7�5���i�A���$�K��/���IhJ8��G�E��<�#��x�8���~�Ͻ�8����5�t`��G��m$�wT+u�tp�5��*�"Cks�iD�o3;�%��u���lV�ݪ�<<�����o=�Q�U�'�8m�����v��>&�^�$��{%�/yܭ� � ��f�;�5�(�T�<���Q.���;�prL̊2I�sgio.0�Kx����-'-@�7VI�ÚHn�۲9�	�hQ6��ͧK��r!!�m�(ҨU�s��s{�$�X9�tO�<6� pp_ra�lo�[�ƊWwwrܤ�K�sr����Z�g	�sq����NA������
U�7ٰOI=^7r���fS.���-�T�U�UeS	�D�i�x�-�#�mW8�3!2ؒ�=�͖M.�\�A������{�f�8=�t�Z7.��TZN��f��k4p����z}H��d�����H��s�,��2�fY��p�C̓y��Lۼ�'y��8�Y��^^9��w���T8�u\�UqF��$�{ {L��9��7��O�hs��ٳ��i�
pf&d$�R�UK=�9D��_/x5�� M Bq٭��(�+Wn㱭�_�87��e}�̦Ne䉄��a�DO߿l}~���<j��Y��L��!�ݓ���2M��Ւ�r߅�s��+�p�w�غ׎�.	]��PJ��(�.�br�p����3_}�>�A���I�z��Ϸ6�Q�\)�+T�'.��}����w�{�5�y�B��I�]vx����Ww�h��jk���:�}�
lC����%Q?��p x ��ӛ,�x+�I�v/)��ܑ�Q��ͨ��٪�TF3,Y'}�MOϾ��߈�A{vvzۇI�qLe	$��M Ձ���~�ߧ�D�g��D���������D�� �-���U�Qtn0�c
}���o�,)�omQ'���z��K$w�d��X��
0;1�F��$������ p�e�̀9��=��2z��d�h�C����ˎU9�h�$���(�L����}{J��m�D��'N��RZ�0��Xf�(�罵��>��۲Ny��d'E�r�h�؍8��"D"�V�y��ק�o��R��/5�eK��v�v�x�6�prQ́�J%$6�7㰰]�nNx�橞k�4�llZ$�vl5g3xwgqᶢ&���^�{m�v�����|%�c�"E���8x8;� ��m
�9'��^$#�Ӑ�ʦ_։�ڥ�ɕJ�3��k��x�a�أTY�!m8�R�9��wW�;��{�3(3�un��R',Բ��b��$C-�� `iqW8i�E�vOq�$�Z9���r4	=��ݓ�iKC�5�T
UIB�Bo��+�  >21��D�w�;H���3�����9��À�uQF�[E2�z�Gu���7�Mۓ��æ�6���&����D�����&�vf�$�1��	ﶨQ� �0��Z=��j8��-,i��w2i��~�>����6z:�]\�vK�46����A�ch���$�1�L���m�-hj'Z��)Y p`<��� �4�k|�֌֊�:ֶnY�TB�Y��ť$]��0t�k�ٷ=�B%�T����%b����+��cR��#�^�׷<��ڴnt��;o��(8�GiFZD�&�wʾ�I>_m2}�L2H=��Uo�1I>d�#�t���.Y�O���� 8Bh�����ƙ$��l�`��Ƅ��iƑ��B��{w����Jԭnk�T��P�G�l�x�4R���UҘ�tqs.7T�{큦I=^�G
���D�7va���I�0E�I�:�Ͷ	2hhw���%\�"s�k�M�a����l���ɚ-����6���ӭ4ѽ����==a2C%�CF [e� ��y������x�P.6F� �}7j�'<�U�kH�=��ہJJUH�pA)����F���! s��ozQ6�d�1�~}	����?\*����g*���w���×�ujhi*R���CF��w�6Q6������^�(�}�y�ȼH�P���oxsZ�kz��I�E`�3�2��^ȁ���or�����p8ei�N���e�Wwve����n��@������K�
���RZy�f�vekD[79��v���F@g� 9��k���N�@�,�,�rO+������￣����豮��������ۥI7d����v�;�5Q&�p́�G�O�p2Q��i*��DiG�e%��A��>�ݦI��eoޙ��/f�lBؒ�tn�BQ6�5�${��2`.9�~>���Ukۼ������]��x#�7�����03P�W<����R9�A�&NȈ�AAI\��(p���0�Ll���gsX�1/E�HBX��s���a�_���ض��Yc�u[�2K�'�1#',��#hZ"�^��"�����
Xِ�� �v�H�N0�b)��8��p���m XXF,�#������LJ � F����3��%$5QA4.��Cf�M�l�q��m��!J6&e@�>�T�[WZʸ���~�|����x<I�� GE��Ӭa�]�r�����H��M�1	%���ηZ��8��B�����#�>�fS��q�<nw]���!��۷l���J��D��EӼ�e'bbU"+S�V"���+M�[�b���%7V}2h��#� ���\AX.ٙs����q	p%�˄�۶��O"`�]���=p�v��X�&�z&�ɞ;>�y֫�c6�̽lҋ�h�u�H^{cq�mn#6 �s�t8�t,	��ŷ)���<�Bvz�Oc�</Kۡ[��*����S\)2<k�vʍm�c�c�#�7V-�u����p�Ϟa:��6��g�@z5+�/�Xj��֧�U��
�ζ���<�#pa2qF��)Y�:5���`զ����X ��V\���,�'9������جK�7'�H��6wfh�F{Pyzb.i+���΢�n�W�Q�J���Mփ�7Lڄ�%�P&r�V.rU���.)NLk0IkZ5)�0c��>v�;NC���0�����S��8Ng�]`�nt��>�nL@/]*���p�F沥����Hs�[� �����t��b)�]P��R;�'�=KY,�eQ='lk�Bڵ��L��괧f�z��T݊��K��Wy��  �/�6��C�@�{�T]�9��C���t��Q���"�����G4)�y����h�����՞պ�F�����a*�m��,ݡ�"w4mQ$e�O$�s�.KW�U�4�)F�4�Q1"M�ٵd�A}�Y.8Ċc�#��v�bɌ��"�4 s�����[�r�$�s%K�ײ$`vc����)�S����`�b,��Q�������]��cv�7�F$�ށz8;����ݦG�y�.�N)EA"0Q$�Vc���[������-{�Ci������jKWv����N��	;��6���7i��d�D�|�/
CI�
N�n��{�v�9��ǅW���^g�kK�y�bo��,��$�,
�����l�ѳ��P��1�Hoh~~߾{;��?�і�<V�/<�����HQf�ktƺ坑��e�c�ZS*�c�c��um�&,V��N��/:I�<�d�X��3&pu��[�&8(8ĄU�q�.y��{&�y����OS���!���/�w�����8�|�i��׭�⑻�uL8���dH���t�qE�F�lȘ"�� *��p3Co<�ȃȳ��d��em��i)l%��T�w�<tՔX^��M�$���eZ��n�'s6�3��G`��I)V�i��Nyn�h�=���>�A�6��j�_sj0�u�R�n�8�No�����˄���4I�V�~��Qj8�N��-K$�ݪV�o$I ���]��mj�&	�����yiH�Q��E*�j8ȢN-Ŕ���m�s����i��p=��q���8!���Q��Ny�v��s6w�Ar?�Q�WϜ��  �C D*�))jM��$0 ��8 ��Çq2��!Ĝ"V�a�!�N�c���]��9 ��M������۟=��u�;`�wn�BOt��+l�ͺ[�@Ůp.徕�e	EҀ�)�`��4g�zI����'�ٻl��E����D��I6o6 C�2堥�0T�kލ�`���(Q&�Z�X��cʇ��w15�V]U4�Qݒs��&� d�^/�#���cv����C%8��I���"$������N�ݖM]��3�͡���Nhk���c�J\E@l4��;�����Q!E� �h���Ѹ�.�<�e�Q�m�;��8y{����݁����r��~6p�G�?2��h���Ѹ[�M"j4��5dž�n�'����';�?���	^��?~9����?��"\r�UڈGm(ۻ'�͡K��H
���HR�� �q3S�W����S� /������5W����Ⱦ��~���4�*���b��?�Q7R�T$�NATO��>�qۋJN�����0M�c6Yh�aAh�뮷�3��ݜ�?/�T6) J.p����s�}L~�I�w,򺾷��4�IФA�fh�$���=G��w!^n'�(�)J��A�P���B���̼H���{,c��h��0hQ��U]  �B�S����]���m:�}�~_�.�I�]��%��d{G�<,�d�j�}��E�
bJ��!��$�t��$���Ci}����'3#L��<�^�ֶ BrGf�ۺ
�D�6���۳+Ҝ��s�k��=��	�y�#�4�ؒp�j8Ѩ�aAD��&m�}�h����D��o�j�f���K����wH�n��ɦ�!2aLԌ6A2� ƽ�U�$w�h뱉�����ֱ����q/�7j��ae�*����D��wG��㌀�pВO��J$���I&����>�n�4�#�3��5�r%p��D�C6�}�[h��Mj�7��+�[�m�3!� $��A�'}��D�������Dߞb�}��[m�!wT�]���B]�h��Ι'@If�>J��̆g�w���?~�!@���ݶڝ������5L:)���d�띊R����M�j�KU���d�����']I)�zN���خ�S*�-؜����Ob��9���Ԝv4B�����
��%�u�;\�$��bػBV3��	� p��������a,�ZQ:J��Q(Uor�Ov��{$�#ֆexP3�Iq��3�� @b+��~��D�f��s�^Hf��pF���q�u
d�f%�	3	����#��P�M��4�1w�Zh�k�u�&�50:��D�	�r �{љ_�%�͉A'��6m��\I� G��>ӧ�Z�jbJT�a�*�K�y�A5�<�My�ܔ��љ}����5��J��(7��.|	��+]ι$���Rz���r�F�p2Q�7y��-Ƅm�l��d�D�Tʥ�vހ\�5˞�NJ���K�L�h�<< � }�ްO��$��������7v�S�EwbA55G,FH�Xdzs�_'~!�6����(��l��d�G�5R<�ʖ�a���3"���H�)����Kv�Ls׵�ͅ����b���D���-k?�f(.�G����H_�ʢO���z�n���H �	�� H�I#-�)%X����*]s=�pҰ����Z*�kM�}�e"w�2m���I���Ji_����nލ�7)ӄ�$�i/o���1_|�ג�������d�D��ֶڊ��2��m9�W�V%D�I	!��E��5�'�q����bɃ���[�ei�H��~h&�r��]ĄpHl�mf��8.�|����y��b�m;Vo�����f�ky���H�2� ��'�{���W~}�ٜ-��,�~�������DYn~�a��us�^έf�~�����˔^�q��y޸���d p#�p�i�����pd��sv��\�u���9����R���>؄� �)�u���I��q;L�w�w�n#�� �"j�ӕ�A�'��(������s��  �w{�����o�����{$h��!�˧Tq*�e~�^���sU����k�"~��@��<��H���%CL�T�uM����1��c}?=p��dtqj�;)��D�H0�A���M����m/b�T���ݓ��mB���qQq��	�'Qbݵۥ������㒅�7�y��G)��/~����W^��vI�յ�F��4�R�]��+��uI��w���Fdo��J���L���B��Dc�GU"UE�W���>:���~8q�>:u����c�1�M(QAR2(f�̧Y��,KĔ01�#�������!A*IŔ�(�@�$(01��	� �1Jʰ#��]�����<����e�����f���M�%�5
P%"�$��f�&��m2ob�O��g4�{����̰L��AL�]��^H�ۿ����Ti!�#AG"$�[W��W!�^�v�v� G+ٚ��J�ͬ�&��C���a�j)n��{i�dq�I03!
@�)���ci�uB
�M��ݶOw=�����G�_��Q���}��=�m��&�N�hU>��k�$����#��?~���_}ÑW]���*D �� �y�}�~6�2��K��S-EQ#oV�$q{�&Y��Y�˴�љH�R^�KJ'DUD�U�8�`����ʨC �� �|F�,�{^�2�/�Fe3�� �FI��Z󬷞�3Q�ެ�x%P]�Q9�,��b.V5�P��p�:�,�1\n�
I�/a��ls�F�cP���rh3�Tc�z�pu�{����d�m�#u�Ƃ�,%`����5\�<[��K��v�a�SA���p`��5��3�Ѻp(Z�����l�H�$��6��?�������e�.��3��<�\k35�Y�kV��O�<)d����� ���d��~����տP�I���R9�x�bBU�^� ;�7\�U<v��&�HS�=�}��ƒ�M�^H�i�뀚�Ua��ÇQ-AuRZ�]dn��>����
����(�*�0//�}����^g�~�
���{6���pkQ��$���AD��{uߛ��3��"������^��$��fP>� �3�:�,(�SD����e~�ڢOq��g�p�O8^�֓H�N��@�j��I�P�D���6�'��8�w��"��Ȅ�[�/`α�7n�X1A����6�6���&��ܣіR�EBS���s���ۏ�Ć_sOj����P��Q�������n��BHhml4,X��J6a`�x� XA��-��d��:ib��`�&�jL�����2+-F4D�1)4J��9n���b�Pj]h֐"$2F֍�X4�kT��GF���p���c�as2�JJ�ǡ)��}ۻ��(q
� ֜-8��p�p���85�1h�b5���IW#�� 8=��Ҩ��W��:�;�Lw�D^%B)EEi�RF)��8����(a�q;\�Y+jff{��7�p�� �c1a깱ڂ�[V�����ԫ�<=qh閻F���(N�jKTeM��GM<S�,����E�n+��F�pe �m��	��h�mŻ
�;q�,��rfʴv9�e��p���K�Rd,\ږ k�<n6A�:��d��[�2nq�� aҁ��0S�0�66�AW�k�&�\I�@�e�U9���6$�<\���+�+NR�8Ok�'��h�tq�yK��nN�Wr��tU��;�kV1N����+un�k`�m��ema���wm��g)=5%b3lzěr�ڏFRN"�t��ݹ�6�ݕ^gXV�}m浥sb��'z�j <@�zѾ��������<�X)�}��!�T��O�'H ;�TA�iA��
 ��Z �h�Ji�B��V�\��9�{�^M7v�wg�ܐ�.y�����s����ٸ��k�L��
�L8��f8wc�E�f�6��F�v~�?+���7%FSH"Sj3��2J��˽'5�$�Ù,�k�w�s�p�8Af���v���~�a��'*��vO^L.�4z�x��;��7���ps�y��k�ۆUM82�9mD�$޸?J%��l���[���@��~��,ơq��'�`4d����8"����~��������D�]�:'71jj������N��'=�B�&���A�̌8A�=��b�ˇ�7YY"L���}��)}�ͶG�-E�m���8���'\��������Ew�����KNl�G{qfI5�ܪ$決)��niA(����r���W^fo<���\�7�P��D���kJ�"y=���C�J���h��}o�|j�8��tH���.)'(�#rHK��[l��歴x|�ͦ	���D��F�fCi�e�qvN�OuQ ���v�K��*���� �7b,��Tr�&!�*$�﵊$��6�I�Q$���#,�)!�jd��1�#1|/����*$��f�'��y,�2�C8��W�SF�ߝvz�ȝ�����<�}�v�F�+]�L�"obߺ -}�G��#t��E81%�%�	��o�^U}��l�ȍ2I=�͉�{�v��;����r��]QP˲}�o�����W�^c)-21)
� (`��v��n��>�Ϯ�w�����]�Zs"&	E�-�"A?.�Ι �k�2Y7ݼ�'��,��!%�7������E�aPJ��=:4��;�pp�ؠ��{\<�"p&�05���]������m2z�5�k<|�/n��L��g��y�\�ຶ}����6v�"�q�I5y9� <�Om�y,�qoͷ�K�!�qݐH�d�_���=�ݖO���Mz����r��s�������b�P1Q�E�d����Gh��lh��nV�'=�M{�6���uUv�sD����A�;8w�d�ߨQ'�n0�}]�������$�F#�Ĕ�`��2CV��u���PR���J=b��ֻ%q��t3 ���F�՞�(��U�U���]��]����]�f��ȕw=��h�q>ç�>vwB�%�Pzy.�qHCx��	l�fx`�8��������O���.6I��L�(��dͶJ�V\�ċ,�����e������#%�qn�h�w1��.�X��"�$���8H���j�D;�ۅ>+� �*?ǿ;�<{��u_}��}�Oۯ�D�r�I'˧�,�^^Uӄ�֣�RR��q��5.�$�Vm| `[/3�߹��߾��U]���Cg3a�r�nVI�hP-c�V�x�Y�i^�m���ñ����"SJ`�g�`ϸ� �� �(\?s����j�~���W]�m2ۣu��L���Q���cM�
�K��i��0$�IC�s�93��.�+M�ٓ:����u�$nk��}���=sa������K�3��H��T��B	g���)� (�
�%����)B1����gY�(�ַ���Q2L\ͺ9����)�vE���v�K�0n�.DX�fݪ�p��)��[�sٸy6���*ݼ޵����~R���j
B�H�)�J
�
B��"��hJ()j��bB���A$BP*if�T�) ��VJ����T�)�	���B��)fhJ���"��������)
%)
�VJH�h)i�*fhJB�B+}p�03�4OYG���"���e�'	���X$�ݛ�O�"��p0:I��N��'��i]��t�%�=�3hpp� �	"���
�o.�~�����cvY4��K#��ڂ��q!8*L�h�$�s'2Fy��]�>oٰ ��vrQ��V�	�NR3)�fA<�>��+,�6���:������W^������8s>�ג�a�$��-�V��`��o�H�,��	�R��� +���n�]����ۄr�7Eor3i�~xrQ�Vf#�4����~?>�/4k%�X���T�$����ɛl4�����D�*�d_Vd�5�d�#���s7}w�g�,3j��?�J�<E0^s�=�$/μ������$�]��:�GףB���S�j]"MW����k��$�n��M�vv�>��E�a0�ne]��+'�^�}(��1��	�y��'��U���0���W-���vO}��|o��H��u-�������hC"d 5}��XI���������ě�9E9߀��У�q�v7=pT��9����n�gi�da�	5}�M)v���#����\�*�ڱJ9vOu��  �u��f}��I��ʢE�����Q�!3P6Z.���m
$�u�[21Y1V è#�ҙ��fc� 1Ѷ�!��$d��,����Fd@�M!AT%E$I1TA�M��D16>z�H ��}��|綉��4�>���"RK���v����~���5�۸ͦN[�S�tps�rߩ��F6�Ҕ�CJ
aQ �~ͻ�|�ݻg�^�\�Ջ����MqE p����<7u��ܠi}~�6�;���m�l�r�z%R��F�1�c��#*"�FHk�'ٳ�$�Y��I5ly��w�O�!�Ђn��AeCr%ʂ��Q
$�vǳ+x ��LO~R��Iwٿ]�׶�f�V�-�!.�U�qt��y��Rw5��'�ɦ�ĺ����cƣe]�ӷ2Y%^z�z�/�!�D�XܦG���P�!H�	)���޵�:�l֧�F����3=��$�(�e���m=�¶8�jA�:�N�����xpm���aS�+��}A@�-��a�+;�{��U��kg� K6QZ�a	�!7c��Y�\.�C��ӳ{���k5Y��d��!���5�i�{�a�aq�����`�)vI�<�D��ƊTn�q�(H�6�(��M�Ka�d�H_}�������H����i.��N�c�RR�"yG����r�=v��Y�5'I$կ\	�[�RI�}�9���;!f�x`S��*)���q]���h \0U�f�'��T�k��f{�@�p6���MG�� �v��d�D�x����c�|7J[�ƁV�R6�;����-��F�7�L4	;�C�p�i͆&
r��H0�
Q&��0׶?��{����)��//G��h�9')��h�5	��I^f�Ɖ>�nݓ�}�M/ٻƌF2��_tt O8?]��~����Z�Y�V�kP8㠚Ex5��Ӹœ9y��s�^C����������5mہ����]1!�#��V
ΆO��w��۽�{�%�L�o�su�c����q�ne�����D���m+
;�}l�����#��Z�������Qe� ���̭�T��k5�&��2P&��D��qj���х��'�٦�H�����c�O�&���{Ƙ��M2����՞��D�©wޛ��m�eV�'|��TI:7Q�;�RQ�	ܚh� R�P�#�%�
�3R"l�#H�Ԅ"@ ��$M���nmZ$�S�|:�cH��% =���~u؝���,�Ґ����r*eĳ��d�D�ˌ;H��fD�{��TM�n�4jZm
v�7g��߹�#�(��!wv{�s�}Q�Ȥo���7�ȯ<�~ܯ�����������18Z��)&�@�$��Wrɮ�w/��r�j� �;(�p�8�֭o}u���:ٮ�u���"%Tݩ�H$���;/6/%LW�6] Ex��I������J!(�w�7m��:?��gnO�o=��<ݍi ۜ@@�B��A�c׻�I&�e�&���{�X�$�%�Wm���$���*HXD4{�� )ثJ�Ć���Dҵo%|�����u��#6����S��MQ��ꉿza�M祙^L��FU0Os2D��'D(qQ
h)	����ɯ{0Ub����$WL��쥝y�~#�<���z�Ө�y�w��L7�1�,���Ҳ�.�z���iIL�;��$�Uk7��|��kf�kznw�j`�I�j��@��5�+�ف�Y��q�m{��}\{����{�n����f��Fm�5�5�֝kr*L��L���M$�1�CX���)(�XD��Qc
���r�2OxpZ �5m,p1L��t ) ��`H;�������U�PZSr�Y���cd�R	@R��-qy�vTwlQ�jF
]^C����4��18���$!Q�g��v5�us^,��j銴rx�P���ë�
�L�y��Vĵ-\<�Wa�^�û�k��`W��q2�Qi�1�n��DD��<��L@p��Z�h��ԽZhS���ڸ�-@��;U��[β�k���Ab�OJN��F66�@`ì�:��A5;�=��ti�����V9ۓ�F�"l�tp0�P��[�Rr��v�U�e��bR��6�k��y��CC��u]E̕G��u9�ug�cb�M�4U�b��R�k�G'$��Ƅ�7#���֝ �Wt��x�E�r׳�N6P�Y���<r<tRӚ�+Ƿf.9u���l\����ױ$�	�Ml����2aӞ�+�vaK��m]q�N��,�]r=Y��C�!��|��ݶ�cR)Js�`�(.�3ٰ����3@ �t9��أ*qę�WH����&PU�tY\%�vM;#3�%<77�(�8R�n�]&�b�x�ONI�e2�X�wi�.qzC��(�$WlDJ'/�:�{.�R��Ni�������{2F���k�=��U[[��tsۮ��l��l�*���k��"۱mgX%���)F1��& ��灼�\���8�$�aqT�^�D���)�s��v�k��a��uH =�ҡ� u�}�o�ZG�� R��� C�����m"	���G���k
��R��"L�D�[��v�q��d�ra�z�9��2/N��h�lӻr\,��}��(����I�R`�b�cN0�L�0�\�H&&�`��ܶOW���7�ݻ'}����U}}���w�y��ۯh8���%Q${|��>��TI�̭�9�I=śWf%��pH�@#�۲l�ܼ���ps��^íu)�7e�{��?r#��[�HdUNp�R&eQ=���vO�c�h��#���D�y��#��t�\h��2���D�Kسe���(W�D����;7�A$@��h��R%LƢ�<�9��څ]��*ݓa���W	�ƀ��su���@�Xt��фz�k�v�/Z�R�A���Z�]��Lv����C��H���*%����o�c�\���C����H��� 
��m�zF��(���	Tj�&�2Q�իD���Э�u��x$���	�\��[���zf�'}�M���Y�(.�S.�vڍ �f�Q4�fC��B`��;D��c�D�3�On�h��/=���س��6�4f*\C��*'�}�9Z#���cvY'��(�H�b�m�"�a�m�v�mXuD�)$�꼗��G޷��;�ͪ'�p�22S��i����|��`�D���(��E�3�{V��;�+Q��Pl��#D��Y�;��T%$��wc߀��d1s8��0�����jB��ۿoY9�U"	�VmH�O����NS����.p�B8��7~�W���;0�Nz瓴��2�ɺϢ��ݷ<��%ɴh�<���X�.8z���G����a�ā���q� � � ���;�-��v���b��?��z��1�$�sv��{�{H��A�pd�ri�|>�W�n\R˸��j� �V���̔	'��Bo=7n@ \�Hk�4���IRq�M�f�$���%�s7�'�{&�H�Vn�DEѶ��]:RQ�|���F�[�V�Y ��v����G��c�f4.����*'W����}�����;���f&�u<퀠����)%��gspn�M��(�{ՙv!����� P�B�4�N�Dr9�꼆n������F�$�\�0On�N�W �}��R�w�e�iTt"�MЄ���+D��6*�9�A�UJI>�Fm2s�gm���-��,T�$��7e�����&sv|h�����'�/�".H㤜2����%Z�4��1�!�M_�R1.�d�{�X�$�A˒�݊�$�'}�M%������P��N5�:�`��x��m��P�u��M��D��Y�oi��.���"i�u_q�]T7:�ͷ�CiB\�)D��A����H����Ü s��-cvC:0h��DULS2(&� �/"ts�����ڸG^F�$�v�)��������5D�"LJ�'��ݶW�{��]�~�)J�k^��
t��f�`l�Iw`d�C�i��&��L��U��3%��g�J$���^ɝ�g>З�T�Sr�"ӍID����$���H�7���Kh��J̸�r%�Q���͏F��̛��N��4Nn��QP6͙W� �v��xß~,1���5��3~��?[�6Q7�̪4�����@i�}��Q�^��p(�8�E:q3P���v	>ܚM�6U$O{�($���I�Ɗ����BHe�>��͔�f�$�dH��ٺm����c�:uT *��O���8��[�,����D��,�'���� �ADH� H����}�ί�߮_�4\dƐ�t�����2���Vv��]qZ]��U+��OgE`93!��u�l�v�Di���v��)�r��p����'Z���"m�	k���D,=���\8x�G���\�����ˁ�����08>���T����gr+w��wd��vP$�5�N����!�AA�@�y���;�b܄�ϙ��WVM4O|=�8#�u(����w����H��upd�c����lf�i;�x��j���A�}��K9��ߢ�l���GvI�ɦ��'b͖	7{�$���2� �DX�Mp�D�	��<h��1� pķ�3m�=�uI7��L�iU7��DU�X��"{�ͻ$�d�D�%Ջ*gؒg$�ʧ(�]��I�}7m����:������Wn*�C��F�`Ȕ�U��d��qQE̜�G�}�X,�Դ���8�� �y��@�63f
 A- bF�{�=�����g��s��7"��oi/!V�gj�n�c�q���]�p`��t�d�=r��;cD;��ѴQp� �S��
��G06�����W۷�� [�q2׿}C����y�A).��$���Q7켪'�9�yƓ��eF(�{ջ��l2ske���f�'1����/yf�Q�ܨ���teV$ob4ɔ�e���n�ݖNw&�&�P̈&]8�(� r��y{��$�dI$��1L��.ڋ���	��#p]:Ҩ$ݒ}�3i�~b�	���������՜mU��*&�q>(b�xo�d�a�I����>��F'T.���5h58T8�a���p��D��{ݘh��}疉9��s��{�(��{M�%�U�!�UZ�ʫ�*�u�s���c��'}���In���d�7jEޕ��R��I�ҢA��ݶ�=�3U$��h��s�)~�kZN"\�%[wʡ����$�M�12ѥ�w,���U�Ah�R�R�` �U�z��4��|������54\�{b ���Y-�5$�S��=�o��A�dշ	L�3DB9-� T�Er��b�m�~��q�N�m����d���)3ْ7��{m�|<���(�2\8m�"`�wצ�R7ln�d��ݖ|��r���8�G�z�&j�øb�K��|��A����F�dNN  �I�v�	�0bmP��`��&���Hs�5^��k|俥��̟����e�%Rq�`��I��d��]����l�߽Y��=�!n����iUBU�vZ�L;H���ئC}� C.#5�<�m�z�q%�C�������	�c6Y5܋2M��7�)I��b.�l\��(��ٌ"�F#��쓛��։�n����{D�A�)���aq���n��DA��}�x�x8����O}q�I�w3*��9Ϲ� x88�|p�7.c�XJI�$����Y=]��$�ޅyPN{v�㙛E�h]�-��EVI�lXY=�3E�}�]m�e*�܉(��Bz��;5��Ƹ���Mkƨ���i*�^D��t��f�[\���N^��(��p[�3v�"�4T���q�M����Wx�x�Q��n��\�<�l[��-��ld㞺�ڎ2�A8`qD ��]� �� s����L��P�$��Jt�d�XG�n��'��a[섂��-�*Ni��!����[7���t0J�\��R]�Ĕ��^P=i����}\K�<��v�:6�
H�����
$��Q&���"��v���;D�(�DЎ&�M���9��8 igװ6Q>���o�r!��jf6Wz��l[�4m�fl�N��v��pp��>4I��ϥ�g3P� q)��!�fB3���>�� �����9��I$�+�g��\��r��Ũ�%:ePH4��Ou��dI#D4;�vK�"���x��^�㬂�F����"O��#�՛.7���-1EJ�+���eh��GV���U��j�w�q�u���E#��CA���ME��<�4'1�������`���B�C	Bq0Ɔ5c��&f$864ZMf�ǼF����|l4Y�f2�Z��Dw�Nb`��8YI!��G���d�%reݖfF,G�rs��#7bm�xAu�E0�A��E�	d�2�HZ(Z%	�VH�2C$bA&eed��(��R�JG��	@@IBQ+,�"F3�C��Y���7�J4[�5�Y��F$����n�h5�� ��E��z��y���N�A��"	b ��9Q��Г2Kk�4*y	�ܠ�#[�Н���b��<�����@�)@JF<Ǯ�zAI�9�q��A-U��A$�!H]Z��������(T
���):<�:>k�#I�@"�m�ѵ5;V��B���Tn����Av�:�n���[����nw%�*낺,AT�\L�U�t�vS��U�������.�n.��P�ט����EDQ#Pk�R�FP��.��9귷91�F�]X��Ÿ�r[���Z��v��;8G�����a��E�(Qt� ������2'gXy�,�[�u�S��8�4���97d*v�j��Y4�;cC�SOKg �{Z���zl�l�v�ڵG���@Z����Х�砻s̜:9��tኸ�հ��3���ծ���]���vS��tvӻ7!�tXtXS�	r6�g2�l����p� ���9�!�ɹE29,���I��0< Z�(f�"w����T��E�<ت�.�H �Y�� x9��[�5L�Z4���0�qF��7U���Cш�Ю�3�bc~��w��j����X��e�0���)6�Z#C.�Cs0+�]�� 9^5ʦ���4�B����d�F\D�i��ڲNk�Yh��@�@|Q7lf�>����K�U4�պP��Q^�6�7�ͻ$��F��v��� �b��-9�"	��ܦ�v�j�K7v��DW|���}0�%�N։�ԫ*㲃d��N��{P�~͔I��h�i.���;�a��FUGUM)M�$�v�H��V�Qq�؉<�O0��cXv�������'��۲N{&�&�pls��܋�p�m�Y����q�ɂ��@Ձt)]$�6|h�.㛻�M�3~��I����}��E8d��S�-)D�w��}�6�H� L `eU�{$u��D�y���������H���3~�sJN"\�$ �#wd��M.��=�ʦ	�$߲n�#ט��j��lHEL��]�[�^D�$���K�:�gL����h�!�n�� ����
�CS9�*F	9��Y�
Ӵ�W8R�E�!f�o�kĝܚh�Iu{i�X�8���p��2��@�!&9����$�7웶���ݠ�7��-�d�D�}�7�&n��p�,�l�=͚kH�~�
�8�}���sl_�/h?1�.I%7R�eG�Kyߙ��u���~�]'ǀb��)�����9�g����Lu��2����A�EC,U*&��P�G8�^oEO��;H��@�&�;���w7�MZ�nf9�4SU*�'�ly�)/�T���DE�v�<r�By����(^	�@�+o7D�O|�%�K��,���	�ᢷ��Y��� e��e0K����1�)UP�g�N�l�R� �ջY}�e�&��mm�p���IӧD�.D�=��D�9����|��f��i��)�ɴY���j��#�'������ʣ���^Zwe�un�=��Hd�e���b�#߲�m���2������Z�+�J������t��-;��K��)���,�Z���)m�:��Օ�np�������e�LzM-t@j�]�\&c��"����3�k&��&�v(�{nB�����@�2�	�;g��d]��@��l���[��]<��ҏ����w�߾�{��F s���ԣ�#U���j�×R\���M5ԏ�s�����3���
NDYn:���s�w���^�����[��`�+>�d��nU}�r	`É�gR3��;�܋�p�G74Y�]0�� ��ݖH�ݹI��NX�'-��>�
���ʺR*m�,��xv����ݶN{f�$����籹	q�fI�\�Բj�1�z��K;^.՟S'��D�}��"1�5.Ӊ�*���vrQ9۷(�'�~���s����sj�����m�*'��I�T�e{�x+��W�d�I�4E��M��CM$�	p����#td��ݒk�w]��,ѩB�tn��Z,��( 0���Z�r ���a�6drl�T�Ԓ�ے{j�.{�'-O0�e�����Z�����t\zyǅA%xb��&��s�f��|�}8�{�w{ξ���>�77�U�hE���f�$���ݒs^�ɼ�Т{�<�Ƒi�N�4��&���ΠO}�2WR=�ȒM/\�� �KX7tD4�RtUP��������$�*׳*5/^ƙ$�כB��b�LK1 ��Sq2M_�D�ݏZ�A��'#��$l����[��	AD74I�y!�����������9zv1ڙ��AF�FD]�{7̏���j��ȟJÆ�XUTA�����Wg�]{b۵k�����r�I�g2Y5~�I�_�I"����9q:�B+6����|�7���WO�H��!p0#[E�L�}TP����_��(����ɼ�ϭ��������!("�A$ݬ/%�]��;� K�y�D�Vw�v��Ѻb��u%X<P%s�5PԀ;�km�d���ֽ�R�ы[GRP*A� �y�w���L Vv�1�� ]������i�'	�]��ҍ�=���a�o��N8�f��6�2,R `eȀ�ʄ��!ˉw��Xw�D��A���_�Wk�ݽ�F�IQ�)��h��(fQ&������ki�o#s��|ޝ�����b�\l]�5d�|�\�����]k����U�1�ɡ#�GC�B#�&�C HNiTHM� @��J	y�o���  s��k��D��A�����n�r)Ã%B���x�{D�����&�{n���so�7�t�b�Yn�n��L`ݒO|��"h����B��ha���^6�E�ڐȞ�sJ�'��ƨ�o�3m���4 ��ο��_���gJY�]p# ��P)d�{TR$wތ�A�w2��s��]��`l��Y�9RI����������8�W��'/g�@�|s�n�f(d2qѕ	N�\rI��nS&׳���>ȁ��+���@�}>X�����4�N��#� �D�ջL�~~�D��`��U��⑤=]qg��7\OW�N��],�u.vx�P���{/;\�{���
p�{+�y�56J��Ig���m�)����'i��9�Ƥ�,#R���U[Z�)ჶ�n0���h�kZޭf��N��TL��7��-��;	`�*�B�4�q:	�����w�n>��ɫ�pj$1'd@�e��Ӥ��&�N/f�'�s8��Mӫ�%�a2C �4h�mL� c1��
CUj��d� ����Q��6� �U�g-c�&"E(�"�2�o=3�ؒ̚j�'�o�n�fD�W㻨��FQ��N�*����u�$��|9,�{�eJ�̼�$���٢�(Ҥ	�I�Y�ɼc�N�W�ʣK]�i�G�o��������uH�^��[�(�(�5H�#���;��? wkc�<��5��s �Vre�W��2�vȸ	�@ӏ9�Kg��(���7&1Q�s����{\�޿���������N��=F@�ubJ۲ˮ�{�{K�A�b��d1D��R�N\8�����z�u%g��"4tЪAR�H�"�P���%{�l�����&�fS$��g7tHӂӅ(�b��'�p�J'��a�I��ěK��YU� ���_7U)�@�Mʢ{�>4I��e�����G�~�h�{��I�̗i�F�I"Ub�Qq'v^*w�{�$ݻ;H�[�k����8d�$��fQ'�ٛ.n�Zf�D$ .1$e���װ& �ӣ��?�����O}��O��2��f���Y�j��V�2��S��ޮ�%��a�g��Ԍŷ%�f>�����T1�����BG4�Ÿ���5 K�X	!��a���Y��C�E{ˬ���'��/)��㘧G8탣F�P�*&E����H��>�M�f���i�I7�Ve���G��*L�i��~�����&��hU$'k%���=�f�p �U�,STn���ݦO��}��N���թ�7qlҞ &�$&D�0$E���Ϗ�>�L4ZW�L�p�ױ&�������Ce�l�>���a�[�	��Lu	�n۾܉$ҳ�Mv��H�{2C�r�GT�7q*X1��K_�l�n3��۲Ny�څ�~�go��ˎ�n�#3���-C��l�',�nS'��,�����z��V�:���[�}�]�s��p���_��W����u� ��`�3Ia��������5�=#3[�:�0�Fke�Y���q�F��C#�W'@���Ma�l��SI���y�$vf�K��$��Ƴ������}��s7�ڴc�-U!���<-���ґi-��qOJ����_�R��rZ�F�$Wc����*��nv��y�x��ΎV�YP�)�b:3�d5ͭ���V]E*�[n�0�t]QHv���l�n��<�#���n9F��H�Z�Znh��I�cs�N�;Z��n���/ˢ��v����a��9+��-�V��r ::cu]!�[��\��<�gs�%�7��"�ʓ�gn�Q�>B�qҭ�5�[����Z��tC� �X�Q8R^�Б[u��܊OV�0`��6)wq�/v`-�ɸ��E��-U u��������":��
��G��X,5���I�Om�\ON�96��A��J�N7�����K��q�z����3�Z\ˍ�T�>��θ�i�h��j0�n��!q�v-�1���E�6yI�s��\ۘn��@�s�(I��MQ<��6S���m�<m&�<��u�nZ��<8��G@:��6~��z�'e���ie��l��<���7���=�����r.D��b���Q��Iz^�ZQ�
����]����v�r03�֚N"wlB[r���n1�Z
x�̓v��ַf�Zֵ�����)��(�6 ��(��TC�k�_4�.�O��^�u���pG�0����:�JJ��F*�yA�]v����������D�,82��tn��e;j�c��nТN�Ŵ�,Y�l�fmݒO��jB�6Ხ�T���dH��"��a2:9��q�IqR.
��P2Rp�����M�m�{�i�ǻ!N�P�O����A��یu�q�2� u��O�iƎ�{܌�p���H�DV|2C=��P�\!�7HJ6
){�ݮ�I�xrQ3^�H�]ř������X7M�N�7�'���L���OV�d�L�l��F�X�J���$�N
 �g6Y6��J ׽�TM�o�u%~9�69O��N_"kd��O2�Rp�5����a�`nkd��1���]r���s��ɶf��O]��\8l�	c0n��c1Q^6<��ݹ�mط\��p�fb9]�)�P�1��䈸!�!6[j�y�����H�O��ڄ�:��XA�5V��d�V��=�����y�9�N�8���6�q0�"F��]�3~�	�1�L�o�6@���)	��F���
`�67����t��sr?y���ͻ��ٴ(���2qg�V�����#�n��i�U��^j��� ��d���DseY輧�����2�B	BJRR�R^݉$ҿ[��%z�7�d�{#MW���P$�ҥJ�*��N�ݦMﶶ�K=3Ut��i�,<�G�H�N�y�6�~���&4e[y�v][Y�dƋ��� �P�0�e���9�y(�W�r	�s/D��/���-������xADS�&&�x:�JWg�_����q��D�"h��4��YM���-�<`�/'0��*'F��\n�$��*���u�#�-��r��d睋�k;Җ����w{�����z>.���b�Eg�B�Z� ��h�S��20�'�َI'�^���{w���j$���"ǝ�0�{܁���(����{�-d�5�����w*2��`Ў�|X��@���l�����$��k�l�2�IM���Bj/ލ���y�� �����/{�2�W��2��K�*�1P0��>��#}�w�;��ݻV,g:2F`!����S$D�0E]��y���D���͗�n�F)I>���'5��p��]���t݋�Yz�}�n�	�z/ts��N��Q(�����*G.��ՠ`��9������@(B�
�(z`��־�X�N��{P�}׵>�8y�[GSr%L��fCR	���ڧ�z�0���9�kgv}(�s��ы��ڜq�Z몲�ƨ���h�9��i]�2o.�'���qw77�M�:�m�&fZ&DnQ �u�+Hwl��c͈Ad�
&(�M�h���\*$�FC�«��u~�۳Լ�i�w}�%���jY��w	/����^^��U��)��N$}���#���@���4�>9��b(��(�$��"o>��� �� .�=�%����Q3�~�k9�״^�pa�T�qD��0�Q&�cO�4������޵��U��k��z�߿n�>ܙ���n�D�!N��((�Qpo׻�$�����U{����⣈�=[u�t��/z����"~�#}�e�uV�W.R�t��m���My��N�&�4���ͦo�1C!p�J?���.]*B��V�\ŵi^*$�.3i�:�s�L>�3���ps�g\�Pm#�ub,|
�j�ӆ]��y�tpp����D�e�R7�nP�{�!,���U)�b)D�k�I��J$�=m�z�wh}�sC-�.T���d2�N{`�@��mM�A�<�D���U@=���۝�Jnn���̓��oj�:�M�)������z%t=c�kn�Ju^W,F��z���*��.,G[ZgM��k��M���AP7c��']n|�3�L�r�Yl����$3sH�(dM�p��ּU^a#�X�&'*��#\p��s��n�#�_�>����<K�R0�d�j1�PʆJ��h�I�^�.�+��L�n�`j%-*�l�NE�D~��i9��Cױ��*}���F�tƖG����ܬ3�d��ݶl���Ii��b�+gW}�F�6��("�ٷV�Y��U��׮ʄ����F\�P�Q'��%���a�:��,����e�煇��TҨC4O����2{lfK'����ih ,v2�HG����F��ӒВء$�'36�Zi��볎��C�����]��$�p��^Th�u{)���۲|t�fCAS7H�J�F̌��]�&�+8h�C8���5J��w}���(�����o[Y�ݫ�z���M�1h0��g��2�S�[-�2��׌"�3-ow�ܣ�-��7;����\k��A��=���&�&$��7m�{�nӥ�ڞ��R�j�J�#�ض�/w�om;��(�o1�#��7$qҪBPn�3٦{syU�Myټ�?��U��,��F'��,	l �V�Cvh*+�{�h�d�=1�$��Ne2s3km�n�b*�U�A@�o���JT�D�(��:�|�,�=�h�t�g$�b��N�nݒz�wi�}'�9��o�?�C���8��:
M�T�@�M��M{훶�� 	�}��s�[GSrEJ,�j4�	/{c+����C�@ 㠍��I��k����YH����PA#�%I5D���rH'��%�8:�Ǉ.ݥ���w��bI>:2r5ER��-���I��q�I=��e0On�D�s��%�FX���P7f��}~ն�����N����6ZѮ®�Z%� 1Td{ۙ�����D�;�v���c����R �d��:1B�q�
1�f6�1�R'�����K�fK �}:7��ۢZ�*	�ձ�*ʫ�������A=��>�bˤOW�}I%�ɛl��ѩ�!R��V� ���I�,�fP��l�Rv��o<� ��}� S�z�^o�����g��o[P�cձ'\(ZR��Q
U_�k�6�s����Q��	��%�ϥwF�B��qP)���7����eݫ������ny�yq�a�"��!iE!��=���I���f�]ư�$_O�"��ºmI�I��Bّ �m�$3����E.�'���Nw�k����c�I��n�9��zX1���U�bEH�{��_���[H��ȷ��nk���A��໻Uw

��d�2i�@�뼪w��1��T�w=L�+����uJ�p��B{ߦ�K��6�5�~}�Wz��4��W �qS<����?�vN��Zh瞪�^�x2T$�꺥Z��0�TN��+�íſ���G�([�c,v���֠�I<��(���`����x�GF]��T�Y�BTC�����j��k��mqġ�� !bv�zƕ�������[�6H0���Brwd��Vm2D�)Q�ʂ(\ �L����5Ļ��n-��#���stJ$���h�]�m������)����~}��B`� .륆�0�$��G.�4�]>�d���[��}�e�z��I&�&��B�$�{5�$��ͶI��d��쯖<�X{�J���E�&I>���H�뼇+J��'���L�`��#M8.GN��9.�=̃j4{�<2�Du{1�?s�ە�{�����0J�Ҁ�P6%m-U�U��'�eP��}-6� �L�.A"���rGA�l����/�O��t��K/"I΃�	�����@��89�k>k�������A�L�堸P\"P@ٌ��C`�`Q��<� M�T�͏gihoF����XXc�w��kM��r�Cn��.�/�h!�DQ4�#�A5����)�Z�a��($�$��F��"���Ɔ�=4�����Ҷ��Ț���+{��{��-�)#3Z�p �����d&@P��uhW�4Z�j5 ��2Ջ��b���������!H��G8u~��"/<��J����G�h�����}��?O�� �(çs�j�ݥ���l����`�����T�x)/cr�v�VEm#b鍩ScU��4f*�\�;��Lc�\P������]�'���9�.<���[@�iG��zKʘ6�0�w=J�j	x�,�]�@G��u��i^0+����1�൦�p��'��l�r)VX�B��[��e���[p�-��{\k#�kf`s��cKP*�*m�a�])�G�GK�;OY�w{v���<��T!У�԰���X��s�C��l�ŝT�cIք"v���q�b�,�������(�w����t��E���\U]t..��'aKj�"͗rZ9�l	ڄ��>j\lm�&�U�o�?ټ��!B�~(��x8({��~�XOh�B��A��u�T4���D�T�u!��.u����֫��q��*%r��4��얷)ʺM6����n�wc�L��屯b�r,�9��avUղE��c)�q�
n`\ @s��"�HX�\�IBg��	�)��E�_�$�Ù!�3�yTI��UPO[���s07$q�R�t�A(�{������i�ջ����L4NwV�B\�RY
�*^u�4J$�za�OWO�S'��۲�T���N�(0�RR������	[��y�vٴ��v����aFIn�W`�D��m�$��ߓ�E������8�jn�smq�!�H��q^o���H��dI4��(Q7卣��
��*�m���l�"!!4�03�A�nm٤��4�'�c�L�u�ʠϻ����R+�D�mQ7}KRmn�y� pC�Gv�>��I�mi�Ü���A��l�**�Jrn`���"KJ�M�Lb^���d��i�z=��Z�nr�BLڎ잭9�ɬ�ʢH=ř!���ӛ,���ʕ*�r(�}ϫo���O��N��\Y�.�R���6�j���Q7��'���L�F��YUl�&�Xh��Ƙ��L$$�4�FH��&��Zl�}�fʀ����7�ͻ'HњZE�(��<aCs$��7���}y#E"}{3����f3S���pfF�����&��2HI���B'��̧ޞ0{�x�	`j4z�8��4D�2�iBi��CG�-{���n���v����:rLj�*���f��y��d�}mc�ɮ�Ȓk���xZ`�����2u���'wִeY($˳���U�Ցꛛ�m#)���{0a'��R&��6����{Io��?v7��v�.0�����h�"5����ɼc2�%~�۲I��e��Ye��ٵB�2��'�̑;�l����;�{(�߱Ȑң�=�#�*�����*$�3km��6�m��$��{)�Ù��"r�mU����y֖�n�bI=Zse���Y�v��E�O��0�X �	m߿ϗ�5(�p:�qŹ�,s�Ƌ��]5̓[Es�`��R�ū=�~�_g-��� 
��)�ǩ혠�0y�uػ�Ls%kp�%�g�87n�܄ėT��nɑ`��pu�5�m���8�۪���(��{���Zx�l�<����g�߶ƳG*���*!&�SF�\�$��U�A�q���<�d�$�X�J���L����I5�\�+K�2QﰼzTH:6n|  pP�)���	"0�	J@\ I4��_I>����7癷	=�ةէv����ȄpʧTQi�&I=�^UiD���,���$�w��t}�$i��%�H�j�����˷'@����U�9��0$���nB(�6#�~X�?mz"��MO{�m��ԗ�m3�`OaE�WU޸U:�8����eܴS�D�M"$m� }��Z�
�6Z|����wq��6�6��'9�Ȝti��gu� xz�,%h�!�ѣu�օ�U,qv�u�\-�dFz�،���톹����!��q��3�dT��F9��Oc��-q�u����t�Eg�9����eơ;D߽7M�OsvQ'����7sd���R�@qE21,�j�'<�%�^�ȒO�}nJK����G}����S��Ӂ�H�Y�贯�xf\�^rf�$�۲��'����IU��Z>ݔh�]ܭ�-+[��d�9� �v��>�Z�܄�R3N���tϽ{گ$w�pz�w�6�k�p�(�@�[�!��݌%��G�����ȝ^ӎ�7�1W��i��@���w۝���?wlg=Pq�ZG��Dn	��%{^�Z=��ږq/l�W���w6}v��;�&�2�t[��i��=כ=�xs���r�I&o|Ug��+�u�����;vI�dH�{Ie�B(mݓ5r;��u�$�vn��o���G�"u}��':�q�ȌUR���$�Ծ����T�۲�>�A����0�9�ڶEVj�6�
I�'��m#��s��F�y�mǺ�::f;s;�vQ� ��B�$=�9�ɼy��T�}��ݮ��rYT�����9	-�bb) �$�A��k�%��wޙ��;��(�ַcN�Bڗrꂔ��ɦ�W���x���m M�m3�32u.*m)D��M�v����%�ij���o�C���ck�]w}�W��x�h٩nܶ�wd���D�{�h����w}�vNa:�j*5TZH�0�v2��d��s��m��m������:��ʉHA��j �[�Ճ�O��I��筞�-�\�.����]0��@�Bx�[���:�%������`�gfe���Y� 9˄�2�}���2㎒�6�T����v�>͚hz��]�"�̝�t��c19i�Qi�ٗd��k�D��,��o���N��3{D�lH�S�GQ�$����p~ݺ4kX���w��l��/�9�q����3p��Q&�8R�%���̭�N�<�mD������U�\�v{7����<փ�vQҐ�S�sHn�.��v�HMs�W�H�
E�`�68�D՘�bM��	n�r�l��A�0�ţY�ެ��ެޭj�z�:�'7ǥD��f�qZ�Wd����\j��r9�`!E��CP)$28���ͫD��=�N��m#��adB8eJ����	O��jչ7n�gP=�"�;w��&���kދ:"}�	�GۢF�pY����m�;�>4OW^��d���*��������`�j���]N�,{崉���I��VD�jݠϻ᭗����RQm��d�?9�s�=��'��'�קv��Nf��GT�"��}Ϸ�$��Ⱦ>��n׎z�ܘ.�R\CV9 �
C�8�}���uwS�f�^����}�"��Iq�h{��y��)�۪�F���]6�̢8ⓧ�%"ܝw�,v2']���G�z?�=�s�C�"�`�-c�֮M�p\��e����&�Üe"iPdXp��00�I���r2��'�-��7�L4I��0����.�n��aʪ��6�=^3(�����W�˲h.�kM~��I��?B˓��I�nE�2OVj�)+�M�Ďj͖O}�0�K�J���&C�(Kj�6��K;9[�f�v��=Y�tN>�dg;��R+�Y��*Ļ'�٦�����(���nt��6��F4!��\�78���n['������7��cB��f��o���<�Z#6�c�&q��	�l�]���}�2M�e3~�-=!����nGVI�7d�es�pp��̷�fɤI&����Y�mg��S.e2T��a9���ޤ���)+݃)��B�{�$B�U]�
�$���8��o��%׋�I�=�0M_g�l��)�UUN�S�$��ͬ��}�z	e�"b�@��Vz�<�ܴ�Z&��}�	>�f]�N{^�5y������-m�m�mF�ND�d�ؒ2BXn-u��!';��I�,�d���o<0��p�Q�U&UQ7ܛ6�=�M4I�ӹL�^Ħ��,E�i�qU&��'�3\�uudK���o�4�}��۫V�\�*�| ����D�2a(;"��N!+���g@a0f�ET���Ao�v�mJ�$���Q��4ƪ�1�2K5��Un�|٨s5m���-ZN�s�,�9����Yaba�qtF�]0�YFQN!��f,͎A�cZ`�B���Vl��K��t�����t��͚�%�l!���5�Y�-�����$<6�m:��"=sa��G�: ���o`	�d�
h���&�{;־���;T%�W_Z��aʰ�BO���p���f� #`)6;=N j&����k@U���,�"-&�*5�4���ق#F���I��=��ݱ�Q��4�,�q��n�i�T�1x���H�*�y �e���Pv���S-�M�[�M�j�s�-Җl�=`�7r��$ �y�vy��2]mN�$\�:S5kuX�\�Z��DkƼh-a��5H�ckn(�W	t�;���
��������,5բ�n.�W��k��"ʄ���n��Qf.��8�U�n�/M�p� �hA1�G;��l �\�e0��g������#rd�-��펗޳�gb�.�7TE��]��"m�c`q��ݜ�% ��*j��+BD�<�tp�����Cf����U�X�kc��ێ�6�� ;4�r�Yy�׭-ɐ^��ӊ[X��1ٗq{<i:+`�iw��x��vݷd��8Uq[=�8�-��*3�E��.�Ɲ����B.�qD\�S��v듆�!��M�v)<�0�u�譖82rnn����y%�<�][#��B���sGm���Oj�N�wH�]�4�jR�ݍ�80i�8��1c�]j�xHG�$��]�
؉��U����[<�ۂ栞��4�������w���<T;tJ>"���C��h��G�C�
 �:�=��������S��oZ�Wi������t=�F���4]j�/<�tIպ�&��2�=��4M�p6Z���Ut����O�������m��;���=y&�0���6"R2�BHڐ�w�o�v�E���U���0PG1s�*H�H��tD&r9 F�lC�m�4"1ED��fݒ{�ɂiw�4S'b�w�`-�N+��]&�b;D��gR�W�\�z��"~�z����H��E��6�$��=�����xa����e�'��mTY�^�B$�Z��v%Sn	vL�;��=�fe�w�����v�:1��A:�4Xv�	�c#�B�ț�*JNw�5��
s��7;e��U̷���=���F��[�����:�� We��\�!������d����Sa�І�s��8��KWc����ی�f�7�-�G{^Iy�$�j��~p�
�( ��oz�~�\�|�в!2�CHюC)�s+m.�7q)Lp��=v�n��k�v-(�!�c�ｚ����)~x\G�70H�N�� T����TKhD!���d7 �Kmw�����*��� һZ���q�L:�I�e7L�[�U$���-+^9�d�ޕ����S�,��[Bj��
��-��'���&}k�^괭�,�]��F�=��Pb9� ��h9'|�y[T����$�ǚ���^��{>i���f��
El˲sڨ�uWt�j��4�	��1A�v��A��fF�����������Q����e1*G�i���8'���@7��i$$�+U��6-u�R�OD=]v�Q�<��`㠠=zu��Q��[���Mm�:9�Mq�V�rA:YIt�qFQ� ��b���' F6�i�a)B�M/T&�������D�x�D�v2�s��M�ƙ'�/5BnTE��L���/���l�ދ�dߞ��O}�"�T�Ռ����%0�*)+ܙ����t|������,��{��(ڂ+IС*K�N{f�$��l��^kݞ�g�ݍ$�B�I�*`�'�ݡD�D6Ԉ� �*&�R%�Q*C$d�Ɂ��cB;�����g{	X�Uy�Z{�u.�����'�2w�`�ax�U��}7���"o��$�i�M��f�mr(�9H�mB�o=3nr��:�@��8�)��ׇr�,(.3�g�L���B��Dw:�,��Uv�$�ݓя5Q1{��i}�ps͜ձ��oöOwN��N*��Ɲp�����e2	�����vn]D|���x����۠U�HP���X�O�����&jX�sO�m��7���3�!G�#۞�d�^j�O��r��^Ql�]N�-���q�������(��e�
D�r2�@��7�K�fزOq�͸I����E�M�n��Hm���%է6��|�hQ&���i{d̶|qb1�)H
ID��G<��"O~�Ϸ'l�J̔!h�h(��H"&"Ja���Xdh�&!�RZ`��(����*�!�G9�#]���I�=�b���Ѯ�R�X��M3�D�Q�ͣ��]�^��g�9� ����)i�7K����ö���'>ٛl���+!� �,"��n$�8�n��ۨS�w|7u�{�D��Y���1��}��u�p?v܈km[�-C*	.��fТM��d��ͧ仙WvH�|Jѡ$��1�	��2{�u:� =�f	+s&�lx��c&ts���z�'&�����P�Iհ�3Wsr�����
�̃k�XXCBU:T�U	���ՙ�V>Xwi�z�Uv,{���LQ�@Y�P0	�L��������z�7mi�1��4��U���4-i�U�R���c���d�k��H�Gv^���(������(.e��8�/P�[�u������N�bN�B�T6.ֈ\3�p�w=��8x�)�-۵����Y�ֻi`	i� sw_�	������p*�w�L�_h�c��00��$$��؁F2H�*H�`��)�f-��'��&�}Yh��9��f������u�U�JLbm��{�m"O��"k��ݒz���9�^��+7U�E�����DGrkۄ�XݦNwЯ%��e��7M�ZR�
�7���D�shz�=���l��[5�f�H��FK� ,���.��<ߝ|���ɫc�	T��n����)����H���J����I���:�T�HA2����\Y'd;]��p>�u�$z���l��m
':=��n9r���x)JϨ�8�(y���fo_R��l^t��J�ڜ��E�h���t���6h0���ZY�ItB��0G$ttK���&���8:���dh$T�ی��������+��Am �I�:	m�Ln�\�)�UE,�s��@߽YvK]f�$�Ӻ)�>G�nrJN4�eW�;�[j�=����fJ4I=�8O{��qE���:j��1w3lQ'�ɦ��j؉����9��cI9�L4�]miݦM��@I��e�-w ͦ{�����7R[�b�e^�Nln"^��T�㝭��#Ȁ9��]�=�T��#!����u���B�=連$f㍮E�)Z��J �P��(�-��N �iC�"]ݙ�qbǻN�=];�ɼ���#�!WU)��<�{޺����܀Nw���>Q%G�p@>;��4I;�p�yٙl�t�Q"�T���!HARQ'���D��^�%^�ܶOV�&��f��@��b唢Wgy�p/nH�D��9W�O��ɿz,�5kؓi8e*����.TH�}7m������?�T�.;9�k�a��"�B-�P�JA%@7��^�_�$�4A'ز#��"��ʷUf��≶a�J`D�a��'�s]mx��&��(�����:��@�R"��I��fJ5�6O�ld��{��=�����^,�&ʊ.iLCTK�fi
�\�{~��Q�����5\��y����=L�[��8G�����NØII����;�֏�Ʃ$߽d��p5�S�>+4NyH I���9�ԭ&y&�iY,9�(R\q0T*M�	@�j7�t{�&��kޛ���<Q�2A�ӣ���Vݭ���,�����o�3�M_�(D�o�t��y�Iܲ��*5Jګ�t�8*�E.�Ϣ���绛�gzǴ}��s��3����"���;��P���E�|���ɮ�̈i7j$�T2�{��7|���9�X��Y'�� ����Z&	�0m9w�ΥjHj@��aA�iI�����1O5!ѝs���;���VR����t�p��ƁL8͞=���Q1yQ�q֢\�]��F[� ��};Q��.�c����u��ܝ<p62UT��a��E�Fp +���Nf�5���p�e�*�z��	��u�n�z8cs�O6�MwXB$�p��{�7���͡�����=:�=?'���N��kvs����\�����L#��۰s��=��3$t�0�QC�������9�c��,��lU��y�8���e��b ����S�w۲Mf;"�nv�k�Gv�bJ���L�| ��ۇ���kO�/$h sU�������$Dˆ�E8;���9��T���x��-�Z%3�[M��"[#�����������:��<,�o5���������"���b�������B� ���+����zè�v�� �E;�RDR�P���E"@R�hE)!X�Q �d)RVD@\�#����EYAA��@HDBdUh��h62�4�� B��J
��Dz�JlVQ ���@��F�";�M@*��Ҩ��#��m*w
	���J�H Ҡ�"=`��]�)�FSH����B�2E*�P� ?Ӟ���α�g������U��8889��;��k��'���g=�_��������O������������������Y��<����#�D������~߇������3j�*����n?������*���������AVg�����3�=�hH:?�b�T����o@������?�������*��'��݇�p�O����w���/��w�������������C�������!��?�J"����Q9�W��(� AIRI	Q%�Hd��HFAIFTI	%P%D� �R�R�VI!X$d��IQ$�d�TH$�� �d�YQ VI!D�AH$� BIAHTIFIBTHFIRHTHTI�Q �!THA�Td�	Q&AIP� �	 IT�R �%AI�RDeD�IP�D�X��`%`IB��d%R�	HE��H�%@��RR @��E�� !  	BB` Q%!T����I	��U!!$HB��!)�$BE %����BR$"B$ ��% HB��	JBU%$��HIRP�$% II	BX	HH����VB��$"P�H�&P�RF�@`$$ea&R $!� �"D�	B )J%$ID��E� P�P��d�)�JT �!%P�BQYB� @IB�P� D�$D�	B$Y�% $HB�D%YQ� �%�aXRRQ��@�VHB�B ��%%	�B!XIVT$?��*����(ġ$�B(P
����Ȱ²#��,,��(@�$�(°�+"Ȑ�ʴ�J�Ĩ�
�	B�"�P��J� �,���H�!"H�*H� �(̨ �B
R���)��'[��w�?�����(
��*���S�:��������/��y�x��������������IPEUۼ?k���w������������?����������?w��9�濵PEU�����QH_���?����=�i���������*���Đ���UUEt�k�����pEU�w��v��ᆐ�0��ul�!QO�8�gI�	����\px:TUm����������?��'�ި"�������ծ��py���:��?�����g����}��PEU�������/����!�ܨ"����QO������?��g�B|ư?����3����������������~?�4��G��������x_��>*��>�1����C�?|������ߝ�J
�����_���������K�_� y�����O��O��]����UQ\������?��.���������?���b������1AY&SY��� ��Y�pP��3'� ax� � ���P    �   Ѡ     (w���  @ � P �V� Z44J(R)   U   ( � RB�\   ���U+0Ͼ[g�;ڏ{7ed��.�.�(郜����/NF��-�S���I��Jݮ�i�  ��H��!)(��]�⡷0���[���]�C�m��R6��ir��U2����vƇp�[��C�  �)UQ&6� � ��� ��M-j�٠�he��@PͰ Z��Q2�@�-�K=.� I@ @���%P& ����m�CbƔ� )�6�@�6�M3Qd�
R�΀5K�E]�٠i�$���1������J�F6,
��r���׽۲[�:zކ��{�����=x���\�OOw�����ݫ���zo �P�I�ǝ�x��#���5,�����޺�X�=�+�zK���6�oUs����X��w��:'[�r��  {������x7v����]{7�N��/N���X�O���{r�or�ө�v̬�����w���xJ"�J*<n�T��SC^�x2뼍�c�;�G<��=oPw+�psݣ�ӳv�5����E�x g(�J�6��To,��a��:�)�nK�k�sw�����Jݮ�WQ���w��p =!P��BS8�op����p;s᛹맽ۚ��\]ނ����`��ʽ���y�{��y����^    S�4�J�  �퀪US@�@S�j�e%*   l��6��~�  ?��SmU)T�   D�LRT*mF�0'��_���I	~��O�?�?�_���}�;]����w��P_k���](("����@_�  *�� ���U9�������K�B����܋��7�u��ͅ�)/$՚��џY+�LL��n�!0Ә֝�Br���(�YP�B�@�V�i� �8l*���hHƃU�1���I!�D�@ �0$���"B��BB����ԉ`�,�6B@j$��B�ctp6J�10nU�Iq��N�j�l�XV�o2�z�B��@�����\��Ie%�k2^FA�8K)���,�y�$7!g(����,�e�HW+��#|�
�:Kb�� ,b��#A�V�ԌV�$� ��$�E(K	�t�}N&7��X�
\����w��Mu+�¢Ĕ�c�Q0�6��D¨��d� ����C�U㪽+ap���ƋaAf�m�8f�ٹF��spϥ?G� I� ���|,�[��i*�a�t"���l� ��)	  @��
+	�A�0$X$#H�X@F�u��N^F�>ެ%I	d�ֈX���a�$ۙ�o���.��r��\6d$ JKa�϶hI_f�{�}��R�0��T�Q���b�0��8�l�Ć�R��>�X���k{���Y&;�}ͤH�$��4�%��/ �%�X!�`ȥ�i��s3Uy9��*[G��Q������sfPr��>�O�Xi�E�
�ns�V��N`o He[��l���I�l^��O<*��W���L|Skឤ���p�\3�U�����}�o�C���̆�}��a*�ß}{4rd8U�6�!�j�&�YKq��!z�9���q6�����f]�|bU�l>�d*F�I$HD%<���w
�%a���$cw
4q��l�^�0�������0��J��_E��o�.�4����CNc{y�+�}��xj�z�yVl�Ûŕ�^����j�!��(�3�7��8u^�Ԅ
�B�"P|F�2�[�Cv�PˁXʐ!N���a��h��l�lT�b�:jn�l�d�7TƵ�M� Ec�6�">���r��?m�Z��7C1�y�~ύ?2��ѿ�-�٣��)4}e%�佡�af�WemՕ�ѭ��cT�)ܲ���el(61�
rA���R��Dѩe��[xi�/5��������ݗ7����,�M���||Yye�B�%B�	w�5x��Ұ�"B) ��,H�bT�C���>��Ur��1�1���-~�5>~7���!��!�"@�P^�����m���0��	lJ PF��	C
��Pc	,����Q���������7�@�F\r���{�Q�u��_��l��Vk�{�i:t�F��7L��;�w>�s�'��s�۠�\iɭ���!wf&�2�Q�2������6k!���B$>�E�F�-��ۼ�J14�53{��f���^���߷�8��^���d�p{�{n�ԋ/����gx_5r�p�G�n]��,����D�谀I�@$�P���#�@�Q@#!T$QXP�B2AA �+$B,V*A�ǉ�<$bQf����)C8Eѷ�8=v�M�a���C�IB}��"��>�#�B�Mk|�KI����Wt��͘G�/$~zl��K+ߏ��ϻ2�h F���og7ݛe���l�D>��$�.�aN��jBٕXo>5G�Z;�,ۗ��J�i�v=���c�ô�Z���Y���I0���B���d F����$
�����@�J�ZcL
�9���4�\*�VNrߌ�I �cF$�d$#g57�������1���
 Y)��Y��[	 ��KāE��D��U�@ޒZ�F�T�Ħ�U.�i�$���1�\k���B�M�z�j�a�Q��ݜ�u��DaE� �Bw�C�WB�U�J(%U�m�N�ї�I
�x4����ѩ
�N06�a��HA�!�t�(�A")nH!P�� q�N�Wu��th2I(n��oB��^�q%�����0��FD�Z�.��K&s�ǉ* �1`BU���А(�JR,��V�D-.��r��`
P
PD��� �!h	K(�_��{�3X��-�FY��0�|�-�B�N�B_����� V���7�1:�����J��ӿ�};��Ԍ�s#�'��,H�e�z6p�m	XY��o���n�0�i�=/4o�$81� Y������H�(�A����R�i$���!Va&�M5M}w'ε��.tִ-f����#�'Ƈ�^B�|�� Q�V���T�~��6�*���]�������ݟi���#
�5&onk�g�)��1ӳ�횉 �Y�5{͟S����*�i�����,���u{p��_?`��4�|}�˵����g����Qy�f�_!����L�4l����6���Ia���)��:1B-<���B���Y����A�(�[��.Uٟ=�l"��l*�ZB�0>`��W�����Ӑ��hv��F��'~ㅺ�[����]�eM���R-	`B��RB��y0��$9w;:K�:��{7x]�<�~��hkP��l0�p���2�����,�
-�[>Moa
�Cj��ͧ�%Y���5{��P����l���f�!����[I�Fw�%��� �?<�"T.��4(�,�-�H��E�B݃�A(�A km�(,��4�ݐ&�.�Wc'��>+e�]%J!Q��(0۷l���,l	�.���to����@�
�\#��Ta �
H$ao��U�Q��}�["LHd�������!�6�N�ZZێ���ӱ�bh!hmt��E���,l2�]df����$�̙#����R|�%���E�*��K����ې1� d��5��Ku�[.���-xs�)����?<�G�$,u&����Ϭ�i��%\*��a$!Wy��l��W��N���Bpܫ)A)	 T$��J,�D$��"F�-4�.�5Ӡh�`D%Hن����F�cm���lԁ�FrC��W�[����kufoiW���tܢ�[�a�����U�t��ƣơi�F�4oEU�}㉅����T^M�n0�
��F�$��/8X]�Жj�!�G�$`�2�SP�ې��@B�Uc[����h�1��o���C[tD���i�jPF�CA�$(o!�z��KdB��6`"h�4?�DѳD���`�%Y Ƙh����B�e��7����}D-���50�������q����Y�ޡ��|4j��i�Y�퐢HW�1�s4B�����¬�e���~����3�O��w��fh�Ha$��i.Ҡ@�0m�Bx�!��B�p]�E�H�aG\5|~XU�`@�Q����-`�Ą�$4��!�]����D��b�Z�	��+A�F�,�=!���hQ��B��`U��IG�-l�J�t�s[	60�66 J��)��`PZl�PJBvB2��DH#$B!P+�h!39��iܑ��A*4��)�Q`�
KSrKb�d��~�IdV�݆�Umo��P"Pa
�D��j�
����j�ḣX�-���)\7����@�E�G^�Y����qQ���#���&͐�YL
24��&*�icRFEa
����y��ؓgنpr�	�BQn��6i��M$(��-@�H$U����),�aK)4���`�)�9����!�E�;�af�g�����Svyy2{:ղ��o�*_!�HP\0�L!z���k�������?^kd�9�e�V�)���vV�����A�#�
�b@�� IBB��*����Ь	f�5Y6�$�̹��I�V�g�+QP�@b��w�^�1MI[nU��M�c1�ݱ���P�0��v3�3X�m3L&/��c1��f<�~-�m3</E$��)��f3�Ic2S#�ĒL��,���a�½��at����l����m�g��c4�b���f<�2ws�nrbE�ӱ��n���5��$�b���Wql�Y�>l!��,cס�!�?�Fi�g�7���K^�(�)�,�O���l���Icu�ѧV禞�&m40)8�n��j��&ߧ��,�I�x۳�̷~�vh=�T��ӧv������ Z�3�_oSm���|�9h�-��I&C+x���L���P��['�3Wz�����#Z���
e3z	$.�Ͷ�!�2��M�g�g����%j�. B��͝mX��qm��I��W�ǚ���~:΢*�7�Fߛs�����s*��pt��%�1V�U6����l�W�<`�{���i#�=��:Ki�˹��� >9�i:l�G>�o�۸Z�g��Ϗ_3�1g����ݣ�@��5�d�3��9<V1���Z��h�2�D*�'5�	�D����9�X���<^?w��9Tq�-��I�m�i$^Q=n�-U�ʹ��m���c���#�Χ�ڷ�~�P�ͶX�2߼i��ܟiYx�@E��`f�\�!��>~t����3@��M��1��f3�N�fٗ�4� O��������/�ʎ�K;�������]���؀l��-��G�w�a�j���$c���o���f3��c1��f3��c1��f3��c1��f3��c1��f�lm3[�6���f3��c1�	$2���z�,���6�P4��� �m6���c1��ͶX 31��n��f�lm3��c1��f3��c1�Z���]*�L�c1��f3_+�p~���C���f3��%�ci�ݵ{�6�L�c1��f3��c4���3��c1��V�u�ݍ�I!��g��f3��c1��}1��n2A$�c1��n��n��f3��c1��f3��c1��f3��c1��f3��c1��f3A$�C1��yZ䔗�*�L�c1��f3�/�#��l��/��c1��f3��c��yG��yG�����}�9�yC1��f3A$�C1��f3��c1��f3��c1��q��1��f3ͯ�ů�13wlv��%B@��iK�� W�H�f3��c1��f3��m�L�c1��f3��c?��c7�~3����f3��c1��f3��c1��f3��c1��f3��c1����c1��f3��c1��f3��c1��f3��c1��f3��c1��f3��c1��f�lm�lm3��c1���[�%㱘����X�f3d0�f<�t�Ͷ �H���)��f?I�$�3�ܶ��f�T���ն��;]m�d�#䥸BZ��i�&���n����_B[I/f�P�f>��C� (��ޞ�؋ݵ��1��I$�1�����n�Q�a������6��y����0�t߅�i�w���*���7c�^Ga����`g�4���Яwk޾�$~�#Y�HE$� GwL^�IƆj�W�v3�4�0ɤ��f3L0�u���_�b��-2M ��X�.���y��[��c6��	�]S1Ͳ�T�/{dH�m3��g#n�s*3=����f|T��zڸ}��&��c��=��͹��uЩq$�Kޤ]6�|��{�4;W�����I��gN��/Gss�ml�m�M_H]3��c1��gwc1��f3��c1�ݱ�ݱ��f3��c1��f3���f3�ަMM�퍦_+U6�	'��~2)��K�
�h�b��v}O�� �o,3�]������~�6���p�sV��H��N�V�Zݚ%j�r�V�BtoRO21Ј�u���\�M̶\3���o �s��'��=���վ��/��[����� {��Iώ�:�I/�㺭�}'�ˤw�+�:��Ԓ�4p��Eށ��,)~��u�$<��Oo����6�/��)ٟ�Df�虑����I}�	��tLd���;�֓M�Kp(=[���'����w.�-�팳�P;��%�$�z�M�
�)уn�λ�����
�=se3��ڙ���`t{Ζ���_^􀯒k�mF���ޗ��FbW�K[�c1��f9�\J| �_[$/|"�l �q�dV���g���xz��:Uxz��K�'���KBjV�S����cմ,�L��-�C�JIi��]���s��trE�K�+�|��IΛ��J�޷�5�w5_�
�%".�b�N8�����Q�[b��? R_sm���Rc_��R����ɩ�"c=�$l8Y������y=x�<|zP���� ��p����[�&����-+�r�RS1$� �^���<��?n�g�b_���o�]ʗsw��������9p������o_hۮ���ʏX�w��ȍ�vZb�s�������n��d���`>GsH�"�Y�륗�e}ǚ��h���{��l���ɒ�qF�Þ�m�Ȳ��ऊ�?�~�_�˘��]�~���n>~�3�����uR~Zܾ��T�-��������}��H���w���xʦ
��)4���>７�kZ -���D�(v �oȥR�]��m���� ��e)
�	�B�y�f^ ����_}Lw��Rq?$��u 2�s�7��۰~4�R��/r_��9����P�Wb"d[���Ov�g��4��>�e�>�m�8�c�V�����HI��s0�k�/�݀�[+�(dD~;�5�i �m֨m��9]��̺P���/o;���p	f�Ƣ��"��ë%��:��S0H�!��ۄ�BOi����2�<{�V����*[юX��7i3��G R�S��]���K�=��{�ۖ���$�-���ZI ��^]�I�c1���'�R��a|cj��d��UM�KI���� 6��}1��bw��g� �C�[�?l�u�Jw�(��� �#1���M�V���$L�{��8�}���r�}p��k;����&jA
�ẍͩ��1J��>�ocR���I]ٹ�[fk�w�n���}�{�v���G�Ӛ��W�)�+��>J�ͼۮ�T��ķ����8t�{�>��_.;7u6���SI�����6g�	~b��Z�[��3%�����C��hA�5�_��I��ѷ_{�BN.����)���sA��7��1��J���@��j$�X�z�qf��I�8�W�Ui8}í7Ӧ������O���z���l�Gq������]��lL_wb~���N�O����A��>�s�;ϹMt�C�h$��� �z�b$c���;�U#�|}�0;��&�O�fL�	!�'��}�����t ��b�B���q �:�8�"~�M���" �T��Q��l>;�ʪ�V�w�  W>�VQ u��K�7�/�>|�o�`SW���1��_�z)d�g�����wV��_I��Թ��#
�i��㱛%��ԯ&��N�2�g:��}{����w_��K��ʺw��OA'I���m����\n� �o }�����I{��IQ��t�c֫s����[�2vRw��t����/I��y4���cζ����{u��ۏ˜u���kD���L �{$�#��OcQ?r�y�n�;�]�6���$Y��7O��I��4[�(��-1�շ�G}o0W��[�+7+gd�$��U�l�����d��ҷ�Y�o�������&�K">�y���:�{��j�_6ٵ�����4L�Ѧ��Ì�=#Q٢*[=��Cҽz�FX�^�̽��}����|�/8U8��}�rI�DK��}'��3b>G~"�O��9�^Q�ZI%��o���[%G��H��'�f�j�3`�۞��n�։o�pq��7 ���ww}ǫk�T��	��=3ɜ���7HTSY���?�$���A��z]��W�4 ����f����]��캽\���b��w�ˀ0rI��z]�T�/&,�{��b���I���z��o g7��ޕ����`/*���iŦ7P�ւw�y#s�H���b�7�6φTr�K�۵S �U��H�+�fÊ��\�� -��h��
!�y¤�$Z4��?��y?t}��������<��IQe�	+պ��m!B�ie�����<y�!4�z�/R.���C��٩K�~�~��U̧�ͩ$��K�x������+gw9��d�k�� bIm+Wޜ���h�3�}�}#��u~4qT���`T I�v3i��y����>o_���ķ� ^~�[ܒ7yl����� W�P�XX8]2�&/2L�%�#��mI#��ԓ B������A4�O�'�)B�1��c���[���g��gY�c��T�Ͷ]3L&/�m�f3��c4�b�I!�m���ƕ�c1��f3��c1��/[����<�I{��t���3�'\чg{�m���gc~ֈ�z{���� /-g��[�GK��I2���o���i�Ƨ��2x�f3��jL=�#��m�d7I-�	Cn�+M<�{�N�0�p�f3�p�/��=��z� ����}�&��J��	�H�v��T�̻n�M|����:��$�+�����i!y��B'SL��]� nx�!��p;m4����"X�W�H�`�B��F�s��I�c1��a��	�a݂����⩴�f3� 	���)��n���ْx�?cD����y�~4E7l�c�c��c	$��~ R��z�IL�f3��c1�̒I �C1����H�9ݳ��$�^�����{a�G���s����>҃���^�ڲ̆��:w^,�X����0�]��I&�*Lžy�Ϸ�&���Q�m0 )��e�,I�,�{���Jֱ����s�	��~�kD ^���n6�F�v�o�L���<�1+���@e��R��Γ���"�\�X�~$�1��~$��-��žm���K���L�C���$�m0��m�-���p�!����n���,�J(m3�2d7�:U6��$���f����Dl)���f2�U6���c1�͹��}�s�tY��f���i���gc1^I)��㱘�p�9��n�>wT�<.����$�&��ĝ8�d +����͑�	'+O��k���%�'/"�HB�'�@,��{B�o�P (�X�����d��c1��mU.�d���6�r�.��Ǖ��r�Tf3��c1��;���.��Hv8{σ�:d8l�I7}"GCRJ��ǚ�z}�H�{n&|}�J�cin)��^Z���3,.�Zy&�sĬv��� /�/�w� J�ĽD��Iq@��'ޡ�xχ�e06�{�|�w����V�~�7W$������/��ww�C���������z'��ޏ���y��������>�@�:�J�<�E�(���k�><Ţ}|���N��5�����py�$]�^I,I(LMN���gC	��0y`��W~�W���O�?�������|��� ty|�����z��$(P
�Y7���ݾ�rQWV?O��H �=~�+�w���HA�X�B��%�w$��E/|ϸ�C�[���W
K�f�%8gI.X:�`Bc�3W�{����5���|Pe�qao���L���cS�p ����gV���^;�{�Y!��X���(*�ֻ�.� ����ʈV^6+�T�!����T�f8<�t�y����`k��x�~˥a������l��]� <���i{���(���4���*Y$�_n�{�LSğD�̧1��kͼ�IP	�{���v\?��x���X�i|q讌�bge�mD�Kk�nu�D�8�[g{X��[,~-�۵���/�^���T{��\�����m�[-�1 I��T�m0:8��{�l�a��c����-��
�S�3�^�N ����$K��������߰ڏ�d�7ܭ��)��U�$��%���zIjq����Ȭ�e�S>�D���f��XI?�{y� �?Q�ș�4��z�;1��>�����5��d�K��� �n�<�ѻ�t2�O�&�A��t���+ ���kqjr@Y}�r���HҀoI;z�)P�'���tnc7�K��`� ���I�n��ǋ�k/�3��3�w���[�i&��'aݰ>��Ģ_���~~W��[�=�D��|��	�IQ���h8�=��wB��TwT�QsT*zj��?��=�ܖ���2T�)Ho3��̶�]��{�1#���ٷ�#�=Q-�=���m���K�ݻЧ�?���\hL�<�T�]�E	Vc���F���j�U�o���z���n<�GA$4���z�$V�2yy@��#(~0&�	E�%�xY$�	����\���c1��$�:^�*H}>��%�%I%�x�i'�$�u6��wU|شpF$n+Ȑ�����3<��^��X
XOF/
�7w��7x7_��N+��C�4�N"Q�f<B�;�^�E�_{�'&�8���.9~����$:۶1xX����zJ�fݭ����Xߵ+�W<�X� d�a%�t�'=�sO��������hڟ���o�!�bb?��/�A�i�d���{�	��f�ݤK|m[%U�=m���i$����f�w��f3�2d"et*�/�$��dΕ<N�^'�l�f3�U����Ǿ�O(L��N��ǋ��B�]h�� sѝ�����8�l�̒�fz����7�üWf�{��udɘHy}�]���׋�S7���L�^�{�w{�����{�g��
��U.��B�|�(��Q?(�TH�ȖR|6����D�mD�EI()
�(ƒ$!Z��x��P4 ���ԊүT TM��b�S���) ��� >��x��J�WB����R&�J��|��&)� ��:	�R� �H#�E�#����˵
6�M lQ�:l~O��$#� � ��$ F	� E�bĐ	"A���H�#��HR�Q)F	$P�F$B6*R;^�1�"�$��a"ă1F,`�BX��`
`�F!��, ���zA�$�bH��D!!�I	!Z� H+��P � ��B? � t*/��=��a#8��uM�+���
4��b�� ��A"��D@�Dx����� 	`�U~[E1U=TA�D��"�j�D�(@��-A DSaH�(b �*n��`W��E>D9rrI��o��Vd��j�2�ƆUv�w�C!i�e�4���H�&j�5URk�DiT2�*��.�f!��tةCm��*��5q#lp�1�GF"�mj9R��B�pd�W!��1�X�\M6�QЩ�ʶ�mB��Y���#e�gBjR��b-tܳJ2��sZ55�M�quA,\;K��hJh��LXX�ف5^Ze�Ep�%�-�As���o]v�3b�1��@����S@�� -�b`�����CZ�r�2��ղ�,�+�6���5�]n��،����c9[\���Ga�L�-�e@��cCj�]ٶ��t���n1�gKq�ιr.�x��.ƫ�+�&(M5��r�e�Ƶ�]����i.�DPpɍi�I�Ү]�2ʼͫ�WJ!�l8��N(| � �D|��(sKA����{=��a�n��X9�m�14j���;:�Wn2�
)b��pJěP�Rjp�7.��ģ���-���s;f��Ν9�ӽ'c��y��b����YT�<��������� sm%�Ϲ}�IZY0�T����[>�V-R^ ��d���l�O�\�$�
���$�H��O���l�a6���uh�s%���$Mr��I2m���$�"Kl��!$�]0��lQ�Pd�x�m,�A$��-�撽��$���O�Iqe�f�8Cqa���$��������䨨�GEڗ�qA�7M��	�clHx��nܩ$���D���d�$�A��x���I��]MjE�p�-[\�>jI{Qlm%�>��J��$/o���v��j9�&��n�P�/�����j����J�^�eg�yR��{ٿH�+�$�ݤ-
L_���x�ZN��H�jQ��;�z��q%�A�:��`Ū��R�B�2�I��I�Ka��>�z����D�L�N��A6��4}�m�z�2K�,�gĨ.r,h)utmɋ��C���-����g߽���Δ�H��OW�I�vUIڴA6)Mq-YB�dXq���oU�}��{̓*Gt,�O���$�@Ii�ϰIC�Y�wh�0�U�N���m�O���2L��$��S�D�4�ŉ��$��n-���K�߳�I{������@�K�0�w�����h��9�PP��>���	y��������L�L�����N���m�O���2r���F6H�M�lD�_z̿}�)�wOd�FˌR��2�hF�f��'A&eP@Q�M\�JTH�6OW�I8��-#�6	�׽�����4�k+�P�u���]<��L���Y$�,=�IҀ��$�d�{�+�n���"D�66n�$��u�撶�$����4���nM��u��:o�*�>e����'��A��e��}�$��:��I:�N�0kH�Q
M�5�mV��߳i�k�!>�~��	::z�>1BYM-�ijacu��Uf�e�gk��
��덲!���-�mX����f�'�V�SB���-�5�"��:E��m�nA3-�b�
�Z7���%�kA	�]����2�u�̄I��gKX�2�B�F�J�M:i6�wN�5�$-4��ug|�h���o�n�^�� ���ي]6/�v�B1m*4��P����*a�Z��H9���|�g�S���OX���[\mc4l��bh��bz������ I�����\��
B쓘5BB{�5}�b}��D��@�$���}�I���H�3g��$���M4md�,���I�u'��2�]аI8�b��$�"Kl�j�L{֝��)�x�t�!vI$�L��$�.��I9�������8��|>���M���������������#\����K��-�K��PX�뵪X˴7���k	$�]l��&V˺	�mFI��>g��2�lU6���*�6���!�kk�\��"���(�3j�2��I�3j�hf�,�, �v���j�k\:�n�vWWI�>t� ��J�vf�*�Z+��G/�I�D��'�'��$�!H]�I>�Oy��E)�n�n�&Y�d�s��w�"9Q��l��;��I�q�$��!$�]1��_��O��2�]аI8�b��$j�%�I����h	F�Q4��nM�Q%�$�_Uo�4��L ����O�Iv���׊[���>�I��=׾b��Y��R���ޙt������spvd��6)u	��'��;R;� �͊�I�PB����d�C��T�n�6j!35�O���+�~���9�P�	���ﾬ�	���X'D��摤����[��ʼ�ouU\��sG�e1e�J! �EbD������j�qR�ѽn�T�0�j]J���}�Nj
|K 6��V턃,;$���y�F���$��z��������魊ғm��;�����C�ە@/�刹Ć���7^%��ﾽ��KxV �
��gg��R4ɨlZ͖*Gk��ާ�Kf�}k�����^����d��X�����u� ���u��� ��:�>Öu�BH��Ė}�,�������q���}�9@!\BdضJ�h�`��`	�]X?W����yb���{����ײ-y75�q���4>��T��,A��Ӌhޥ�6l�<�1��@������I�f���V왴��[��6�'���}��/up�� _���6`k��َʊf��٬�6���b���_�}���3�=��uW�}�E����9�4ݒآb�y����B�ڠ�� ���i�Gf��[�o�5��Ԡ�̀z���/r�zِ2��V�&���B���W�W�v>�6 � a��wy��&�4Yu�K�(�&vJ0Ɍ幘��l	�bl[e�� E���1�8�m��3�,M�lD*��h�%l1���n)���4iu�m�����.�{h�l�G\[�-à��c<�Y�Z�ec �&M�f��ir�̬�ͨX+�=�k#�s��˕wZ�5���@9x�h)�b5�-ǄG(�p�I[v�5��\e�`��/�^��[2�9����#^���siu֚^�܈���4X<c�fF�f@>��Y��ܹf�ם }�U��תĔ���¬���f@9x�h�٧��eX�ᬃjlպŐq�,A��V �u� ��:�=PZ�&�(�a7fjm�~Q��צ���O{W'h�{��P
�}��$2��%&�Z,4��SV�N���ݦ:͍bT��fFi�R_Ư�E�!�Ht�4+$� 3F��@Ð�"V�-�ݧv~����Vv��aV�M�����Bmu�r1Z��j8�՗5�m��u�C���\&�ci�6[��96�m�
�bE_��s�X�nЗk�A0f���`�π�,A�r���@<�u�~��$�5�9��f�+`M�]_��$i��h�δ���eŝq,և7�<i� yz�{�̀{����˖iJ[���#M���}_Qբu�2*�h	�+��m�r�%���0�S� }��vt��X�1.\lMHU�eؚRha��ɂ�Z�U�O��}�������́���6��5�u���.�=�v�n��5�.0���R��=�Բغ�@�U:���Z���n��F�΁���}䓒�r���h}y����P=m��	�MN,[1�١}�d�] ��C펥�+64U"7e3h'I'`E[&���P��`��i����(�y��co���j�h�ıƥ%5.̹E(��K�[�5�35��:��^� {� {l��A���gm8�T����~�LǃoZ)�,A�� ��u��c Zv��Q�(F����[ :��C�ΐg���yx�?�~Ư��=�f��EŹ���_� ��N��%!��)�u(e�aa$H0�%���f!D!�-u�A(n�F&�,e�H#Xh�U�(�� Haa�*ʁ/f���6Xf�ѯ����SpeXʽ!+Ƃ�R�B�B���!F���*�e�Y��t�X\oZ�H�/T�!*�@�,��$$
(!
�M�	�%��)�Q
�B$F�hIn�$H�Q�R3h]X�(-#E�
���K�-�6�ƒ�4���L���j��c�Quv� E�%5HH��`@�"���$bȱ��I�j���H�H��!9�KH2�ysmQ���R�˫Z��Eb�X�78��M������x`�l�,��Pl3�A�6[�jj��n��ƪ��a���+Zֵ���[ut�\�V�Zƪ��V۫Z֨�j����n6�Z���A00�&1��c�1��l��6�mK�KQ�bԢ��
j�a�b9ÙS5�i1+���}��j�
Z�� -Πh���I�ak]������a�.��8K�r�H�pL ��-�η)�li��Z�a��LC<���R3�u�j�0�2SL�L]q��*��M3m������pU��Wl��UK���bCn]�ք��z�Nf�A��e�%*K
�tU�)�-�@A�e���R�]c[���\j���,,h���sA������+����k�k�cu[��r��MƇ4�-�t4n�Nbu���Ƒ�	��j������ܥ�������z�z:�cC�Κ��¡�ݬ2֋�c]A�6�3�h,��؛m[�KU� F*c�\��d5Xj�(VM7)�422���qd2�`YPE�Y�ܑ����9�����l��U���[e.�n&
cA�6eqB�&ѵ٘)p��+Ze�4FQY���G��`@��ݥͥ�s0ǮɪP����M�Cp#�T�h��1�L�ĸ#)p���-�.T ҌQu�,k4�����Uj�ܓ��s��0_�]"A�
�h���^ �E ��q�"��(h"������w��I����3)kM�o
a_u��|�� :��C�ΐ/��M�$ȱ�(M�o@���y��;Xk5Fƙ��s����lTV�aŖ�g��}�@>���W��|{��ZX���fj��F�Fb�6�f�� �t���6+ {��6[�����=ܬ�:��fղ*�*�����j�y{��>�t���Q�=#z�lѤ���ʠw<�����T�=�sjԠۛ�M��@>W��^��ΐ}���1f��?�����iK�+u���)s�[͹�E�m&P�A��ft��V�R]*�`�*�]A��,��T��)�٠�wV�+��d�^R%�7+Tm�D�\-�������ֺY�6b�KS-2:\�6W<��k��<���cnΜ瓓�yO���������a��qFu%��}~:��x�!-��a��@^\��K�E�V��˷������9@>�<a0�#���҆�=|,�c��nҐ2h�I����C`	�-� a�gUyNVlB�ӧA��ݠ��� eb���W���ΐ{�X��S��%�Q7����Z��^-�]�@/��@�����58�m����m���H�nu�^�`{-ڄޘ޻��k���_����Np�yZQ]�.]��l��j)�ėM�H�B�އ��=5Բ-��ߨ6�zt�S�\�h2�n�\b]@F��׶A����6-P�*fnu�,Mv��lH[ZY�`�Z+���jQ�.�8"��ү����${��I`�����]����sf�W�u���|���>�@=y�x�q,׃�7��שn�^د�UQ#:> ͏��3#0�A! �7�i͘�5�yx�4>�����g[ üz���R]�I�Sv}_ӽV ��]րÃe��|rK��6��k���kOul��݀�9����x��V���2�@MXʷj�r�w�������/����:�=���M�6D�SLE�h�XїMZT�W�Eݝ�k�;Ǭ��Z%�6k���@��S����6u*���+:����g^s�4A����=5$�l���N}����@��~����H"7e-'E+�7�w�@Lخ�w�N��@ȸu�^��)4M��+V\��5'�P�_�=�W'����X�.��9��XB�h4.Ҫj�KAH�� �?f��(nn}���\��Es���46��-0�����w�@H����*���jY��_8����El5����}T�A��Eì��\ ���uy��D�Bp�9� Z�[b�Xٮ����`gs�`j�������[d�];-Ѡn��l�꺰���uY�$"B0�*�ND����	 )h�4��
`�D�A���!����}���������~}�Lj���������O�K�v{��O߽�F����٩? �~U�ˡ߭�����F�����6B ��߾m��E-��-vT�#Ȕe��J���즹��	?ܒޕ��@~���]X�%Ձ!�L�,ۻ�|�QP��j�ۙ�e�߿�>N���J�~�_�����Y��W� B)����F�?{��fd˚̼�]L�y.�I7�����/��H
�'}���N���թ&�g{��@?��7������.��35f�̹TV������I7��wU�_ȰF�߽��T����ӡ���}i�7z�9{������'$ӻ߅�6w� {���4쀬����wVꢤ[f�.��\5b��2�s�T�m��˄�����Ԇ�����L\�])�-��C=�DذI[5��&�s���Ev][V9�s�..	�ͨ�����
](3j��mY��A����W�r>����F��#��M�m�	�-��KV�_V��Jkl��.��T����Z��,�AQ荒d� ��u`j�Y�B��N�ua��t~%�<�͕��hJ��I���yA���ŢY7\_x��:����ː�/��]��o����������?.�l��w�@{#�/��pq��t-]�*�)��������W�_��T��X~\?Y�j���eYT�VUQ�;�`�Wu�<tIhw��q�>��~����WE���=�� �Ͳ�f�j��A�fc�9�Wh��i[��T�����guhր�]K"�	��M4͢ϩ���������CF�s.�X��Dךe�3��X��5b^#vo	fGb#2r۝��W-%4�b�iWWcWB�hL��\�e���Ny%̠w\te"�E����H���mݔ�g��Yf�,������Ъu�q�)��w`�Z�N�j�o�����!��~6 ����rO��vk��"]��I���2jV������k$���~�Iߧ3�S�/�`7�~�l?s�,2Ja�Ң�'v�e�U���� /����ԓ��{��M�wU<��-�����'W��5�ə5/ZԬ��� ��H��@X�a�=��zk\�`pb+]WM�����U�for�E]ր��Բ6V��Sv�ç�:Q���Z˝����*�[D�:> ܎ {�z����
�@i������~M$�-�7n�V^Zԛ��L ��B�}��`	��X�lW�W�UY�k�Mb��.�&�'�;��R}��kS�D���s�?���?���v!A�f¦��TK+5'�C��=?~���{ک7��kRyD?�o�5'�z���.�.����ˎ��y~���:c۶�H�C	AEL��Ф�t����m�������Ov{ک>��>䣽�f❷;�f��+.Gj�r%�IG�C��7z��B}$��g�&�/��I7\���X�'=�?j��ŴJeӰ[4�°�9B��_R~P?�  ���߳�jI����z�}��~R(��������VJ�����wf���$��߫RN��٩h@P��@AF!.��g�'{/߫Rn}ۅ_jfj�k*�*�RyD?* �[罳��N��~�I���&��~@`���!�{��������oU㺖�z���@�����:q�@�[AEeltlS�[eS3*�aD*����� `� �Qz~��?I;��?j����Hw���̙��/an��nZ����H�Ĭ�~"$��@����K+> l
���<sb��]K fGRȭ�Q|���V���[,�}������9��A`$����ߵrw���jI�Ngf�'�,bK�t�����eZ�GZɅ]�R~�hԓ��vj~�"���%�~�h3��`z�C%0�6
r�Mu��?$E"A�����ک9�g�jI��;5&63�J�)!D`�P�2�bS��"$X�%
�R�˚���W���]f�(������+����&s�MG#B]t�u3+��Un�5sHM�B���fb��LK���j���V�P֑�ݝ*J��x��6���kC��D�L)wX��!��:W��ݜ�h��v�RXl��e��'�p�r�
�I�~�hO܅~4�t�Zv¶�h }=���	��k
�.��"��.��с6Q�Y���Ct��$H2 1�w���~�?~���w���I��p|�Tץ;	m�aݵ��-�eL.]]\�s��@�$B��n�I604�ߕ�2-�������"1X�`@�P`쓟��P�4q���n��n�L����_����b*�� ��X��{��թ'����RO������A"�)"�$DH�]_���%7�7h�cor���� q�l��z݀{���������f�Mi�?!���
�#����MI?~��F�����W?~Q�H���K��~�Z���O~*��+VVaWz.����_'}���Pj
�}u6���������)3�r���e�K�S3%�]����E�@c�������%A���_픛�Q*%D�f�RnD�����Ѹ����p��(�D D!O�H��A^=����8o�����.�i1�����4aY5VP��2#$>�D(�taW�aXJ�V锾�C�E滭n��HU��c�IN�������f]�Ma!�f R^f�I�°2�z�0��RB�F��1�J�£k(�8PY0�� �,H����E�,�#�H�Q��,� ���+�C%�`J�R���h�)�Ca�тG0��S	d)��Q��i)&��6�ʽh0���M[�)�	���Q�WЪ.�U�d"�! ����B1�i$��r�T�`]�0m(i E�,X�DcXE�)$"	�HE`�	E.$H0",� ��E��
Vŀ�|x�j	��A"F0�" ��0!�E"1b0`B }�0� 1`I"�"@�����nUډA�9���%�4͚�c6�p�&h��@��P�)�l��, *�k�v3�:�TZF�hl��AUڳ`]�TUۦ٣�!�Lv�4t1�i5,!J����S�˵��(�j\K��Z�0��WA���դc�7.�it,cG��˶ �b[1[z�X$����c,Ք��5�f;M`�Lmf�%�����E1LJ�!s+��W���ae�A-Hm�1�.��a555�����)J�4QXk�.��5�l�\�r��`��u31骘�ȑ��"�@�+vannph<�t�b�R,5 ��+��@�6t8��dfH �l����e�Q��jK�Vit
�QF�!��s�Z����݈.B�^a�dˬ�6)��i>V"6�S@�&��+h	��M��8���w&Y.�����fR�Ԧ�����X9z�.�ڬ� ��8e�����3��m����F����u����gQ���˲�-��
X�iYY�
�[	_��
����y��������?�n%���wFz�\J�P>�u�h?>�q*%D��~͐7�TyG�?I���F�U�^��^��3A�:�Q*'������	��"n@������4��Q*@��_���ȕ�w�~�Xn%Ĩ���L���	�7W��̬��4��PjD�f��p2%A�������~"%ĸ���_��T�Q9��?hw�T}��_���VV������^����O�@������q*@������M�ȕ�}�;�&��
���\Oǽ�(7��=�?���6����}Z{O���|�kЃP;����pnD�o$���0��X��ծ�%��:�,�.��(˽ �����ߍ'��TN��_����*%D��W�Pn&D����a]�O���{�*�ٗv�l�Iy�P��iU�֯U2�q*%D��s�3�7�TJ����<@�K�Q*'{�l�n%A���k�������S�S){�	/�ǚWy��9�J%D��߶PnM�����)l0	A	�Je!bbC�>[>>c	D�IA ����n#VL� �M�0��Ma `�i"S�DH�cŁE�BD��qU�jD��5�C���s/���pnD���o�(7�A��<W�߲虓F�^�5��UaZM��J�P+��~�n@�����҃q*(��}�h�D��Pj��M����e���J��^�Ve̻4��Q*?�.'3��?@�K�Q*'}����dJ�Q<s�٤�J�P�d�������ȕ��~�xandѸ��K�^���n&�TJ��v���q*@�l�2�x!o�~F�i��i����Ư2U�3!zy�����D�5��z�prD���o^��Pj�{֫nk�M��Q++���9\.�2^U��� �Cf��7U���T���џ��p*%D�=��q*@��_�Y��A�b�Aa��Pja��I�9��_���e������¯��FzO��gB��?�}�����$T��cq.@��{��p2%D�����4��P*%D�f�Pn&A�}^�ʗ���73Utoz��U�7"T��{�M&�TJ�Q>�_�v�Q�6�pl� &�B# $T"!$"�
,
,EH"$RQb)
�q=�������~��oR�T�k��˲�2�n&�!+{�U4��Q*(�G�Q�!B*�D���_���ȕ�{���O�ĸ��}|�I���D �?�  E��Yq=�~��@����e�2���fd�jMT��	"'ܕ��j) �~��)'�1�+��04�Y��QЉFQww�*U�/B� ���׿h@ȕ�w��~��7�TO���]��T��(��%�.^����U*��Q�oĆ�GFnq���wQ*@�=�M���}�߷A���TO���Ԋ����w���M����^���3&��޷u�3f����TJ�Q;̾��p@�SQ.%D��߷�q*%D���W�٤�J�Q*%}ʾ��qT2%G���
�O�����I����^����wդ�J�Q*%}����d��{��oR��
�Q;���t�Pj{�O��������f�焉�OȐ.��o'����r��e��T�Q=̿z�p2%@�kw��Z��iaUbS4�[�����L壆eK�J��7Q�aF��vmLAcq�kay���J5CM�2����YEn�\���C�bjԩH\��!m����[���+}���v�50:-m�j\ѹ��Eq5�ļ&��*�����@�~j����I�5��{-��mS���|�����W�|�8����*��M�ȕ��(�􁿌v�n���.�%lֱ���Y�d��?�����p*%D�2���J�Q*%}ڿ��L�Q�o���6��E�w�� �n�ۖ`^�T�҉�>^��^���~�I���TN��7"TJ��N�'� 7�TJ���}zMĨ5'�����#����������%�{��� n �@���ڿ{V�PjD��^��p2%A��u���-������e^Uz73w��W++A���TJ��~=I���s�=���Q*'/��e�T�Q9ܿz�7�Tgy*w�e�Zw.kE�����%��"TN_;��n@����~��d�Q=��z�7�T*/��f�q*%G���T/+F�o{���u�&^f�q*%D���u�ԛ�7�z]�'ȳ ��eQt�LA�Sm3Q�d�ev�'8s�=�'�d�Q+����n%D�5��z�q.%G�zO�a�q+{�S�NK�е�*Ԅ[�[v3�Mi{�2�l���Z��p�k�aцr^h�M�.αe�Ʒf+��F6�9��r�t&p�D�U��w����jM3B�nфncY|���NJ�Q9���I���TN�{Y=A���TN_%��� A�
�Q?_o���xrRr��}��R��K����ܻ��TJ�P9}��z��"#�.%D�~�~Ն�T�Q=�h����Pj9�}���Q�o�~kʬ�����3f���T�Q=��'�7�T���k�M���4��L�����a���TO�O���I�����;�aM��ɷLw3ŗ�xr'%?Ӑ@d��;���7�TJ�����H�Q*%D���y��q*��\K�}�4��Q*?�~���j�+F�kz�n�/E��7�T��0���pr9)�����қb�h��#�oiq�#M1�K-�-���~?���v%A���������r�/��xN$����ԟ�j����;�3y�f���K5�]H���rNr�w����L�}��
����������r�=�&��
�Q=|�{-@�%����~ޤM������&d�;���ݻ���n�TJ�_s��Pn
@�8&2��������q*%D�0���q2%D���|{4������Rd��K�;�Ò���K�c�xrc��������Pn&D��������Q�D��Q���?�O��Mĸ��v�/����
�;,�{+&V�ĭj��6�h7��
��w�4;�Q*@���y��p*%D�����7��$���~��Ĩ�~����*�&�p.�oreV�pu�TJ���ڰ�J')%"���c-XF�4��P]�"M�X�-�L��-!����Dd}�{'�O�.%A������d
�Q;u�{07�T9�Y�Ud�����%v�u�Ҵ����T}'�ѳ�!z~?k��I���*@��&�TJ�Q;��6G�@�O�\J�Q;~�^~���ʟ�_�\�Ѹ������u����Q*'���i7��)a��j�a����*%D�_���Ĩ��w�צ�p*%G��z���ff��޲^���UVh7"TJ��+����j%D�����҃q*;S  !��U�RA7�z�?~��D�5���Pn@��{����^F�^ky���xh7����6,��D��W����Ĩ5�{�����
�Q>｛ n%A��2�w�/ߩ7"Ta����T���|�>��`��|��d/B�}�ۿœÒ������xG*��6%V�3]KV\�1��/2��b�y�~�I���Y�ߴ�����{����n%D���˯Yv❞�w��rY����6a�3
�������g��,�:�[6Uރ�7�TO������ȕ�w���&�TJ�Q9}��z�\J�Q+���n�oB�����&
�z|����_	��n%A��þ��+�"�d�_ߪ����*%D��ׯ�A���TN_'}���X"j%���O�fI/&��͹����zM��
�Q?{�����q*@������7"T���ﴛ��*%D�;~�A�������aT׳Ò��gͻٲ���9)8�K�}����q.%D�����4��Q*%D�;�=q.%@�� ����9Ϲ{��{s��+(���!BQ�,YWFݪ�8���Sn4UgJ��
�ɒe�S �����1�W�]+1W��A��\٭��mD
5--�]2),%��m-ɳ+*l8���2?��JG�!�K�5J9��nvy��H (���&��rr}99%��D�������q2%G��_�.��	�q37+{�U�M&�TJ�Q9|��Pn&���n�n��檵9�n����4��S0����?>���:�Q*'��׵V�PjD��{��ȕ����+2�p5{���5T��%m.�e��"zw��>:l>���~���Ĩ5�r�+���D�5��ߴ��7�TO��f��Pj���ʫʢ�F�^f���kW3I���
�Ǵ;��D���{��_���J�Q;}��ԛ��jD��_�A���V)��L��l�����1��dϼ/��Ǻ|�ЉQ=�����Q*%D��_}I��TOs���n@���9W�Pn&D���VH^V��������e�W��MD������> n%D����k���D����^_�7"TP���u���q*<��x�+�[�R�[�+	ZMĨ5�}�=��dJ�SO����f9��SWER[�r�j�6�￾O��?�
�Q;|�{,7��
����;��*>�.k$˪�;�Y��=H0X�r���%$�~�����&��K��V˱��s�K63�ah*�e�T�W�4h���W�Ib�YK��),ւ�M]ٔlDvh�V�]N&&�c���jb�<���xs�,��jD������a���TJ�=y蛁q*@����&��
�Q;��U��_]��M��ׇ�i�j�kS�n�T��wG������Ҧ�dJ������7�TJ���_���dJ�Q=�k'�a���D���?��M�7g�&��㥽���%9*'���~��L�Q*'y�g��q*%D�����4��PjD�r���dJ�;���-�̭;���{�޲����P*D�{��~�Ĩ5�W�����p2%A��u���p*�������Ĩ5	���P��s2f���蹻��ԭ&�n%A��}�4��p*rRw�RX;`�g���˷��.��Vj1r#u�=����t���TO����M�ȕ�{�צ�p��^�����]������`@�D��TY��L�ʺ�T̟�� ��5��ʪ��}�TJ�]�_����*%D���� n%D����4��Q*%D�wמ��ȕ��e�z7�[���[˙W��K�Q*'����p�bm+IM=h ��%YAT
.ƛP§�9"��TL�}���Pj�~��L���Q*'/��e��~D������p�~�مd���Y��Qw6ևp7������Pn@���d�{,7�����ڿߩ7"T��{��&��
���̗�a�q+{�aW�4K�nD���`$,@���~������j%@�}���q.%A�_;��n%D������a�����|T��2�M���oZ�f��M&�\J�Q9~�{I�7�T��+��-�m>L���u��"$@�
7l��h���;�K$����BE{�K����5�wߵ���q*%D��s%��a����v��ݽ>^�z��j��*;V.���T�=;吽н?ߟ�ߡ&��
�Q=���@�K�Q*%w��f��"�R"��\J�Q=�k'�'�ѽ�߿���h���d��|��U�7 TJ��r���?1.����{����Ĩ5��՟�n�������q*B}���Y��4n&kz%l˗y��
�Pj��;�&��
�Q+ܿ{V�Q���0bȢp %q`P.��$���D��� ������%B@4�	���7�&[� �*����FYIBD�A!E)�QMB$A�"b�U��"��P��4@`@��1��fM%$BX�$!rI�A��VK!E��+aE������ @����D �AB0��h?�t1�����~P�?�L;	��1��@J���5	GW7L��U���sb�\Kt�:eQ1T�u����u���.��SZ
�q��$x&��lp��1�{7l�c*��u���P�1Y��[�1�cU�f �4rc��1�`�͢�dm���˳e!]f��cU��ia��ÃGd/g+sIK
JUZ���+[�
����\b��6�!���\�Z�j1�S1��d�h:�\,���m�P�i�sb��+�M���Ӎ���[l%	cfG����	�L�5���h���9�Qƥɶ�*Ԕ�L�q�E�K��M�]Nmh9����h�P�PDla�Z@���s	�*˶�m�P��픋�m��p�%D˔�llc�:���îqJn"�B�!5�\sR�6����F�f�˲l�4֍K�h��[1�2:�UuƬc�:m�KZ�e�j֥t��m�����X�e�^ e;1,�Zl�l�fF��֛*��Sc]�h�J��6f��h�lk��.�V�R�U��M\-���Y�)[M�Y�bˍ��-.�Ś�V<��am-75E���-0̃�,k�M6(�e�;hd�%l���i��Z6-3D�ڨڜh�&C;�ZV�bh�(\���M�D�E������3i� ��14�5
�-����q��Gce]2�\��3�ueq����4�W���M(��аJT�i � �b"� �E8�TT�~�hA��� ��7��5���p*%A���~�n���ޯU��%���[�嗼�U��7���Aq=�o'�ĸ��r�/ߨ7"TJ��sޭ&�TJ��������jj�q.%G���u��]��Ѹ���Y6k4U�7q*%D����&�TJ�P�h��R��2DK���� %��ʪ²̹D�+O=��h{�T�랫��7 TJ�\��ڰ�J�P��_���]�O���|�b�bf��96sub���9��	�|�3vs���{���A�5�TJ�;��Xn%A���z��B E�D�5����I�9����Ւay4n%�w5�j��34�PjD�;��j�p.%A��v����Q*'y��]�TJ�Q=��=T�5����{	Y��F�V���w�y��n&D����{4��Q*%D���z�7�TJ���Y��J�Q*%w���&�TJ�;<z��s�E�y�]og<$�%'$�r�/����Q*'����q*@���}�4;�q*���p!��	�Ci��ƈ2�*��%�I�B0�:�04P���B���\0���SUE���	R�$��"�� �(�PJc"�STJ%�8:~w����֩�9�t�*\۩�n���E�kp��4�`�5U���Tl`
�1�
�1n�.ۭej�+�i��Y5������J��6jkk�YMS.1,Z������:��9ک�")P�(��&�f)2eeJ��u��+2��|�U:H��g��p*<����Y�������Z��&�q*@���u��M����d5�B|�� in�Z��3��(�Y�Q2U��NW}���Q*%{��j�q*@��s��U&�T!?���%γn��L�i(�xf唗k0d}�W��q�,��Y�
�=��Xn%D�����҃q*%D���K�7"TJ��p�����*0����(�2�n&o7�^�5�fh7��
���k=p[�Pjy��i7�TJ����4;�Q*%D��U����*<�����xaZ7{�]T�욺�n&��
��;�MĨ��s��z�7��WyW^����D���o^��Pj��x��7��T�V�*aZ�ȕ�}�/ޠ��Q*'y�f�(7��
���k������z{I�7�����˕�7�7�����̕��J�P*'nr�����,���.��j�V5���ҊS�5ux�J�U�|��>�����
�Q;�߶Pn%A����I�������̲e��M^U�4�O�E��	- 44E�#�KJ�RR"��@�M�?E�-R�d�k�0sun��<�ͳྵ��R:���l�K��8*4�3�x��,���pgqi������3CU��ũ:ԘlĶ;2�%������5XU�;q*%D�����n%D����}��dJ�Q>��S��3蚉Q*';�ۓI���￷��u\a��z/���Y�>^��D���zg�np*%D�{��Pn%A��9]��p2%A��U����/N���������:�|�>{�>~k��J�P*'��~�����WyS��n�TJ��v��A���TN�%�ԛ��*3����Us34��Mn�ݓI�9��)q9�_鸞�J�P*'o��?D��Q*'y����q*%D�{�M&�TJ���z�%d���3W���Ԫ��n%D���U������Y}�|P��j��MJ�7�k�U2���Lv.?��:t�����I�J�Q*'��g��J�Pjw�u�Xn�T|{��e�z75S={姜�a�1r]�(0ת#�����J�P*'o����D�5�a}���
�Q>�oے��>�pjD���~��Ĩ����f��&����sp��	��������A�P�� �I(	�D��F1��b"EH�B$A ��ZCH�L���p*'n{ן�n�������I�9���������'{����w�7���[�h���J�Q*%{�u����j%D��w;=����$.%���_�Pn&A������q2%N�����fr����oK�����мT�~O��2'��`�! ���A*!"w����R@����w٤�J�Q���X�0���ۼ�zk��OD䨕���A���T?��kr�R�?�^]q���̴�V�r�T�J�.�?���߯�����TO��~��D�5�e��a�7��}�z�vW�Ó����R��l���o�}i
���A>I��8��~�~��D�5�{Y��p*%D�z���"�.@���~��&�\J��~�2�+4�k{%o%�ޓpw�TO_���Pn%A����z&�\J�P=���I���TN{�ޓq?��t��޳�����a�oO�����Z����*%D�r�_�7�TJ���}zMĨ� �1,ș=�����*%D���z��\J����e^[fh�M�W����4�Pj �O�����Ĩ5������z�]�j�q*@��������Q�e��dA[�xI{�+�޳vO	�INK���e�T�P��^��w�U��ia���b���ٻ�ғ/��z���O@ȕ�W=]��prD���_}��Pj�rz�L/'����Ȱ����ZW�c`jaJŗg\�{��'�%')'�~��w��.%D���u��J�Q*'��~�+���TOw�3�7�T~=rx�^VV����n�����&�q*%D������7�TJ��wY���Q*'=���Ĩ5�Wݕ�hwȕv{Ɨ��焗yv��]��8�S�������J�P*'�þ��D�5�wG�&��
�Q9�޽(7�ԟ�o���4w>�/E�W�5��>Y5�@j���n��5�����7��
���s�I��bު��̍ �,�M4�T����L�+���j��
��XZGl4M��2�
��Mls��qJA�D57����J��IV��i�v�(ذn�Q�6����NV�lH�\��N�`E�tɈ �:���Qb����g4^N���}��C��w��e�e��q5���L���n@������OD����;�!Xaً�s�ص�i�4h1�1��#�Gz�ޠ�L�Pjo���7�TJ������J�Q�܇}RQveh�M���=�-��@+��,��VҶ�+(�A�7�TN{��U�T�Q>�wפ�J�Pj9����dJ�Q+ݝ��ĸ���us�U�h�J����+I���TOs����D�5���A�5�TJ����Xn%A����;��R\}O�ğ�4��tn7��3�<'JrS����I���TOs���p.%A��u���Q*'����q*C��h��^�L�1|u�U�xH���s�&!���_���p*%D���~�Ĩ��w��z�7�TJ��wY��J�Q�����Y]��ȩ�ǎ�y<9)�bTO�����ȕ��7���%�GEIWG�l�-�s;��5&r����=�;3�=�TJ��g}ZMĨ5�s���C���vz�^�W7w�n���G~��,�Ȍ%�Feҩ�C^7���7B1m�� ���CA���p]�G7&�̴֕��j<ii���n�1Aչk�
e�f�6hh.)Mp�ͩ���
�Q9~�{,7��
��a�hw"T������7�TJ��q�5^Q��Zj�M1u��z��Y����7�T��w^�M���Wݗ�j�q*@��_%�ԛ��*@�3��M���N������7���e��ZMĨ��s��O�q*%D绬�Pn%D����}zMĨ��s�_}A����ޯ^�$�+F�kY5���jUe�7�T�/�R�"w��V�q*@��������D�5���A�5�"!.%����V�P��������O����~};��*@�3�=pnD�K�h�Q�ǾGFԣ��m���\�(�r�2��ʲ��o;����9��
������I�������n@��y��v�P���z?>?>z�uA�l�ªV�,V��m{'�%')%9=�/��M����}����%�����}Z�>�p*%D�k?U�T���������/C罱k�_A��/B��5���I�|�Q H��"��Mĸ�/W���TJ�Q;���D��Q*'������(n�O��lg�����}�l����н5߽��T�Q*%D��}�Xn%G�(����~�&�TJ�Q9��Y?Pn%Ĩ��!�%d�Ӹy����K�f�pnD����(7��
��w^�����Wݕ}���
�Q�Z�5U��_]'�2�N���]�VVd���\J�P>�{I�7�Q;�x�pԨ;md�Hj����ډb:m��}߿����1'��A���Y��
�Pj���i7Y������������5�u��>Tb²�9M�k95ڽ�Ò���}��d��\J�Q>�K��7"TJ��{�4��Q*%Dﻬ�Pn!z�����?a������X��xo��L�Q*'������Q*%D�3��Mĸ��}�h�@��Q*'/��A����{+יw�ٚ7{�͙xU�p*%A�_e����*%D�2���J��v�qj�}����Ĩ5���i7 T}�}�� (�xro;���u�����TN���U&�TJ�P;|'}���Q*'����q*@���vg�n%΅����������/E�ɟ��>3�>^5�TNs;ⴛ�Q*%C{�w.j�kjQ�m̶�YPX����ªL��������P}�TJ�����q2%D���wդ�J�Q����5������OY<.((��u\j�Ќ�1�e�焔��$����Pn@�������q*@���u�7�T���/����Q�g���j�;<96�o<�н�Ò���D�3�=p.%A�s�=���Q*'9��A���TN��͑7*%G��^�T��sN�]�V�s*�hw TJ��r����Q*'���z�7��
���_}A�������l�%8O}����t���]ڏ���n%D��(���_�RnD����~���L�P*'y��i7�T��'�w����MFarkE@w4�����Z҉��k�홱t���i5�ҡBn6l	uڍZ�)b�.mn�lEJ�:�M,xܐsNW� K�2��5���s�h�J2�^L����͜[ds��:�nf�RPn �#F���ʻ̼��x-�$
�g�n%Ĩý���Eٕ�q5�k.�z��&�q*%D��ｳI���T%�7.�U����M�I�e1�ٶ�r^L�,���ޗ�Pz&D���������}����Ĩ5��Q��4=>^���~q@�3fMq1�R�����ó�'%')'���z�pnD���o�(7��
���;��dJ�P+�W}���Q�m��a��ĭe�oz���M�T�Q>�g�n~dK�P?w=?M���{߿f��PjD��/����Q�=�3.Vw�l��o30�&�dJ�Q>�g�i7�TJ���_�A�������z�q.%D���}�]>^��^�O��]�W���{J���CfV�q7�TJ��}���
�Q;�޽(7��
��=������s�ٞ n���*�Fd���y��a�5RĨ5�}}�{C����N����%�0�������Vgf%�Cfm�H����?�����*%D�{/�(7��
���_}I����^��//&��޲/��t�@�S���@��P�1	D�T$��D�"�i!Hh�
�bҋ@J�P�
5�T��(�n �JE�">LR��ow�}o��W�K�E��Ҏ���\2�T-��]e��:M+͛]�\��vU&�ƺ�3k��R��:�+��+m�����Q��ڔ#%��R�l���u��ڃ2E�TK�,MG�v[mR�(���`�Q�J�6�(�fը6hR��L�������&�(7�!����bѕ�eue��jn���r,�t�ae��tBA����Q�-�h�1���u �"��ˍ/&ٶg�%�Kf�fm	�tUFQ�ń�\��(m v�M�f���E�g6چ[�k���,3(",,�5��3.�q!�m�:����Jm�pq\��\�k���#�q&�Hb�\ѷ[�J�mp��r�X�*c�.������.+���eU�f (���J؅�� �"@�j�
M
mU��J	�@"	&�Gj2��q�85�F[2���2�v�A�1v#�*�0l7��C��Z�-���QZ�m,t5+1V�sZ�V1�������Գ0�]�)��L*dɗw�ד�7�TO����Ĩ5�v�K�7"TJ�_r����L�Q*'y�zi7�Tg�:W���d����r�e������}}�g��q*%D�}�MĨ��}~�g�n%Ĩ5�������5�����|F,=>^��}3�x���zqB�r�?~��D�5��}���
�Q;�߶Pn%A���{��ȕ�zK�/Ӹ��W.�yw��@��A�q=�^�J���퟿j�����ȃ�ِ>�+u�c���$A�&� {�O~���o�e�a)v����D�j̘a�V�C?�����({���iN���y�چ�
2��Z��m�K]-�r�-�ܺ��t�}�@�\�h�i��SX�fH�̋2�y�JFb��ĉLH� IU�CH���5S����C�s�й�t�{;+���pNh�I1��V�y�˲݀yu�_uM�hlq�q4٫6 ��j�|��C�ِ+�`g����<L�o�5n���$�1a�4�Ѧ�P�{Mf�8�\͇C������ �]f�u� ~��%X�z�ZX��H
���*L63,V��� w�Y���,A��� �qr�2DaM�T�ͻ�M:.�f������ܫ��[ x���ĩ�A�ɱ1n� u�d�Kv��~��#@ńVAD�@B��#B�I �ؤ▫��g���M���{jM��(=���������N� a��7u�{*��18�����w���d��BY�mYZKg,[�i]�Ae{���߰}�V �Cb�=���˫�}���z��'��%���ͪ6Z�fu�ؾaz���>��P�,���"���E?��m��F��a���GV���twZN	/�g���Qi�F�n��oL�[���m��� �ۖ�?}�U�Z�ɺ��n�j�ws�x�2��a�=��U_Z�Y$��٠��v!JX	�-M�Z��E�ҵ�r6L�+u��ۙH��D�ֹ���M^^Q�K��m41��,&,6.�-GZ-XM���S<	\.�l��q^���(�^kv��(ذ��y�jc�-*˪Q�#ug9s��yﴁySu]ů(=Op�M^�`wS��H�6[�u���65�c,�]n�~���<��ꤜ���I�)��a��^���ԕI	�8�f)Y���l��J��Y��:�����{����X���Y��u�M�]ZWFдۦ�+c���$a���B����u� |r��F�"�u�M��׫�{��;ۖ��\���l׍l[ǋX,q���CݽT�WH�ųO�Uz���L�<vۼ7@�߾���[ôV!uA6l���L��KtW3m�n�w�W�z�{�X��\U%�wy�|��{�?=���U#�2�+0A"ָ�l��(�-l�ue���^itT�3�:n3)(���2���P3m�� ��^֪�F�q�W��$��b�D���u%UT*���feB0)4��>`a��Xw]K x������N6p��T
�h��J�C��	/��S#��V ����wA�D��( �:v�ڶ�M4l����7Ik�|�֚���Hg�-�ۛ���Ƶ6uQ�Y%�7a|,�D�������������T�	�]5N�XN�2�
l)�wsubҬ�����0ä�%��+}!�@��u`�RZ�R��M��6�@#e&�a4m��6F�9����C�}~:���hr�[^�́n\�����d�V���f�N�ӝ���q��ЊDu�L�|��b
���[JŨ�8�a�b[����f�.:�C�� /f��Uwǉ�/�pպ��z�2�ųB�f��Y�?_\Im���l�=Ȃ�r��J!~1�c�S+��A�)(h�b���m��ib.-&�݊�km�Oyzw{厵<yv�kh�5�,<M�h�./�Ы=la�"��٧x�ucՃc�A�p��3$�����HY��� fIu`W�FԘ<l�cf��=��hw�vjX������c�������$$20��H0� & �T�4�� (B1 Ȑ�H����h�X���E� �!H@�!AH�qA�A>�ns��*�u��;�S�jRkƖ�(ˋf�.:�zِ�Y�g�+{�s�����Y�=��ݝ3���M���-�й�mҊ?��K�G�-�z0`��� ��M{�X����������|[��05�Z,z�{}۝f�����$_��8�:��vpD4ӣh�V� {�W ��X���d�� ~� 	 ��6�J�)h�u,���=��Z6:����H(�t��Y(\u��t�����������9s��瘿��f%���h�1�tTkV�3��(��aT�`�-�e��(�&�6�T�C5��%.k�Q�٢�J�R�W\*]5K���ji�r���"/:\l6#IF�e�aV˔6tYp��#7.8)����������E�32�Ch
uP�w��w�z�Ί��s�t}����qݪT�ٮ.&���4͋4�L0�@�$�f�|��k�dج	���O{{�KK�	�@uCJ��$��SZ�q���0�>]n�9Q��ꯪ�������u�!*��Y*jm��U���u� �s� �]�i�qSou�݋c�x,q��v��:���a|���*�����D�����Mz�@x��x�4;�f@Ϯ\TKG����S5�� �]�hs���t�K/
:����V�\F�P��V6��I����������Xګe���R�U�wiSI�D�K]B�є�\�0�b�c�6P����T;1l�f��T�Z�ՆU�!nV¥��V�UjK�t%����	�6�;��d��='�.`Ń.j���M�ڞP�}��^:�z�@x��}��q�qF�y���z�@;���^ڦ���,G��ۯtǉ��<2dֵ�>��zلA�A���{:�ss^$E$�7�������}�� ��RȚbR�)���۰�M�����:ם5���6���
���p-+k����P�wϟ���{��@>�Y�G\���OS�qk(��m�M0��I�ov>AW���ֺ@����/�����Q�\�ڥT:��g����Ӟࠕ'+��I9���T���;�G��ʙ�E�6�ʰJ���:�Y�i�+�`z�@�}q*��M���i�C�UW�K����??���� ٰ;f��i7�uv����MY���n�=/f�@-S˒��.�)�C��I�IM�I{rC��/��yX�x��ƚpR	#6m�4Z3`�u�����J�è�����Y�_up�] g֢�C`��M�� u�8z�����������vW 9�.ҷd6�T��T�W�^�I�_;Z�\S���؝���@��ɚ7��%U冁h�e�X]e�&���"s(�r1�H�` ���a�e�p!u�eB�I��&�*��ղ�RYe�(fJWIP`�$�!@f����T��(�
m�Vʲ��!	A���f�L��$�5(��Q�ueFJ	! ���M��`��! �`BcYA��P����B�K�p��5t\���-խkS��A��2��Gmkt�·�2���%j	�]C��
k�j��кk��3W5k �5�s�n�%��Q�X�1�c l�檰��1Y��n1����1�ck�����c�T�s8�Kq�Wc�2��cնո�g�mqQLVM��8˂6m�5��9& 5Ѵ,��]�\-9 �b[�4r�m�L�j���3�m����֍�К��y��T��3�b�+��x�1�0ؕ�X�]�8eQ�m�3^v��&�hX0����eR�6�&%64&��q��A��%�ݰ-�uR�ky���6�T��*�D�)m���ƪ�x�FY���B��^k������pv.���	�x%X䌳T�fƺZ6d�4�m�6���@W��֐�Hf̈́5ŕ��
q*�`�q�\k�l���9����نU6�b�ZԎ1s�J��l0��cM #��i2dJ���ܭ)r�9q�Cf��W]r�+]q�.˝Z��v�q�Z�]`���)m�YkVgY pjn"
�v�S-k�3P�h�[b�� t���lK�YR����gM�q�)+k,WF�ZS%�j�SY(l��b[tqJL�mB�bge��B���W�3mR�VX�9��VYv�0��Vh�#.����bR���0ܚ*QF������&]�:� N=U��"!�-��;O�S�h:��6���O�:�g�ԙ =E�i�����<��,6a��p�] �� �z���.�?��~�h����}���k~~3��a�5vn١�X�W��Zm(��4֧��֘c��hpZ�A�m/������9��{/�&�Yjܿ,�i�t� < �δ �vZ�%��@��ÇPJ�����@�`fk���W��#�րȪu�=� w�sM�����G��ȉ��m�Ű��D��gZ v�ք��R�F�6={�,�w��W��{����&�n���ӎ�KxFV��%
j���ML�F�.)[Q�R�Z:*`�`���٬����kB,�r��uF�PÀ4K�h�[t�sZ�RgZ�.��C\��s�R�i^�6���f%�i�!��Z��k.�`���
�xL�(D�4"�Y���{����H��D�n@����	Ğ�h,1f0î�g�QѶh�P`7A��O�̐�3W��HlC��$\�g]ҽ����1�.-��D�7���l{�0/�Y�}�d�ΐ�]v3���z<{�l�M�F���V����Z6>�`�Z-�D��ƤDպٻ}�@�
Y��;L�@N�u`W�J���n�WL���GV���#�`b����ܶi��խ�[��G�l���}�t�$��4��4���``��`ː�kWq�L��?�{�{�`�B�G�5@�A�wi�_!� ��*�JR����n��YuU��ңk�����CM��
�i������31�1x5 Cj�cFkBA��kQ�fe.mf��sG��H��#�q���;�F�=FYR���,usMCx���z��� � {^�����"���[&��E�eXvZ�]�f��]���H��b2�u��lQ��<r�Z���4;����2�����ձ�Q-�4����,A}���r١�s��8+0l��� �5�@>V�CZزå0]�U3,e�*�KTh&���-�S+� �@��1^V#�ά@�ᱭ�7ty�6��5�5�ن���������բw��}���l�Ƒ��ŝXj��UY5�>��w^��v��X	ր�GR��ٴbl�[vSw��z����:@=�f@���H�-��n�$hںJ���C`n�C��,A��H��ǫi�A	��ޯ,@�ջ�	�CY�2k��dQu�t[�ùJ�����qO{��w�_WH��D<qNݥ��6���9Dw6k+%MP� �%�����C�}U^ g*�2W 9�.ջ�m�Jf��ྪ���Fր��]d�#�%f�i�x�G�7p�5����}ΐ�@�bҵs�w��$�������ef��ź��'�=�}v� �s�}y�>V݁��B��ء����)�{�����>}�v�mMMN��MR�F^7Kri��f��﾿��y�ޮ�3�T�����M�?,���lՠg��+����x� z��4;��}v� ����v�$�:j�wF�VI���X1T���K {5�}��U����Ք��O[Ɣ��� ���nu��ň͑:4��ۺ����n����rK��'��zjI��{z�k�� �!gڗ+w��Emy�J13]
�i�M�V�;
;
��;V�V��"k\�,4�\���K,]06)	��h�\�M�j�L.T�6�Z\c-Mv&�̂Z�ճ03�S!���t7Q(Yi��3���@`#SaK1���\�j}K꯾�6�Zc)��ջEm�ۨy���n���Sd��e��]�5K��ڎ�\������ޜ4�υ����膒t��|��{SX�u!�ėhDD��4;��}�� ����?~��C�>N�0Z�����i f*�����Y6> ��|Mf�M"gU���{}������rI9-�V�d��X�l ��7v���iRB��UTw���V �[�=��``��Q��n�6nn�y}�� ���.�c���%��:Qj��M��3L70����� �۰�z֤���o/*��z��=UC�		PE
H	P$$�
�)�BT$B0BX��$HQr�$$䇑��J"ݞ8t�t.��B��(�&�gYX2��r�
[�e(б�"+-�Z �K
�˖fW�\��][�m`�B ی�':�w�<\�͒�ì��'���tuy�}���ΐ�:�2�-���)5�7I�p�] {r٠{d���p_礼8��I��������=v�(^�b��b��T�@��a��P�:��.�ڧ {#���[-
��(�Zv�{�\�t|�t�R$bն�� ڃfձMb�*�˭�%�n�}���m��ܬG�)�.&x��5+u�-�R�4n�0k�� }�t�u�Hʝf�����f��(�ݴ��S-3`b��mbB��4�7�{�RO���ԓ���}�3�g�i�n��F��T]�!ؿ��x��ΐ^t��
��mcM8H$�-�H^�{� {s�����܍�5����� ��ﻃ=�e��gki*�Ĥ[���V��+e
��}���y^V �^V#�.��1'7d��-*n	v0,�1��6%�	uz$�V ����86uUW���X'�Oǒ=ǺG����:@/�� �D���Ѳ����gF��N���+Ԭ̩�'��׵Ro�ú���db��",`4� � �@0-�:������}_N�W�SlP�!���� {r١}�X��:@�nqp�ŭǬNkKt��������α�,�g�ɪ�2��8�P��KEM�Џ�NO��p�������R���H(�t�	:B����d4�7�JW%���b��f�޶d�nu�w,࿌l#qů[�Kb��?���ʝրâu�7u�����vB��,���4�i����Azِ��b���OՀ�m��8��{�����hw��u�H����0/�`���sjgf�F��A����ٚ�#�4p��J�35C]��������6�iui�,x�Fmmh�4X�Z�$0�u�:Z$����3JK�&���3�4��sJ���j١vL��-��Ae[cc��T�r�fp�Z�NO�'���'<i�����b�*t۴�,���wɌC��Π8�݆ �M1�О��0�}�?�������źm�	���ݍ6�a���h�v�v�M��e����Y��u� �۝f�|��3�e�-�k׺F4֐\[?���T��B����ުߺ�!�dQ�%�z��f˫ x�2��'5T�@f�]XEH:*¶�RM6���'�δ�|,.�`.:�;<�ׯ�ůf���M]�~��z@4��4�;��m2$�D��Y���
��&�|���� +�`S�Q���"D�g@�RPqI!	 HPZH�PB�v�Q	0 ��@�Ȭ��E$��F�)���4��S,0XU˶a��m��T�y�U�p�V���)jFA"��"5a,a@�*��*�%%kF�Th�j��HIA�F@$B ����ŀB)$���(��E� @�#�F	 ��dB �dHD� F,*��"@�S"D��#
%�((h�$�A*J���	RƔ�H����$`Y Ū)�41	 �2�PE�#)HQ	L�`|�dDu7�5��L,6�+&ų0d B0�*Ԗ�H�H�I���v�L��#*P���$�I@PB��$��A(PF�%��U��	V��5M�Uq`PݎQ�i40X��b2X�[�"G���+�+�S;.Tr�­�L��%��5�F��c�7Z9�%��UT���4b1]�m���H*��ک)F�6�[j��ز�v����lnرV��eڬ�!@&�.�A*�kr���-�\��nm
!�������D����P+�H��Eb�Q��)��m�\K��3	WMN5�&����w	�d"��LY��b����u�����W8,�D��+�IEi�3\W��Q&�v,��A�f�*B�	PQv�U��ҮP��Zd��*&��Pڕ�CJ��5mʡ���Q\M�!B��T�(�����+��^<l�i]m9�80E�j���nV�FY,�	m�̲�[ce���0x5D`�L��cb���w�����s�y9�G��u���p> S�s��>��}����s�SV�ʸn��4����c�cr�e)JƆvL���Vf�L�9�+n�Qs[��t�^+ʍ��T��uE����,�w��Mj(�U�ٮ���Q�ށ� �)�ó�����u`p��Y���=��=K`.:����{z�ݹ�i�� ��_��܆=��@>W��-��4>�t�}��gݝ����<��'�C�l�.�`v�Y���,G�(iq2-��dx���������-!;pdm���3M1eV7f`3uk�u���ϲ�Lج�U���٦�)�-?����y���]/u��f3�X�4��-3�j�l 3�@nIu�UW��3�X�qh�����_WEv���j��r����$��9�\��u,��dJ�4�.ŻE]Ӱj��C�s��� /�Y�}�Eh�x6Dۂk��ު��T��#����k�ք����I�W�.�QIw���Y�h`d{F�*R���ūs�2�b�.��ϟ��v{z�ޮ�/����䉊n+-�m��tǴ12�q�\� �\�ِ��b�z��Qt�M1i۲�-�db����[��� �^V#��j���D6'���RM���ԓu��u~A)Љ.{��jA�>�D����vEYl���_}��� n�]db���U|b����i��<�N$���8���١��ڶ�&K�]Z�V`hmb�%�Ǐ�lI���{��u� �x���O�_�L�{ހ^jy��bh(kI$��Ǣ5��=�w�� �z�}�j�w���r��&��#M6Y��د�������u�0��jڠq�m=ȶM��n��>^:� nlv:���&ouՀ0�=d{u���+V��*tذ;���뮲j��@i�~}}k�󣟌�L�f��ô��g�X1tS`���Ul�b��WmP1f��E
0��٥�48��F�kf��2�m�h�0r��t���ʚh���rbڷ��c�&���,p���ib��i��e�Y��l�m�X��8�U�W����̪Q<�Os�5����Vۭ֬�v�{���߯@�NNs�|��5�L�k��ƙ*(DD`6��R�����_���F�����<��>�Ç��5'Dt�p��kv��FX#c6:��������b�Y�{s��ߺ�ѰP�65�z8{� /f�,�Xú�@��<݊1��խ�&��]f�zِ��X���X�ʭׯ�ůf��bZ�����hr�١��H�ųJvZ�/͂!��M&4��� ���D�V�)vn���`5ڵI2YI� ��F���Itl��Y�2�RLY���63?~zh����\(�Sk�H��J0�݄)�a���uN[��ٶ<&&�.[�+��J"��C^v��av�n�Y�L��Ny'''gS�n��V+cI,Ѭ����+���̀{۝f��f�r���5�5�I�� /f�,���z�@>\[?�߳3?5���vU���l���:��ŢY+���f@��4��o1,�&��f�{� /f�ي�u���_�����v{˙\'@��}�pu�L#��[	�[���H��F<i�n�ٮ}����Y����/���>�;i���"�t��b3b7^���y�����@��2מX�ˎ�C��H�ǫ��AE2�*��7�9�M���t�@�0 � �� ��� @.�!E��;t��*QK�#ca�qw�S�+;/>�������f���R�x6MLC�蚰�V�@a�e���神����?���A��qF`�����<���v�nu�����V�7�$K���Gt/��w[;۴���VU,��96�e*�LWWH- �wu<��P+��x��=\���A�mD!�������V��kFڀ{��Wf���,A��]��޷kM�F��Y�4;��>]n�>\u�^t���Tj�5��b��<�u��!��?~3�!I�`�D(JEi�
 ���٩&득����._k
/,�vM���;ꪣ�g+ dU:��̀|����.I�bm�$�>���Fk{3�Y�v�s�1M���-iR�l>~����*�l��u���.&��d�Xb#u5xj0Ϋ5&�vj�l�F�@nGR�9�uW��}�ES�$�AՕn�i���<d������HCS�:> �-n���i�h�,.�6��������}�:`�h�u�F�P�m:F�@�i�l�z��� +n���͛7a����qmtw%	QL�\�h�]�[kT�km4�ִ�;Z�ٱ�,xk^5�lЌq�ʵ%���nDrfR��Z��Ѽ[�91	Q��]]�8��j�4RY���n�W����b��i�`G`&b��D��(a��V5�Ԗ��NK���UU�e���P��4��f�E��<�����v�ê��
:4���1��Qƪ���?{���t�}���_��q�Hz���MC�0pjE��@���|�n�>���f@Ϫ��n�$Dm�o\��w]�z��U��sb�6���TSVʰ)UӀ}���]n�=���/f��Tx�6�j2i06޶d��A�� �ΐ2�RLY���6bOr=�P�{��
Z�Y4�/b�kI�r岌��+��0�#������ybV݁��b�k�8lw��*��-��j��Q���s�[f�d��a���,hfۇASU�e����Ҏ7\V����<z��	����q�"mY�KQ`��rNMj��j��;JE�M�
�����[�}���C��T�l���X��+��47����"ם ]�f�����G�����������i��T-`{�Xs]K x���հ���4�:�#ݓ�^4@>^��w��u�H�s���.���o�Y�Lx�� ����@��RX�4�";.�8��"]v�ո[4n�Ay|��~=�oU ������z���8#��`���cX�\a��������w[2��V ���v�R����(β��<�O���vp9$��P"�d!�P@�b�$ �()(�A�d�!H���$ib!P*)H @HB$ E6 |�:
��s�j��{����H��T=�6`���� �����Y��nu��́�SǸ�E"�jk[&��r��t�}w-�^:�<uʓ��z���7��=���ܒrn���Ͷ�*P,��RQb�tɫ��$��eN�`l��<tl�>̒�&[d[w?�'9��%9ݰu)v���č�*�E0��w]XشK a�2�5���.n���F�dm���^:�2K� {u�`5�_W�_Y��I�'d�l��I� a�u�=��ZT����w�m�{\~X�a��������%B���H��MϖQ��bO�H�%���F	���� RmJ�H$~!JJIIB��Rʅ]�ۼAp���`�Ym4Q(HQzH~	d�"H�$R$� a�$P!����y1x��0R��W��[�e�Pfuf�Bf��v\2��F:5kkMF+�sC+�+bmbKLȎ��� �@ �GZ��P�t��1!ft�Yc�)q@�q��Uq�1�a��1�c�6aQ1�ccc��.M����1�oxj�1�c�A�hg+���f.΂֭ldљڌ�J�,mڹ"&���t�m��E\�����sv�����I�V�40�GBPΐ��su��V�	[����!�-�Z���\C��B���h�f��m��l����5��
R�f΍zt�m'r�F[Zڳr�#j��if15-I\@�ZDd��Z2��pۯF���L�P2.�2��Mv,R��	��óu۫IY*�CFR���a�nQк��Ї��Q�e]bV�dlp#��vlukv��`%.�F6�[��4�3Y*�����D�U1�A��Z��v��qT�P�֪A[�b�V���ivj�E���v�����u&ee��W(۝^Gb�e�iuMj��u�U�ծr��Tє�*��c��D�����-��ck���LX\DP��6�c�]�e۳v�dh�v3f[[��b��b;P �jT�µ�.��Ld0
4�[�Ӎn�PJ���R!	�8 � *����0�+5��lv�w�%cyZV[�R��p1��˜#].(�9����<(*b�u�C���"lB�:�`(�(/�
u:"A�H��u���7�~�d��v�b)����$�rb���y��nu�^:�zِ=�Z���h�6i���u��>��j�U���I�`�� -m���o>�ߏ ��-�]�f�{��F47�nș�MF�Sh�MF����Sig@���� �{��:��,G�+�����&<of�zِ�:@9g[}y��7X޼��ٚӚ]�f�� zِ�r���.�螎<���0���U���[2�$�|����c]��*l@s/D`Jbg-K�n�ZЩB�Y���}�WT-ڴ�����HM� ����fD��A���H�5%k�1MCm�lL�!E�l��hL���Zd�&�X�cxL;J�Uۭ13�C^�5m�m��]�}�Q���h�|C!Z�T�lzԁ��,A�"�V�5n�1�Y��ik�V`!u�a�JJ�Y���w]�u��4;��}V]�y��B�нR�+��f!k*DZ�V��d�ܬA�X����{*�n��װ{Y����z�_ﾪ��FE]ր�Pu�!݊��0���l茚Lû� zِ��X���b3�Ԟ��mn���5�q@;��}�� ������4�ݢ�k�qFcZ��Du� ��#���Lj����<*,���fU���q	'�_�qlо�H޶d��ҦT��fKq� 2D E!B��	�h ���II R1Đ#C�JaL��HA ���1#�1X��x"DK�#D@�"F0!"I8����7���3	V4�ՄjZ`���.�3�ٱ�̺0�9�
$��\- �j	ԺT�#n�Rgb����. �'w�Iяi,)�fӴ��vn���Q�K��+PˇY28,��K L�;����#��V�ֈݹl��ۖ��j�|�l�=�J�֭{��d׍j�}�f@>T�hu�,A�WHyvW�[xܚ��lǋv@����t�}ۖ���Y����m`�a"!�gl�/�}�oo@t��qm���B#̥��n��h�k-L��wS���H�ųN=�mK5��4���$�4
�\�`�ei��M�x���] ��@-�O�?g���7�u��� Ra;�5t(�]�<d�uC��ńF! X(�.I��gک7]�oRNs�ٯ �W@MS���m"�l f��`pIk���wy�Y"�l�b��i��l�a������W�޺� dS��<`�z��������G&H���ws��'ugs-��t.n&�!��A�U��v�5sc����~=��j�r��i��ꅺ�תD�Mփ�R�@,s˥t!��)�{��V�`���:�_U}�E�l�G�<MN�رe�Yw`MZ%��}_"0�r����8/��羽(��]�ʽ^a���$�rwڹ>��٨��|��^�u@/���Z���y٤z�ddw�}_Q����0���u,�����`A��d7VRiZa*6 ܏�w�;:׊�̺8Ve��� ��I�mTZo���O�ߧ�%�3#��٢5A4�l��﨔6y�F�kK���c�nƞ ������Yڤ=�����	���m:Fڷ���d�������� v��`b��nH���[�f��z�@=w�_[2��#;�t�4l��8�� |�� ��wU'�_guP]+��a+A���@.���:��*K6�u*�ʊ�J2ݥ�h�q��6�..Bmcp�L�f��͹��!�e��%0Vٗc.��:l*�E�%K�vqJ+]�mn�:�(a�:�9͚�H�X�Ku,����2kP��e�3�vjm7�.^�c,3�Y���Wƪ��'z�
уB�:J�}:��z������IIzi�s��V�
�m0մ�#�1��z��Z� ���i쫐��c�a��Ψ�]�bԃ�V ��hzǐ�yb�:���`���1Z����[�G�aݽTޮ���l���vw�I1f��dnj������C��2}^X��ųO�h��Z�[?5�jJ{�K f-��a�?W��Q���`h�J4^���\�����}�^��H��p.��ƣ�07DR��i�)�VV�N ��%�&Iu`��{>ˣ���6�U-W8�ni]Zj� t�!�iX����.Ҽ�M�Ђis	v�jjb#��r���md&2�-�Aծ��ۜ�s��Y���ݳ��4
F�A�Qݹl��z݀^� ���#=�M�o#�0��֨� ]�f��[�z�@��h���Ĥp�60[���d�] ��f�ˋf��*kՃ̈́ٚCqk� {�Kz��Y���l��we7��l��Ln��� b�f�OD�����u�b�1�+j�"lRZ�����:������_WHgv�n=p�,mC���ڹ��5(�m'B�F�Zn˫ f('����� $Pu��8��L�vQ��lՀ=���m��v�Tjj�;�Xws���Y�U�A��=dOT�m��28,�F�]U_}TH�{��t���qh�i��Ѭqv�b�f@/��<��i��Z�6�6�Nb�" ���hd[��!cE���l�����mk�CGo�֪ut�|��i}ۊ�z����%)����ҸS�7j��Ri��f@>������?���[Θ*P��s�wF���.� 0f���d�㿦�ݹl����n�#xn���hUl՗�?a��H��1�"���V �*�hA��!1e'IZ�V���u`	�Բ-����z�_�=��xި��L�Ġv�C�i����(�:�ci i�KaҦ[h��;�`�j�&��.�N�e�7�5D���bF=��6�����QfU'@���� ��X���d�� ~�UV�'���Y�T�0������ݹl���,F_��!�fǎ6ǭ8��X������'5N6 �U�h}!�!��m�^��<�{�� �S�о���lXz	@���0F4A����8��Jo���ɂ����H����E6H�-�s��YfR՗��kDsLSm��h��]�u�\b�T\:�biz��e�WYb\����n�W��n����h����]˳t���0+��!��9&f����F�i�iJ��yXXFѩE�l�idh�xHz̀9�տ��#	Ca��4�\��73��Zś����U@=�١�ΐ;�V�?nl�W�9Z8٭2�h��nic3t���l��u� ����>A�	օf�D�h�HݷhڦXV �͛ ��:��f@>��@��jEFksu��5)��ΐ�����l��u�������oV�.-� �͊�諭��u�hIP�铷=�.A�@���נ^��8�2&P��^tl+evp��ceD�%�N��28,�[�Y���̻��5Z�G>�4p��S�U�Xc��BU�#`ST��4M2��ѥ�FAM�9G�	 �d��"�@�#(F_B�EE��j�@! ��F�H��$g����1�P�1�!��-'Ґ�$���PK����J��h.�!I�0`H@0�2(5P�,b@�#!FI"�;#�0#�,�h �J���K@@ri��Ti����;���y�e����Z8�4��������A7mu��sLn�Z챹2*�i���k��]���]�����JUT���ʂ��J1ʦ�v�ڎn09����LhR��dѪ�V�:�Y��.!�T���t�[�!���k7)�mM�t����5��t�RX2�ftة�If�%�Vd�4�ϽO&�%�^���Sgb\F2�"�i�ܫJ �Nq�CYj�U"F�q��&+6��"1\-��M�̑g�<a[O
[6����5�.3 ^v��R�sW*�ݱ]�c��]�f	��R0�*iP-^&ib�{p�3�L�6�C�+v����F[5��E�9�b�`F�b�WFƔ�4Ə	J�j5u̮s��b�x6��\4� ��@����`��+�^��Uw���`�)��
���-u$k���2����4�eF��ٛjb�Үi�P5ð��-�q�,�+7(�W���Һ��MT��t��N�?d�q�E�e�]4жV1���*6����,A�WH�u��t��]�mO[���A�ݹlз���] ���[��u��͑l�,Z�8���4/���w��=�t��;�����l�M��Z���@>^:��mP�f@�v�`n&�[3E�������o��|�L��hA@�X;b�2Q��鐎��Y_���?{s�����Ԩڞ=a&Ǳ/�.�uۋK�l�A��O�s�r�v}^X���Ӫ�����u�QY�@��~��y99$���h�@û�$��}�W�O�N��e4m���Ba�@i��`	��Y1V�@a݊���!�[,�n�wI��6}�Ţu�3�q�͗VU}_Q�뮲;y|{^�4�DG�5�y�$�롲\閍 �I��J�Wk��`�7R��}��4;��@;���~�ϡϐ�{vR�F�+�Vh�Hm#7G��Mv�P�� �x�4>�@��F�������B�{��>W��-�H���~������9P�Y	�E����a�lu�d��;�_U�!	!KBR$@�BTR�$�$R���_�꯬��&����(�&�2,�L��4>�@:�� ���|�U���P�f�x�Z���'��nu�	��z;v"]e�]�钐 I��F�������w}}j�=�� �U���6P$�ڦ�e*�*�N\i3dqz�߾���~�$��T�U���Vw�'!D2�s�m��|�U�-�d���4>��f���������Ml�d���4*�[_WH��=���Zړf4�4n�@��2�m,A�ܬGٙ��BL�@:�摒�0�ˢ��*3k.�h*� �1�� &���+(�ͩ�U�C-�1�sl�يO��ނS&�9��.+���h�@6�k�ٳ��H��gSU������s����p^(˰]Mmwgi�j12(�ͭS)�Ii����I� )`��}�I�����f�0�a���<��}��NiC��,���<����9*�.k��l�VZ�7V޷��w�:��[��A1boT��s�rr^��{v���CJ9���2��h� 4��hj�������{�K�.�
��-q,�SJ �l��^X��ųC�ΐ8=�IcCpo&��oQ�@������ĹQ�h�����J�LZv����yx�49w+_[2�s��uM=y7a�8Ɩ��t�n���̳c�W9�,�CqK�m5M�պЅ�������\[4/��O��b��m!��˙�E��J�i�+]N�:T݌�T&{GiaD�8뙠��ٶR*u�:� �6�h����Й�
�2�`�ɛ9�$���+næ͍Q�sfH���|��hw�����~Ϙr�Y�L��*�Ӵ6X3\���H���@M����a�3��M���8'�l�/��y[v�n[4/���������#xf�� ��2�$��f�,�����8��7�S��fw�n/sv%�߷�^�M)��n��`t�-�f F�z,Ы)�`R�3��@l�R�d��߯�L��9;oNӰ8Jm���(�%��I"&�;`L��0���١}l���5�ת=��Y��Ű������~��yb{z�ˋf����oZmH��n�h�y[U�!�K_���{c�`;9X�~;)-�8�j,#�f@/s��ųC��,G�θ����H����~��o�ww|�3�FaQ��l�h.a�sh���]uկU�{�� ��<`�Й JL:��hL�rHm43IBWD.cr =���о�d�� Sݥi��F�ǩ7��;����ڠ.�`[f@�rݯm��X�F�/N�M�g{����vjDl"�Z-}C睊͎�rTV�AA6�N��������,A�m�g��=�γO���!=�x��b��ِ����=�@,E�J�%�]ss#biukX�$.&��������vo:@�����4lM���ź�mV�7W8���G�~��E`	���}�y�w+�����Ԕ1�4K^�8����4>V݀}m� �/Ub=��Aq-mIh�c�[ΐ�]f��\�}ΐ>���d�ц�5��/&Vf�yU�}��RN��I��s����A5�n]Ʌʴ��t��&^;�͗k�i��
�,���a��$%bԕە�b��G���6��Jm6a450�i"�L��a\���o�+L��6` �[vT2��S:���j��7j�],���s�M��ii�9\�g9 �+�]_=z��;�Y,�˚�fj�ǉ�ؽU�$S�16-bƘ�I�.¨g"Cf�ָٮ��w�~��H�]f���
�7�߽�:N�>n���\R���R��Y4π��@ò(g����T���ᬛ�׺��vڠu� ��@{ָgrZ�i�&�?-��8�]f�޹\��X���H�����ɻ$�竤�ųC�ܶh}m�԰]V�V�{�d޵�zL?=��]�v#pS&���[�ĒXkz�[��s�=��h�f>�}�΢�[<����u�X2�Y���f382ցf�1j���#�iL�5�w�v^�L% T֎qu
靋R�&u`��̌ئ�͂.�&β}��${�B���2gG��է�1��<l�pZ��Kla��t�yx�i����q��n�q<�0��2�^���v���3(��8�T:��D�m�-�h�z���� ��H�[z����&&	9�n����f��s����ؽU��[��LoY�Tx�y4-�N�;���5U��]l
(�R��J��>�~�6ߟ��4/���hkm�7e϶E�`��K(�W�b"5���z��m�+��2��E���@^*ݴ>�h�,�V��֬�ԓ��wT� ��0@)���`��_��~3�(06H�	5�0�����] la}S�rΨ��� �D���h}�f@=��X���lE�@.k���Mx��Pz��`,��(3[�W2�XdjJ�ڤ5�Ź�9�.���Z� ��́N�+Zd�A�����9�XJis�]����m&�IH��b/���Y���2{���m"nG�Y � ޻bw<��] ��Y�ׯ�u�M���MbxD�Y��:͹�b=e�H0�GP1�B|d�dP�a���,$�#���tsx�Y�a
�IL�Q������c*�L$sssD��a�(��/��mJ%^�Va&�4�i�"F$C�1�B��,"$��U[�	"�ٖ�aʕ	$0�XLQ�M(F� �#"A����M�@��٢��`��vHC�	>�
M��8���D�	�P�4E�"ޘʴ���`ABB�[*�a���r��Ր���$aE�
QkB$haI�PB����QKj�kw.��P`� }���E�H�E!�nU�.��4��!8s��ղ��l9Q�\E��Vں�Z�� �Fj1�չ+�v3�i*��h��-M3������&�[@�뜴�-�DMS��j�c-sl!�b[Q4b���65v�b��1�c��6��1]�������h��1�TLc�0�M&���.�\;m4c��\(e��Qn�Sk�!5T�v�j���&e��m�B�Z��e��l.���5�Jћe��+9�b�LjfX(�֛qFZӈm��;H6�c�+]6 T"W6Ya�-�жv$�U�#��ɣ-"���,���3hČa��\�aj�����[�.�&v�L�MIBQ�f��Y�F��c��J��e�aj�Pc�����Re	l˔��fm�m�)+r��ȫ)l�T�,��YX�*�²���p[j�YlB!���]4�����\74b�`�&��jZ�5vƶ���m�WV�;U�cJ�[sKr�-�m�6768��eö��k��9v��a�
9`ge66�4��bR3(V#��GcE2:�jֺ�2�B�M,����6Ə�%i��� ����/d�`�X���A�nԹ�B��� ����`�R�`���.�T�%�+���� ��.�Tkh��!��er�ZᚙԬ��R�^�(��V:�����a1d˳.�Q �4�v��5��S.m٭��j���i�����PG����Tڠ�~Tt(&�L"�@�g罼��+n��֫��L��CؚQ�ם �s� ��lAo<�߻�Ś=6���ǫ`w-�C!J�w<�X$f[��Jl�u�֭y�Ǐ^6�/�e��̀|��}�d����2�ޯ�1��#�s�X8j��/�}��i�����@��|,�jGQM�w�&Ѻ�y�;�� ��m����}�ׯ�ԛ2L��y �q�hyz��C�m��s�Ҟ�7��odı�m�=������y����~:�I'h�����y��T�+Y	�Y��!�2�%�eڶ�:l%2!�@�	r*��������L[F��h���1�����B���SL�ڛ��2%n��f��Eچ�̆�J+��q3���G\Ϊ�Q��cep�,�]^\�ʼ�y����Pد���@�;u�p[Cm=�sC�^^нv֒��`�l���c��B�p4Ʀ֎���߳�m�}�Z�KCD:D :n�����'�$�av�
���P����)S��S����2�8, 3�CպN��פnLŰkI�s���\�^X���H���q(a�H�SB�U�h|�݀}w��}y��`��Ŧ�R~��ۈ{��_nu�{�X�˻k���wF�f��B͆����HsM�Dš�ԙ���Tlh�v�.cGF�,Gޒ/ !�*Z�i�F�� �4�������xث�n�71sLW+]m�5�vmC	*��K�-Eڙ�&�VPvÀ��\�g C6�������aV-��l��8��\3l�*c0�1`�Prn��\ ���Y fl}_W���]ֆB+�C��J�m�-Ր0��3]H���H˺�uEi�x�[Z�׻�����X��T�:@=��,E=�X��A1�����{r١���ywmp�yb?}�C[m<SwdÆ�y����ת"�Jj�/-�T"$	l���&��6�B�[�M@i�2��a�>ܐ.�=}쌅��m-�E����CW����yb���w�-����u�Q#?���a���-Qa��gu�"�'Q�+'5��ԓﯝ�W��4�������5dC#dpX7\;磌羽��]d�9�\�.#X��)�V��s�˻k�w��{����V�3Y"�ݖ�5�_�o���h��.�[EE�6,�&
gkE���0�6:�@ٲ��̄��6�7�T���I�$ŻU�ԡ��(����{z���H�x�4���n�I�E���kb �:@�[-1E�<rd}��2U'mɂ&��ï:@;=�,S0�߷��~j��S﫝���_{Z���+�7XV�f��l���_WHz�@����?b�y���ȿ�3Q$��hC���������Sp�Y��1F�F�I�Eu�.HA&�LYv���gݡ���竤��rH�֔�'7�
�h��mG�cy\�s{��m������u�;���uz���7j���N��[/��F���w�Y2:��_R<7�6�j�%�m��y�Y n���R {5�a�ڑSX��QDli��q�z�@9�s�RM��wW,�P��Cs[����-İKy,�6]f�˗]V��l
:anu��v_��ަ�U4aw4�9���F1�V�P�B4ƥ��.F��ү����LGi6I�d�7dQ6��e�L�r$�k
�j��]])�!6�Xan�������E';��I��r�ja��y����U�h~��>�w�������x��Q#v��0��%��]��xų ���.{���5�7RR�1�kt���my��H��ku8��H�%la����� gZ*�z=���5Fb�ܮY��� ���z�䐺�Ŧ�6L{��@yu�w:���d���4�rλ�z3T��$3TG���(��z������eK@zk��ښ��9צݛ��h~��}�]{,WB�Xl]�&�:Z�G���囂o�u�@=ˬ��ܶi����N��U҈�b��:�¡e�L�R���Z�ci�pS"ٲ�\��Ϊ�o9#mk��4��Y[��Ն`����3��!
����Gr��]u�v��wM����j�[Z�=��2���h}�/�� ��[4�TV�8-IH��l3f�ם �<��<����ubY��56���&�0�ܶh}�f@<�.�C봱��C[m<SwZ6h����s��@��ր���3l�?{։S��$xfǃ"��nu���j�C
k��,Θ8<�uc3���6!�~�����߻��l�p���f�l!�	��`h�V�Tڶ��km��_���� ]�f��+�i�Ÿ���
�Z5S.���}g;�
 EШ�駻�X��[2�ܬGwh\Ik��,Sb��>�̀y���[4/��٥i�5�)�Q��ԇ�W�U��u�2G���a�Mu,�a�}�ev��u�eN����۠s�r|���B�$��X9�i]�,OůĊv�"��E$��+�D�,#�\�\5�b����妭���qlckN,�Wu�|�t�mP�W,���������NF�&�Ln�n[4/�� ^�URZ�`��Ⱥ6t��*�Flw$��w���#�0�Qb�N����/3�5$�o��H}\��f�I�[1%�0���{��@3Ih~���h��2 �ɱn�5Í�?}��w e%���ff�l�����ۡ^��l-�׺�G���V�>�um`����sҲ��Z��.K�X�]���붨j�C��,A�����6j5�{"��-�1��\�$�͋�$���,�O��=�%���,Œ.�i*e�$��{��IVݙI{�S�H�{qCW�U����U2�t=�	�.� �u��b����I����W�Aa,��i �5��*B4ڸ H��!'���ԩ��u�VKm]�.֤%���j-,r[F��5��F\�T��]n�L\��K��t�5K)��4�RU:R1utF�ՙ�VĴ.��+�.�f���3 A�.�]�����ٖ�ș�*�<��2�\B�ƒ}�J���\W�NP��Rj�(���)���}�����ް)�Q��4�7S,�qZ�������hЕ����A,�ESN����(4��qb²��/��f���$�s�8���Y��N*��d��!�EiꊑD�A]�Z!�d�qf��uS(�7\mw_�$�ȯ���6�A��	��>��$��~ �����$�K��"Hݕt�L�u=�Nш�HT�FѲ�,�-����UT���x�{�]аI8�l��=�}��}K���;�Pt���@�K����>���zI?zHz|��D@��Q*�� �-��cR���{��I'4�d�}��y��$&
�_�  *�� _�  *� �������W��
��
 � DP�����
�P��`�D*��X��`�A
�D`�D
�@H
��`�@E *
�A��T*EP��@*`�A��E ��*T��DV
�P*A��DB
� �A"�X*��EF
�*��* 
�*T`* �@D��EV
�`*��
�P"�@�*D��D
���A`�A`*H
�
�"� *B
�@ *��
���E*F�
�Db*D��H
� *��@B*���E
������D * *��
�*
�X
�"*D��@X
���Ab*� *�"*H
�B����@�� @�"�"�
� ��EF�b��X
�X��DU� ����U����V�]�
��� *����������W� _� ��� ����b��L��zJ�b
�=� � ���fO� ��@
�� "�@  ( R��J �(
�  
�[�              �            
              ��  ͉��ի+�k���u�-��Wv�;���O/___n�{�{[�]�q��\���zkՙ������ P  �g�S��n��j�r���j��/�]z�ֻ�m�����u귲����s��{woXW��m{�m���  `  D�z��^�{��ݳ�=���x�u���v�v�t�Z�휽u�uu���^�ò��x7�W��w�m�ݮ�v     �]�\췇��װ����*���ګר黫�n�-\�h6�;���q�k;���x������� tCs�νdP�+m%(R���)K6�)JV�bԥ)6�%(�JP����,��JQP�&R���QJV�)@�@  i[i)J`kIJR��$�&���fJQJ���,�d��*I��R�V�RR����T��)Vm���m    �e)J��Wz�i���5]��L�gvڻY��]y��OsV�=�u��7k2�����ux��  1�=��(�]�ݷ��)�]��Wz�׭z�w��փ�\t:wV�V��׵�]�xz�Swo \  ����ۭ�ӻg������7s޹U�un�.���;ٻi�n�g`ˆ��[]�KKe�      Oy�G��Qv�۰n�t�ji���O]��m��k�`ܻ:�׺����{ں���[�u�� �LԒ�F� ����R��   �В4�� �'�T��Jz�  T��6T�*   Ԕ� 	��<r�9G��NG�������l�3��DKt��
 *�u޳��@Wb��PU�����ʀ
�P@ES�~a��ȅI����f�$�09�IBHZH����
f�<.��>1!\fi��9��Şm�"{�����B��ӳ6����O"������� ����6|��4m<|8xO��{��Di$�� s�q�H�>���a�!���H_�%�M��}�B6)5�{��2	���L1+�4�S`CZ!�����K����I"H�@`�AS[=e�ٚ|�SE���41��)Ǝ�U�H|y�1< l4c�H��5e4����4ą�$sG�F����9��JS�=��9�y���(��Đ�#���4)��f���8@6��Yn`�5$&�� X�r- ]�9\IrVI�[�7��ÐA5d8�<|�ս�t�Ȯ�\������y�0Xc�x����#/��4,���d��qڡ�E)�M��$��&xs�ĝ�/*Ą�t�qyឲ,�RW7���c��'�p�b!��K�Ȼ|��|�טs��B6f��9=�u#P� [�_f����0����3EHF]�℅cnK�#B)`��9� I
a�\�C�x;�sＧ�	�A�i�J��
@��XB�F����,+�-!T���_Y湴��1�8�0���R��1��BA��%�I�Hb��6Gd>A/����PǞ��F�#4y<����Bp�4l��7��XF!ѣt�'�"T��G6$�p�6�;|��0�
�u�xb��U8 ~Nqn.b�PQLB�f�0�P־���,�@�ׄ)���
bWA��$"А� �`�b����Ȑ�FRh��Ą��x��E�fj�!�ǫbWWqQ�!�w�E�c"�<BDTI	h��4ʰ!�
bB�)��+��n#�r�l�W��pL1�D��0$"4�Q(dD ńk��$�HE#$�XB#`I��,Ǆ��w$�:�k�������V	�F4X�l
! ��@h56F�IL*d�iH���`B0tm�NH><�O
���٣�s�}<�4j�䄒�l�g��|8{��E���%ҙ�6���y������&���d�����b�l����J��W%��M]�&�=D\Z$��7ڸ��U�s�\��CUa7�`��y�H�%���/8������,���c�aB��i��*��G"CA�ˆr�&�L,tZ�x��T������Tȅ$w/��0�ш��Ď.�H$�R57tD�A���T�����0�d��d���!�,�)P���oL5�k����b$N��D�� �=�b� #`X�4_v?|}�9�Bgu4&��T�T j'���B\�.o���&���.�(�|_asX]XC�|y�������}!X @�0
s~��!C� BB.�g���a}$�\#}�7$vm��!��1�,#�j�LIϒ,Y��<<�$|��X�!�b�� ��1����� �6�Lc)L!��A���2C���_9B�jNq�Y��D�W��d!$�{�䛧�$��6aIRxyVȵ <$ �XI�v$��h���
�lB��i ��"�- ���+�"E�x$��!"/��|@�O��1<`oYϽu��p�0׈|z@��aW|�5��,� �R �!"$$����bcɻ��$��{��5`�����y���=�%:=�o��E�'��z�׉�����>%}�"D�q�U�Z�h�<����`q \�o��:�(�6� ��;H�P#V��M���.t��O$��S-vq<%pѾ����L;!����#Lt��L�6p���[8X��Қa5�����H�thܬ���K��G�*�*�p!Hx`���E�S�]$��$.�=���#
K�4\�����	���!LI�� �	L�b4`	�%V��/*/��j&��#n&�Ge7<4�D�<�xx�ތ)�
��b���y�y�rSD8�?��[��j� �x�hD�=#��$7p�%�^�H�krk���B���������HI�R[�e�l���<ʢB!5"�V��2g�]G<R#��:V���xb���X@��Ӧ?<g�E���(B�K�C5�q�1�;��$�I ��`�D`I#�t���,�f�X���x�}>'��i��BV%bT�R�FT�<ٳ:�5��Z�Fb��r-R��S.ux�=���y�.b1��o\��^���s�8�f04�b1�*�-�-�Z��Z��r<�a�,i�O�4����fߧ�wy�ԕb��K�U꘡Us@-e�@���A `��`�"]Q��6M�܁�#H&:�z����:6ry=ѹ�A�u��Q!#%Uj���*'7���ą\v쓏��S��#ne5
k���+a��<�׉)º0�F�2�e4�ᧁ�0�����5�HV�]Jk��<)���ׁ/(iC���˲m�L�O3�#x)�6�������M5���
*B�&��f���#����@a7�:X�Lt+	4i�Ë��HW��%!bBM.!��B�+�Jb l�P��1$Y"شX�b��RPb��Ebd!#�!" �$E�# 0M �����t@�MF�HC�1���X2��<Hr�%ĸ�"��^45�����;"xzx���k��#ONy��0�������$!V01��x�}��18��y����"�V��{=�V˘����,*8kg8{�e��ɔ�7�3	����$$`F�̤�ܥ�ns�������"*��5��!��7옺n��m��4y��4II
2��.0�����)�l+�ĕ%��c/5��=�S)@!��*V
ń��L1��C4���Si�3��>�"a b5
������C�rS�ZD��*m�L=�lVI!�5�%�B1�gnv#]�-�7��H��VO�<�h�'���`�b�bW�yս�D�Ģ1!�H�����;<�p*�	�dHϾֶ`ƌ�� bZ��0`X,qaH�a�C�~}��n,uHD�#4d}=Ѷy�^B1*�H0a�6�B0OS���C�	�T2IRH�<S�!(fd����5�x��M���>I�Xȅ����#t���}GLj8Da�,���vb�c���#�H�
�`h�D�a## &����HBR�6�$
�h�Ec
�md!I ���wE��V!�A��y�D��>�p���e1�4���(F�X0 BJl�Z�2�� �E��	 D��3D�N@b�P�&4L$R�E�,x��k�<����燳F��44h�7�������O<)���<HP�Ӂ��А1x�C�h@�&��7�4�|k�B�f�l8���i1�1с���
x0+���Ӂ��:B0֍�)�$#�.v�8���qѭ���X��9O<��y�-Y��C�l⫉#Unb����paM�x$��CZ��i�B�B��h�+��4n%����x8�=M� �p�F��LM$����Bc�ӊ�`1ف��v�Z�!3��0S�HL1F�� ��1�D��o�9�K|�ux9�o��Ï��Źf/*�#*D��<|<<5�~%xP��D�+�j��|����r3�Ii�|��Bxhp�l�g����O����r5 ��M��Jc)������$HS��D����N4�S3���x�$#����#£�Ȧx�Yp�Zk�#	F�\{�UA!vbH�Q|:>��[�1n�fU=�Eȑ�M���wwC���t:�C���t:t:��$J$C���t:�C���t:�CZ�w����p%o�������5WwT&�Aه��;΄1EP��wwf��o�
�rt��d2��I$�B@���/r��a�VVLBr��ԐKRH/][��e���搆���>�NEe�tS��#nO-��I�o�N�{�wu ��$|�D��m���=��s*ֻ|}�q�� չ49<���:��&	ؗ�����]T�� �;�Q��FB�C���)}��҄�۪�f.���H�c����"������}��<�#��9�ts��l������u�H���|�S<d%�`��M�|�|`�H���e���J��y!�;8� �*�bG�� '3$!˔~$�I&�	<�d�C���tHd0�����9�is�o"���͞����Il��Z��%.Y	�q�� 2I�RS�� �<^���V�$�͢����Ⱦ��i��mp%�2LC��$�C���t:�C���t:�C���t:�C���t:�C���t:�d��$�Q'��>��t:�C���ty��t:�C���t:�C���t:�G%�$�C���t:�Y$��� t:�C���t:�C���t:�I���t;��^��AB�y��"��0�`�:7w����V�-Ԓ	K��A�L�Q� C���t:�C���t:�{�����t;��l&�C��wP<HtJ�C���t;�C���� vKh�:�C���t:�C����t�*
ZH$�@���E��! t;un��A��u�D� � {�Z���-�C�M0�L*-�|���a$���	�IF�V� ���*�C�Y�yiG��n�CRN�{�=R���A�����m��&}��_z�����b6�I�����WK�$<�t�rC���C����Wns�bX6��j�S��l�}�� {�n枧�9!�g,�r��w1D�ZJ$w0�H���ƛ
����0�ԑ$�(p:�%�(�,@�a��ƇC���t:
���ty�$��.H���>��a4�B�-�-$�����a��t���ؔ:����F�&�� �	��a���(�r[D�������Ϳ�f��� �$� N꠽I �p;�-��w>�}�ό���2�� '���I�(��^i��x5@ 4�`���$��	$x:�C���h�y���"E�+�'6�;�����t��s��t���1]��8J���W�@uN`n]��I��D"ݵ�yiq@�A���t:�C���t:�I���t:�C�ѻ��C���t;uZ���t*-�I�wXl:/u��Ʉ������F^'[9P�C9Bѝζ�W�~�o.�)��V��������l���_�^���Rv\���3MG�I���D�ۛ�v��\�[�g|v؞O�I9{t��ͩ�P��b�����H�K���v�E{kP�o��u�Ig,z���.�&K����r�K���I1Z��A,������t:���C���_6�y�05�$g+��U�0ȗd���MUm���3܂��ןw
����H�I]��ʭ��:dP7��!$6�GH�m!ٻ��~�  $-�Aû���	$��t6���F�*�^�ܐ<`RdK9��Kɣ����X�8���'�
�΅G%�+w�z4��ѦEM^0I�����a�%Ƙ0�`�H�C���I �f��BZ��ow1i� ����\�C�C!�i,��P:<}"���O$���4Ŗ����2xi�פ��lz�ȮV:�=̚���|35E�������'���|��>)����/f��rx�����v?<Xy�L�=�	��}�q=��=�'Zad���0�i���A7W�6�[����wU�{͡��@��d�1��e$���}��)�:���!A&sK�'*,�{�pk���j�Al����w&!hwj�����*����hPT��5��A�8M�#E��7{�H\o�	&j���Qm�j��]Pmf�m� Er��Rp9�  Y�꫻��v=t;t�6�c��͘D%��d�Oeԡ�@�`s��SR��|�^�
D��SNw�̙��M��[}B� 6��$q��	���ZVu*�s9a��g���$ &�/����͎�m=��p�8��;{ug�;۠6GMu�4��$�9�d�Oe�h��n���;2OJ�w����8v� kGD'k�v�� �X`���}3[lJ	܂E�|��#��ãi�M��H {.m:���L���$T�K�# ����3!��J'�:6ಷ[SĭsK�&��#Z쵺yj�.�;6� �?�t�oF�a���#��;}��P��:Czy���nv�� p�Q�����]�#����!.j��g5h�n�cf)
%�P�I%U(�/}ڵ,��ًRy��5{��"S|l��gVw����xׯu����ns�i��X���	b�]��u�nD�ԗ-k�%���amw ��!���X�������G�e�<���*覎7��ͫ5���$��j觢\���U��wq�E�3�]o	..O=���kE����|T�Ħ&�t�K#�@S}RL��Ѹ��9C$�8d(���C�[��A�%=���v)�5�0�I�$Hd�x�����$��Y��^�#��{����~��%�a7;�B�I��yvF��N�]��x<rD�d���x>)y�WU�cww�&�3���>��h r���|��y�G�[{�q�T�{<��4+�q���t#1,��w�}�t�&ܹ���^{E��wRn�wI���R,��"���o���s���n1��)L�=�� @\�6]�i�G�{ٞ��4�Y�g�0��m����7M0�fqNz%���C�vO_s�T��x<��h�Ы��䐀�|*ݷ�i�{lU�=&�v yi�\°��0��F�>�d/���5�����<n��:	�ؖ�ݫE����vta�yd�_ ���Gt�!%L!�4�Õ@� ��:wt�������z=9�y�S4H�wx�^�)��rhA���OM�*�9�u�H��wӦ�x���]c�۷��D q�;�[�C{٣�׉���F��/"~@�������HB�0ٯNx�6mñ:�#�X����T�Оk������#ZN���8`c�{�&/v��B�!$�s;~}ܨ�Մ�:x`[4w%(k	V�U�<��ǝW�"8>c����[�q��s�sn��{�$���L�  N��9���rXV�O��	4Y4�ݘ�����L���C�nJs��{�j�s!w��DHSV�5��:#���]+����M�d�ـ����ڑ�3�@]��B�r�o��wr����ݜYU*���B9��Z��j[o-��eK���*�A���\3�����^�;�7�� ���y������X)�B1C-�7����K%wz�a"��S�z���ȴ^S�w�B����Y�����:&Ja��C�ȸ>m��J�j���A��$8�HX$�t��]��1n�g�On:�/wws(�e�r"J�U�$o
��r������	7�o{���B0�rA={!��F`��f�I)���̣M�ڦ&�/�cl��8H�[�V��v�A0��{Q�0�g�2_�*�;���Hi��$<����d2>n;��t:�C��yШ�:�C�����	ww4بP8�C��yZ�tk!pĐp8�C���tf  t:�C���� �;%�J�=J�a��c٪f�>3��d ���wD�$��~�P�k)�>?����{�1
���7k�7�?}��Ϡ=�IF��·C��l
�w-���KgMK�ާZHX$�u����^����RQ�m{C�ǀa���&�"郟:�M�	����0H$�2(Imէ��j̩��?�ST�=#-��MJ�|6�t:�d�R꭭�V�@�xI*3�@�t:/+]��r�A�w]V�%�C���t:�C���t:�I!{�y�ʴf`�h�S�	���t:�C��wP�M�+C��Sf�!2N�l(W��³`B�>cA�(qyWL|{�,��<'�9������s\�*���$�n	�j��� $���a��jl���B��I'(��&ww%C��� u�TZ �Jh�:�C�[
�E�k��2$����0 A�e]��Mzr�rv$��hA�]�Ԓ
L��};2^��|<5 P�~�,.�(&=m�t��;�2kh��rtZ��䣀>�IW�s,���Ԁ}kұE���/c�F�J��$�Uh7}�����A�$�����4+ǰww��3ո�Ly�Ry�~�ה�����
]��7:c ���k�٦��=�,�F��G`�e�Ll����Ʀ��[���az��fve��{\<��ك�ن��n���?���{��`��K�v/>$^�l��C��M	��A��h���:L�8�Bs�|NH1]D��hG�Py���I U���ΰPPjk���	�^+<���ޞ	zt�����6s~�Cfz1�Ks	�I�[g�y��ݰ��HU�{�q��x�sv�
�ݘ��--7��B�k�B�Xi�1��O�<�+q���g���mɎ�wI�G���,��c��9E�w���t�0JM��X��uyE���6�2���M,���7��L�?��|�y9I$V�;��w�@ uHJ�8z��[�9����I�^wA��que�J�l�d����ٺ>�S=�fs��E�ִE�ٯy����R�ްg&��ӻ�3��H4HM�ǝ$����h�a�Z�#�Ǩ�n���?vJ2]�%�83�he���q�Z=���\��x�^��(���ެe���
(sI�O А�Ke�l���d��I�ܗusRm� �$w�	����^j�rA��Ԯ��3x�"�8@���-�X*MGt�%�fd��f;�����-�a=��)� ���Տ�ybǙ�t�?=wb�a|���� IZI�M���V��" �7az�������b�vn	>UK;}��6
�B�Rg��s���M�͆y������myl;2d���	�͉��Ǳ�̻On��nȗ�c�V!ݚ;������}w�|d�BzwF(��`Jj�6�S�`չ嘑�>�Y���$�$�n����0|/�V�҇j��n..�ĒA���f�y�H{���w@��u=�I'���P?�Z�p��$ԁb�ABjHVV%r�q.m�@�$w�
�r�D�Q7�E�;���JTX�iSv�oZo�s�I��� ���{�����Ȃ�u��4�r�ː\�hx�P�XI"�'v�&��ux@�u������YI�dӗ���Yslè i�;΅E��7 ���ȵ�v=�M�MJAӪ�Ы7��ʓ'�t�ۖ�����G�W:��L#X�6GI+o�]@S��a�X%Iy�����p�Y��s�G�쒻����u3$��&�;�,19r̙,3��wkЪT|���>~�5��o3E�M�:o���q�Y{H����;��GR=�I�TbVĺ��	��oWKH�  �a��S�����5�u�C�|d�uR@�� -�O��y�m�5��B@����C�r	$
����a��a��u$���2�S�Ҥ��Z����I����{Y?���Kw������1�py�KR\(|R�F"����䐁�"����V��A�!fY����7�֛8���'BZ.t�L$��[4� �t�����w��+��"u&�����7�
���D���$�w���+�� [5C鷮�y�v��
X���jT?;!l�@\PY�w2: ��P��$�pəzw�tn� {�n�rK�j]y�hR���U�y��%6�݂E�֘	pu�b)��I ��H/@9$�ݭ���9�����k  ���N�Ѧa���t���-��e�������`Q�����#�ڶfN4vy��BG}c�Q�r�	��iwyt)pCL��y��#�>�O�%�P��.[j�� �� t�� G�Ho���MY�ڹz�A��W�U(6�I���+J��p�Ӷ�m�@�t:�C�-X���T:/+o 'k�'{����s �(t1�I�G��;�otS;�,��V#��vo���f�8�KݺhsY|OJ;��`G(����`آRѦ���;�n������B����t;�L��A�oRJ��,[s$�@�I����@�Uz�.��=ݣ�H2��XD2����s� T:�Ē
��਴:�� ��j�d��0P�8Lp:)ցǸ�0>u+��Yh�:�[m�á��t:]B���Vl4�@ѱ5RI\��E"���ȒL�Q�:b�3^�𗻩�:�:�C���t: 
��I � 9]��v�����q"z�䓛q#��Q&�$���5$�$����y��!0%������� ���}�;Y,I�Hl��f�D����G.e�H�C���$H�i�C�@���@���A��P(t:9!!@�2n�G�]�*���D�ʬ�&ٻ+� .�6n�H!t^QNP(�C�:����iڊ�B�T�ڻd���T��6�(��(ONo�|�O��w�{߽��T�@*���ȭh��;�@R��|��=T��	E}?"z���1'�!�4��@�Q�)�	�U>���0U= ҩ����"��*,�"IQ>_$���BB! @��`�iT�A(���Ȭ`��H�`�4���M�R��  	�ҡ� �z��U(	��iA�'ȁ���P���A^ ��>�����@O��CJ��V ��#HH1�HI"l�|�	BD���@`B�	F�����o�B!B1�d, �d�0����H �����H�"@	 � ! �>��1#"�� 0D���!HB��TP҉�A�$@a
�/��X�� Sp�!����T4��E_QG �'�� MD�@��(���D}W^(C�TL��(�EB)�(�`��$P>+���m��@���4���؅@�1QQ  AB�_�
 *��EEP��z��"� `	;����cx�mv�`[9k:�쓨�3��@��j��	]#&��
��NkN�Ov��(�6�z��v�D@Q8�J�%��E��E,/'n�`�dHk$�t ⱋY�[է��ۮ3�P�}��;���s��:��ִfn��@��Yz)���z���-����]X[�Q���xՕ�-x�M�csۤ�@��W%����Ǧ���v�i7��n)��^{J�21�`��b��p��{5˸�azB�dT�;��;e�#�-OA�z�5X��9S4e�ڶ���.�l�s��݀����9R8<n|Ev�*rZ6�̎6��;n�W�rNٞ��O]�T` ��:���jG.H�l��egsԇN������k5�rf�]jv�Q\ �z ����	�C�t��Ř�QVf%���w�v�\��R�W
ԅ8��F]�,Y7Wo%���S�/�qY0f�$-�Η8olm�;�3�mE���ȝn��bK�Qb�U�4��!Br�&y�����ِ�T�j�z���2G�I����n ��ҁ�us�=��(�yP����L+q%)#�5@��\5!���A�Pڠ�ۆ��{���)0VH��r��@��� �˺�ջ���n�I��-r8�(�N�2���12ƅ� �"�T�ԑ:1U2aƛ���{�g@�ۓ:��x���R5!��X��=lj2&:1�P"��tݸj@�t�P9�t�{����+NZSn�BH�.����\ؿ�K15ȇȋ���� �� �5���2�r�����>^;���:�fu@{�WX}��s��v���� v�ܝj�gu� �#���� ���5�	�����b�T�y������;���F�G�.�������bHϻ�s�A�N������~�;��K)WE?p�㞜8a�LO��sr�=嫬[���8�ywVw.�rYdM8\��5���R^�@wv.Gp��ĤV�D��$e��>�@�}���Iy�1)��%�'��ݡ���hs������e��Y4>ř�����a�{�:���u���wtDm�2�ŖEݡ��L�!�e��,�8\���j�6g����gp�uU̖�A���n�GcbY_Ȇ���� o�X2tQ�!]�. ��.�R1���P�3e��W��ϼq�MH��T�$S(��Ru�R݆��ѵDdd�vL�I*�%�#�X{�q@=嫬��٘��}߶��}���e�nX���k�A;W��7vq@�zuG���������ہ.7��n����;
�ob�Aew]��9˭�%^0VS�7/l��fq�ˎͤ{7MN.�uz��B-��w���HPQ�U
Go��]>1�Z�gu�|nኃs�4���G��n��ft@��b� ιͱ�p9ۼ�Tg{s��$+S+N��-�ӽ�E�j�"�M�}u[v�^7�i'f!;<nݩ�Ǳ�v�7m��N�G\9wRIsJ��>�฻V姊9��1�!I#%���r�n���W���޹CMָO"���V�'��jꃸơݭ��mQ�tuqdՓp�H�e�" ��P9��X=mB �]՞�c}"p�Fex��n���hԆ�l�!�ѨA�p\��Y�wT��������%�8�;�3�W]�9�����U]Q\�(&h������ƶ����"�$�Ko�bi#N'K5En�wY�5=��F5���:�nl�tv��뤵h�j�yu�֝���)�r4�hꗧEJ�f.����{.d��g-E��2�F��U
�&��q�@l�Tz� 2pެ����sen��d�)P}�u��Dɚ��=Q�*�pԑ��uW5*��vD⎁�y�Xn��}�ҁ���Y���y9mv��M�@��@l㖤;�j��(5�7WfFIb��F�V�ݳ:�C���fEn�gX͝q���ͳc� c`1(9�_�oN��z�����{�H���n֮�G*"�@+� �$2QO�(�o���(^���A�y~������L��T(�ѫ�'=�~��`z�Z��F%F%BFaUHP�4�A7g��z��tΨ�oJ{���i�;S�U7W3JïZ���@d�X�f[v�I}�}�s�'r�����KW{- n�*�[���^㻻��Z��{��H�RLV)jQ�(�K���C}��U����h�1Ӵv�cpjLiM���S�x;�"K���s��{;�u���l��-�7��38��WDX�N�{���=�;~~F�û���������Z@��.U�.F�S$�;[s#�G*I/�gw�~������nI%�;������b_r��ⲇ9yw��#�8�g��w[m�hػ|�Dx�DDU�{�&I����d�3_DF�s)nTݍ6���͹�����F��M�~B^�
�ϳqw)��}K�#�!.L�v$)�meg�k���YS�wf��ۣF�rbl��؃�����H��΍%��ÿ!f��<�I �U�&�<+i���\m��l���������}�޹���������V�d���5����j��y�˼�,U��{��oS͕!����㻻�ʼ�p�7�F�d�db�$��x|�[�hT�u��R�7��;����p�w'r�y���,�;o[�dm���Ϝm�;����`-����.�W]GF�p+u��1v��%{���	�� ,!��k�x�3�m���t-��%kv���_m�.u���&�a�g���6��)�8n:+���8���\�c�η�HI�v�b�/h@0�m���)h)����z��s�wG߹���.�Pn�R���n'RI}��g�$�ӷo��.�\.!m�c��Njcxۑ�!�$�]����������K��i�g$�1�}����`������{��߿�����I%����i-[*4/t�_|��\I)1L���
�$���$����I/�{���5�����i��@�H�u�Էwl���ݜ�U�Ij}�Ԓ_nm���pwysMz����7�1bII��ߟ8�~���h�o��󕿱,���}&���_�V��Nr�s���J���=����[5�S�#iX�v�z�ÏcDvj9R@L�T>�qY�L�w
̓����߃]�n&����4�dq�ζ�=��a�E��AIy�W@.r�B��պ��A*;8h:`]]b���ֺ�I��w<����G-��	qz�bZ�h���j(��RJ�����(�%�f�/�K^��4/t�_|���(T�on�n_������6�"�f��1=����żcg_�M�yv}���"dl��+nF�*HZ�o_�KS7�"K�ͼ}�IN�.�V� � 4$G�
��C5%��s�[�.��ffq����̺�m]��^���$�����!e�hj�W^{˫���T9#T�6Ea)Tb2��$�y6cưP��}݋RIs�{�KSúȳ}�s�l�������ӖZ]#��=���)ȑ��%�I�i%�����t�T�K���D�v3�mHӵ0�Z�$���<��\�%�f*�[Y����~�z���Iv���K����Bnc����"Cwf�����n%��:`�{wu��ﾩyf����&��T�s
�I}�ʐ��ݙiwS�y-�ܝ3���6[Ke�[�^sZ���.r6������ F�ҩ�·$��h�A7o,Rg��w��^O�"Kw6���.F�S$�R?�r<p �-�k�@;r]�����?_;R;���wwwT͕!���2����qYC����E�ms�m�=;v6<��p�S2���3:�F��G95�h�4�R�(썶��]�����KV�l�_^y��1&�4`�_�`�!#BB$a HD�`B$�Z���p�@�E �	pHjeb����B,XD�0t��Bo\k��%�ZFUfC-Vڮ(`
 Cʎ����C�txe�q�aX/�t�CEnB��R��[X��P�BkЄ��L��R�V�I�3&�7���F��+(@#(�*D�%X�e%�a+��� ���F2�B0	G3f�qZ� B@�{0ZCh�$@��*`$C�Z�aB�i!5���	'��Ek��e��ȝ���Y�Vë��6�pu-�x$�[�P�뇥�!9�t�.6!�J��D�s!i"[��I�E��%A(���$���n�+�t����͔]Ke"[��l�m��f���#D�ݎ)���vR�� $9v9�+i��/���Z��\@Xq��%�-�nLZ���mu��FS��=��V��mœ�;a��P�b�M�K)nM���=�ٞ)ǆ�6��s�_\t�3�yn�;�v��QB�����"��N,r]���H��<�8��nw�o���:N��ś&���p	CX^��t�J{y���8��n�VG��������-E��7�-�mm�<c�v5�n4p�I�Y��+�v� �A�a�.��8r��(s>$��(�h�'���@k�:�],��\c����QL�ca�Ϯ��}}���+�͝�<��*g7i���7�]l�{9���]uly0�]����m��ht�*Mr{ .Um�-<��v�[�*��tt�Ϝ������v�F���A��n�v�v NwM;qN�`���ڶ���ۧ����v�i+�^r��٥Ξv9�.�d7 ��mW�o�~�=�e-u]��a�;�^M�+�Y�ᵦ/�Y�f4��!���[��N��m���W�%�CY�IÒR��p�ѭI�32�=GB>�h�E��_�E0T� z�����i�@����� ���EP�R����<���o���f���W\�s��o)a7�o�{�����|��i�+HZ�˲���ӣc�)��V�"2�%�7��	}LY�5��>tZ�<#V�;r`���lB���a��$�����%�z��ר��E��m�&���n��kr�(�
����B�y�m���F�~�k��fe�G9Υ39�x�fgOz��/�V�d��J$��r����}QD�ޛ��KSú��k�����$����6N2�d��m�w톶��ʻ�r������nI%۝�}�H�5���.	WTu�v��Y'����m�w톶�|��W9G3����.t;�KK�в�;.��G���6�v{q�g�">h,�,�qd�]���p���Nd���g:[�I�{9�tv܃��̰v^���R�Z���y��4��ɸ	��c�S�lHv1P�9�u@��qh�xWZ��֤�]�����W(��E9�߿3F�;��t$�9f�#���6߮#��[}�\\�j��GS�RȀ�f{N���%�ͱ��0c�g�����|�Z��*I/zf�����qw�~�ݦ�n�丧A�ܜ
�Ye�-|#m���לm����mm��w��X�%��[O�l5��ߣ���/�@�^�w�;�gS�~���w�/ږ��<?~�$�snw�4����p�K�q8�RI{�;��$���(�K}�Ӝc}�w�k~���F��M��8�J7Y~I-{8tHK�-�����P;^��u��Sp�5=�)]{C�W�wX~Y���߈�߃͓v-���H�c�,Cm(�hI�f�~~��^����}ðn�f�����ĉ��.�'b��7'�kEm�#����c�c����=Y��+7j�C}{�����͸�852.zW �q9�sl�6���ݕQGQ�X����q�jb�W 啌`�EIGk�h}�^���l@d�t�:ۋA�l6QsQv��v7$�v�:����7��ʁݝ3�A�㺳�ލ��A�B�9&��ڄKؖ���׶����PrIjaF�w�Z�ݒ��l��uuA�������9�\q	�܉��{�>K0棜��#R:�����;��Q�q�r�Ë77���p��([���>��mHӻ&Z�Dƭ�@Q���@�DUU��h�� 2p֨����|P���jM�tV��G
���+c9��A��G�ǔ�K�e7+�bK�d��~�Z9j6It�:��:��'�!���D�o��ӧ���N����ݛ�D����1fb��S�������@7Z���p�yI��S�&�mT��K$���'�z�X(�6�8H�q�{D��h�JT�)�L�73U_s�߾�:��'�C� q9[�%��E(��A�8�b�嘤�Ű�|���� ��-���DGd=�� n=^�,���$���T�2�͍�/�r"�r�|�5�{����f&׫�����*����WF����ܓ�}��͇����1
R=F�	DQ�Qu�x��#�������'�^��s�N�]���6�m�C�ŉ~X�_?w�����Xf��}�s�G9���_#�ߑb��vȬ�Y�<�ա��7�<E��zv���������� ج@Q�����z��ߦ~�>^�t>��q�R	[!p��?�2�c�����ر(���恞��T��@<�g�#��; �<��^����7j{j�T���x�=��X�?+����o$��߶nI������/�q,�~�?��]nin�l��]�����@s�j���9ɓ=/Ш7_� ���䶛$�ͬ��C�Y��/����+�yxެ��vcy&	�!$g/j���UP ��5&�h:5NKb�m������= q��|Y^��O]4k��Z1XkW-�7k�S��1�+eE盩K3�B<�v����������<tk�v����Dv���먲�+ �M��W��,=�������X�o�J
�9&P>^�uA��o�-�b��i�� ����t�0���g����0��ߦ����Y��7�I�(ق0��шQ�۱�d�/�-z��b�}�ڴ�l@l�����~�A�{�]VZ����dܪu��}⡿�P�������u����ow��G1��Mۢj�@?S<���*���9_?|�����P��Ԏ�0MUrZ�"q�~�DNkQ�T:?*u��r'u���=��~Ɖv�
U�(��2l҅LqVB���$��ʄՊ6X�q�����߿?ް�g~z_��[y�>ҕ�n�s22������N��jH��b�<�Uc�v��������6��vB�.�7HE�vl�ׇ]D��/V��Fs#��mff/Rʝ�mE�5��lC �ىI�6[|�{���TkT͸���AȈ��������$%�j��6��{zoؗ�1b���lܓ�ߴ~ݓ�߯��	�B(�5�}��mwfʛ��I�~�����o�s��b������rN�����{��줊U��G �Wf��$��ؖd������ʃ3m�>��G#�G#��>�!w�?���یU�0��#v��yuA?����a Xڀ�IQE\mV펐��4�a�f,_��߻������:��t�����G2eh��Y`�+[
~K1/�+W{uaΣ�*�������s���#�7�����L���1̊G��(�ムs��o���� �����w��Oo_�Ý�����_�I��ߪ��l�I5��wj�_����֡�9Ȏ~��~����ߔ�?��s�\�C�wl�l�������rs�ʃ|����A�r"#�"+~���Vo#��M5�H�y#QV�y�	���lN�#�mi��! 壅��@0]q��b��w�=~���g;���"&Yn\CK*�Z��Rʘ#Q�K�b7o'h�����^>Ru�@uֹ����A�f#<�߾������]d�[v��UtM�>�}�o�G��� ֧����n�����d���ٿႄ��{?F�G#R�dAP~���P;�yQ�Cj�D������~��?�F{�w�$���t���~��}�DA�p� ��������@9��@C�*G=����������jK��v�y�W�~��@�ĳ�Wy����t�ݛqmpu<\[p���Rk3/�W���������?�� �������%H�I!����H�E
6��%��X"�:ѾNk5椝�s���7�����t�{�5Ȏ	�]��j�7$��{��(~@�0 o'���������s�j�����I�g�����Z�6�c�;(�ݟ�=�Ν��X��R}���=�>��=�,�Um�d�Qe�C�K�F`O{�����ߦ������� �B	B)��I4���*�	Ҳ�de�1I$=����v4i:���y*�0��B>�]^���{n]��ȵ��bkǷ\��UbW �	��d�';���zyX���d�s�%��3m�k�[�ix!�C�qY�D\샊\��Y@���K�f�����C�ߘ��I��an$�n���Ψ&R�|�m1������;]�ݴu�j��D��س䐃~��~<y��*�zuFw���q���	����B�.6�!_�$���1r"����!�}(� ;�l�"9�0d+�I?}���'{���Jf���h�l���}�7嘒��bBX��?^����{����'�{����E"����;�~3D�wn���.©�����MH<����P�s��ꐶ;�����f��b_�,F	 �"�������Oo����=��}7'Pʐb�?k��������5i\��7G��)�{緦��bX��rs�~O!�۱:ي\�0�����JCY�K3$�_��R)�~�������� ���v����ږINǓFR0d�Ą�f̩�hB�(�2���Mx!JV1!o([�V\�Ȱ�*Ѕ0!�hb�!bE�BB�d冕y �uaLSP�a�$�ӸP�z!��V2H#0� `B�V) Iõ�H��!�P��:��21��y�b'u�a�MH� HX0 ���,"�h�I%mY�m�..��R�p
kE�i%�\	9�y/�9�)�%�¤�yD��܌J�9�R�ԉǆ��|1���e	W�ad1�!�R�,%M&�`B0bā$ 2, Dd�d� F���NqB�z�^qߨ��C��Ѡ�1��aRV5H�R%	H�b2bB.���FHBI!	K��!p�IQ���J��L��ɨ}�~mm����|Ѹqᶻ�b���<�=̤5Z4T�t�J�Ō����g.�#�M�#F�tqn(���n����!��ڹZ+���I�m��v�V2�n1��/D����s��8`j�����#��P^ ��7l��n�F�re���Vt�Y�ژ�΋�3�Wct\�ט�m�xrv�燛����u�j'��n6��JY<g
WBmm��q��xCb������+vz:������_^�#�;{r�;]��tnn��z68'-�"#�7�bI	8���9⽭��^��d��uӂN���ph�x�2og/W6ګ�7/m��q�1ћG=�ޯ'F���#N8H`��a�2�]�O���m�T��*�bu6�!�!����A0y�PGh衤Q`���}
}ϲY��J�@n��͆��i�-�����$sj��i�F:��.x����m���nV�Ξݳ%�&i��ՓU��	g��y)m�B{>j�ƂQf��I���~�߿~ՠs�oD �[�s���b��� ���*n*��Җ��J�����$��Ŀ��S��_���_� �Df���,�B�1T*,���Ԇe1��G#�*�}�����Fn��nF�J6�#V���1z��H��@n�g�"'^o�zlnR*9M���y�X;qXЯ.'B�m@�s���Bs	��I�b��~�t��}�=�zuFx�H��mmpl�yA �D��k�lwe' �����;�z��v�n�⇍��R)%t[u�wC��zj�dX�BY�QD�l�a�"��P�CXH�`��).$�6S7���2�Z�җp# �#��f*ks���G@p@�lIR���#�m� 7jʀ��k�Tk��|��Z�VD��?����os������c{߿�(����Y��ܚjI,�A,mM��Dr"[k� ѿ+�7(=��/����C���8�L��n��V�O���ι;}yuӰH�V�WI�9]�\++a܏{ｼ�=:��n��s|�&YdX؏� lU�vI�`�31M���@=���;,֨75����}�s��Dsh�m;���\T�X�쉧v�{�����?!@�b�L���~�Vr���>ݜP�h.�)�H�n�W���_u�;�uiŹ�w1gX�
	��!T�($@(�  1 X� H' �DfS����*N���&�D�(��\�F��O�� ��Q��2	 @��CZ�����O�����O~�훓��~ �X#"#X���W߬{��mN�s^괶hs��@�Io�,B�-v���\g`ó5Vҽ5қ/'i4K�	�Ą����ݲ~����'�޹C=���n	��vb 0	�&#"!�k 5Ț�>\oV��@���s��v�v��T`?zK�.�B�ңV%�כ��g�D�����߮P7�N���3���ÆF�en��j���5�B�l�!�f�A��B|;'l�Z]�Zz��Jm?�_�,���}���|��Q�Q�"G-w�$�]��1��V��30�˺�'X0t[+����^����N3gc���3n���hNZ��j��sUyP;��I� �tu.l���L�s�v�Qt���ň�����ӬO���6mɢێ�)mn=p�w�s�yD�T������}�}�V�f�ݻ*.��h~�`~��WM�#�J��ht�}mٲ��J�A;�$�l&>��Dn���d=��8�7����lsQ����
���
+,Fc�nF7Xn�\�{zP=�]��3(w�Ƈ}k��)P���]��© fN��Ds�&y�B'_���]ffcY����5-��F����o�΁�M��wg�oJ�WGW)wf�ݖZ�O߱$����~4�O�= ̝j�s��N6� ����wq5Sj�$裃�|��1�D��I"i.;uo]s��k�q��b�=�~���z_�H�5�늚�-�떤���Ur��k�,E����.	�ͦ�ז�ɝ��od��Tc�^z�p��Uu�^-�u�<ѕέkmui��mz�S묇a�'6��H �����.��m�_��Pڠ��9�n��f��J�l{$N^��ޛ�b�����:�������C>����%D��e����j�wm���9�U���9q��Vok8J!��-Q9$����(�￮��׿��s�t}�:~F
g�������2F�«jq��>��ɮ(М{�[�P����D����`�H�۽>����wg<o.�&�RJ݆2�ǖ�EF���Q��?,�Y��v�,��A�mBv�ϣ�s�r#�_�ՙ��7�Ĥ+��Yj�>�v�9��;�DATd�ڠ�����/����߾g���Y-�,u�Mu٠}���@�֫�s��9�r�����@���E��CQe���p�(ݽ(�pԇgj�r>9����yǧ�)�,���u*����C�%�.��n�-ш�r�v.��i�������+��9����7}~ru�}�tl�mZ��cDP	��d��<�3�&#�1���r�����}��1%�w�}�^��}[��l����]�hq�����3�,JC��U�X���.�t;V�q�'k���F�9�����=�74�H��@��Ow~�@�|~��v�I1GSu���(=�G"q�R��e�H>�mG������;TUW2&��˷�맾1�z�tE�Q�ҫ�#8�\#��60B#o��ľ���Ǡ}>�P����]Aw7i+���5W��T�*�V�V�l�!����g#�HU�4����@��h��5!���g�xN��2��N�M�@�vg_��ߢ#��=������� v��9��G1[���O�-��f֞�v��@����}��(�N�ot�����2(�J�����'�r#���|�6~�Ԁ��I�6�B0�%����FrM��~S�p�ڍ<�N&�!�`I���7b�g�4g-�p��ʛ3��]�+X�|�+���7M��F�y3�Ǝ��d��ӶF��f��G���q9%{;pz�$�=��l��8{�d6���6wt�yiKU[cQ7�A_��T<�v���O=���)��]�a5�r�m���� �IlZ�������x�I�ZG�]�&�e�V����@�w�P���Y�"n��c��уts#��X��X�����P;���Xs��V�{����%�b��C����`��߇\�vǶ����y����bŉ,���~�l��{�rI�o�o�����~���u��T��Ŋ�������\�r�]P�}P}��(n����jT꣸)%��� gu�~�����_���/�o'���b����������F��nˣ�T�@>սXd�l�q&F	E$Jcy#2*��H�V��8��n�Q�x�����bgvZ�7FK.+�q�4��H+`@��#�os<���0
r"p۞�Lˆl���bL�7�-��A�W]d���A�nbr��fQ����ۅ��x�b��[���#tݶ�V��kwW�}��(�;E۰���B ܝj�g������������,N�H�Ɍm~������;G�}���|��}�رbK/�����T�7n��l�����m5!�ڄ�i�":��+��k�Y��Ct��fbS���@;����<��}�O���VE��������?/�C��+ue�
EX��#�F����l�چζ����x4�i5�ۼxyoV��u�����r�ݎ��2S��5W�e�f�� e?��	 ���34z��Z%����5 fN�Fd��+��wE%u]������bX�����e0�HIP�Tl���(�մ�?
���D�T.���=�䓽�����}���?(D`�k;�g�a���7�����M�r�<����sZ��DD���h����/=^��	
���#�Y[�f �E�  (A3>����'�ϾT�b�8߭8u��wuR�S;��M��;Wu�Tkv+j"�Gۗ<y�L[y+�9�����E�U"�"�E>�������R�� ���5qWH������d6�k�.��[D�e��{pԁ����r">�9�� %���:�~�������uջ7s\,�[�N{�����@�.d�����O{�?� �����	&%#��#�R7*øڄ��H\ ����9p� ����@� �&FHJ�J0�0�4D�����K K�r���f�|)�'�P҆*O��`��t��&����B���)Laf,�.�t@�d!!:֍jH�%N�@����1!$H0"�BVecYYR!B� �J|
uCFC�;��a����F�X�B��A'�֒S%���R�B&�"b��_���2��R-6��%��/����F�ٍ�|��/n��V{]% ��v���`�E$DDDQ�".͌�G4$��l��3�i؇�\a�k�ý>��Ș��q�;`���zX�pB�d�{n2I��e6�ne#j'vb�g����-�s�!t�J�3�5q�1�'�-�N]��^�h�p��cm�NKn�{��ۍ��
�\#b;U��n-''<�2�gs�;!�wGX���v�۬�lR�Ӏ���f��jIU`z�,\��u��=��E�u�'z�ܗVQ3iL�<�2c�s�XrhF��`�Qͬ�:=�on=��Ϯ��P��X686-Ѱ��y��fԆk���qہM��i�t�)ڻ.�����F�\F7kkC�ڶ[kc���Ѫ�Y�dy�ͰE� EV��*�+2E�3���N��`d8�r�e*��K�Sr��'[�5����v인�Y�!�;=��m֖�+sN�'n�50-jr%qg�
ۊ�C�ݟn6��
Y�]sn�Xy�82����4&Rl'��Y�#�۹{�k`�9���Hm�v,*9��]��\Nݦ��pZ�n_������%l�Ҽͳ��;N'�En9z��֑�A<2��m'9"�RK�sMi�Fh-)q��k��S��f%�bĺ��*P(	���DP�!P�Q=OT�mx�.�OB
:?��E� ;��g���w����/O:vT9���WX�?�f'�}���(@�v���r"�~��Ti�>����IkpuH���(+�Qg.)n]1�܄ic

9  	��yok{����:���K�E*�`�kDD�m�j�� ��Q}�37v��^P�{W����{hʆ�G"9r#��7�P��ꊯ���%v%r����}˺���8�y{y���_ٙ��f�%��H*�����sKs�!�f�A��H��wF��]r&��r�M�b~}��Z�gwd��ﵹ5�ԯ�4)Z4 P�H�!!A��R�
���}�!3R�}Lq�1�)b�0)�O��]�Z��ѵ�j�/d��d*��06��HCl����of�/p����H[��sϓ��·�4b�ӧ�8�֎�V,����Ԃ�z�z�d&������Dq�@tݴ�sj�c���Gi�y-+H�c�K-e����$�$�3*X��}~��{0]V��荄��h�{t
+�D蛊���
�H�����`
cCu~K3�{��P��T�y����pjF���\��9��2�Uј�*�̶�ʺ2@n}�s����3i�3ݼ���X��9�}�3����hէ�Ձ�߿J�ٝQ�ù�q�ԩ��2b����΁��:�ٟ���V���C��b$ȣ�T婨9��{�MH�������D�h�������+n�##����gT%i7��m�zAۃ�	��0�FchX��1����A�΁��:�9��٫�]���B	�+�J"��@��r_O,̚��� ���]�~C}�%�ū���Hֺ�'j�73��&ڵ��r���u�ۧ\j���m3�C���9��h	�|��s��6�R;nQ��x�~X�������������w�B ���9��h��h5����\MUʫH*�Ur 2p־��E�f�Z5�}�;﷦��g�)3����G)G�m�K�@{޸�H��PfSr��mBOz�]d�[v[�M�t�|�~XbJM���{��5��[TGu�;	��u�0V6�Pv�‿�W��&��S�4#%ȝN��6]f�"���Z0���ņ,3}�����;����<~�a��ޖUl�\�qŲ��(�J!��L0U�Y]W`s�� ��j@�t��G>�G ��De����}ߏ�*�+[���\v`u�w�V�d$��(A@�H� Eb�A� ��+V��*T�r"r3�~�� �k^��~����I/*����-��U��oa�O�ʃ2��_�"g}�(@���{â-�={(��Urm<_%����\9^���`}>>��6cv�;ܽGM��Ԫ�v]�l,,�Z���嘮����3�~`t�l��t��Wa�fH�C��Y	�g��}���}�;�����x.�����
��a	e�J۸l�%-�5�y���٧T.��3�����;���$Ģ�S"�	V���n�(���۳����,��n`��+[�#a�^~��1�P��G9�G'�����֍I���)-�c��	C�-{��A�N�X}�P7vqC�]�s�7�e�	*��6�=���&j�EJW%+�1u������z{t@s��2z":���A�Q�*�jf�*�]�k���A<y�Ry9���uWrLZ�hԇe�H��~�s����Vg���<�WRF�(��1����5 n�k���y�⪠�*o�*�&�r����(���kӪ�r�{��&*9RLe�:�TݸjCwZ����9���U0���)2�=��e�d;�dL��Y�����P�Lj̴�]px"�
�7n�e�%:���.�
���w.�yƺ�)���ą]���O�Q�q ����Gm�e����m�q��.\�p��ޭ�M�w�{��$�?W~�/{�KVǮۤ��`{�{t��)#0����b$:��q��x����o���7����B���]���ڕvO�-۝]�ms+z�k�n13b��-H9�t�s�j���H��`㉩Z�̘�Y@�<ެ>ݙ���(���E�ߘ�!��,UB�.���kF�;-�R9��F�r�1"e+J���C�lΨ;w�P;�7�����{���·!��$q�@�<�#�
�Q14L���j��>�9G��p�!%���f��mB��=��̗W*�|~y2�Y��f'm��3s�X�X�b/
��M��n+!r�Y�I��&xG�,�ySz.8�a�i�a�E����"�5�Y0b"���$����t�5���5!��Bf�,���T��l�b�>[��w�P;ϹP=�8����nIc��(�oV.���o:/w:���s�Q6�)��%������;���q����Y��M��}t>=_|Ymr�r������<���@ȵ6n�Q;(�-����9�O<���x����F�~:N�Ԁ�Z���\UDw�T<����ۋ����v��]�&�Ru�@u���7v���Gd?k�ʆw����ɔr������{��~Q��`A���X��DDdD.s�͈��tԠ3]�����M�|�L�Q�ޒ&��@��w�@�6Z�r#���U�����)#�XNI"��cj�$�w��|��T-���퟿*�9~������e�b�{�8�W�c�1ŏ#I&&�3��F�\�V��*�mc��o=����W�uFoo�#�:��Zi��E"��M�8��6��{zgꃷg��T������ 'eu:�$eA�}ʁ�l��36؀s��`���nһ.��Rn��{zh�{٢��ǋV,�fb�ȏ*��R�3%���&�*�+J׍H�庺��v��9{y�>�Lꏼg<o��B[e��B�@���C=Gҷ+&�MvN�n�*�n�YP�D�9�{4{��@��f}��c���Y�Ȇ��m���x�<dDU�c8� ;9����jN��
�.�$���n)X}�P;�8�r�Xq��f���}����ViwSp����=,��[� 7v؀s��Dnk.�VǶK�Qڦ�埖,�߾�����۲r��ٹ>V0X��Nne�-�PgfwGe[���-��\����4�WM����Vy�N��d����B:W: �JqV
g��a���X�6��R�lL�1�U�ݍ�&a��lStz|��D9�3�:�>!3����lv^l�/K��M���՘�K�^��]��rJ;k����V�oJ<��4��	�X�;6�g.�m�/d8��s��"#�ߏ 3}�a��b�������O��7lsۥ�*��oXd�	Pr�Xo��|�WT�_T}�]�p��jR�Q�>��/�9��9G��|���Zsm�#c!˻ĉ��ĩ-���v�ꃗ�j�r��fq����ԩ�ݐM�>�z��C'�� ;�l@9�Z�2Y.�Ye{&�kr��|���>K[���c8��6��s݄�ܰ�0�RE#xb�q�i����}ʁݳ��s�~�,��%ݸ�x�A�����TEH��XVXVYIm�+4]��4�t�DcT"�bU"%B*�P(�P�'0��[OE=x��E����w�.N9p�� 0��Sb����Փ��峭U�,t�O8"���;��t[l.��^��񝳞m��W<�n��ORAr����q�ζ��la�l���qu��m�ˎ�;���`��p��b��W��Wav�F�\⸫n��$��69c����^݀9!j;k]���h�*i��B�w=��M��F��Y��������Td1��s��g!�3�[:���N���܋�n��8wP9vwpX��h�H�cu4Z�Z��N��9:�:Ô��o\���c�Nv/c�7'��+F�b\v�n�nPv������X���q��p��u�4�����i��իl�<��>���=�غb���5����E}�(���D>AvH!����]�TQ�"��t��"���̧Ʈ�t��t����%�`;5צ�F��30�l���!�N��r�Y�X��6�Ք�x�;�ʁ�6�mZ�n��G�+z�[�55�����c�P+AO��Xo=�@�n��5{WT/w:��H6�RK�6L��^5��T�l@kk�Ȏ)���V[�R�뱷��w�כՆ���a���COgq��+r&���2����=���ı=�����,��{>�ǐ5��>����9P,~��튩�\1r��odbԸbb�ľ{s���D�l���sM�Ը�d6�s!m�	��=����\�o����O ��b{߳�(r)��1}ڧ~x�%LLý:����*����Mq�G·�[�ȋP!(�C&]]fm9p,KϾ��"X�%��{��`r&D�,O3��v"dK��w�ӑ,K޽;��k-�����)��K�.����>'~ip8	�����a��$dF�"I!��P�Ue`�v=<qȖ&���6��`�%����yQ,�u����	3���ն�f��9')Ű�j\��,N����yQ,�tgݡ�:�bX�}�w�D�l����pJ��~���r�s�N�n(�UZ�r�X�'�����,��=��brD�l����9P,K���ቘ��{�ϓvY��'��ȹ�Z̛D�K���d�p9Q,K	�]��cz�qXy��C�rVV�Cr�����g�������V%��tgݡȚ�bX�{�>�D����~>EQ�W[6m'���D�uWf8c嶖�Z�LX��/�߻��D�l3�]v ���߻�9��,N罽��Dfu?W~����	n�6�͔���ı>���
��9 X�߮~�S�5��=�G��NA�����x�\3�Ͼ��Yj�W\���w���A�,���v������~��"X��T��tJ`���+�C��`i�
�O�Obj%���7�Ȗ%�bw>��brD���R}-��W\��)mc����$��)"~�߮�@�L�`X����C�5ı>���
�bX�'���͙�&bfuu�'�h�WSj�"恛A�����]�9ı,6Y#�Sw���e�kOl7��rP�J#3s���=�ቘ�����;ݧ"j%�`y���mA�,|�~�$E�WVl���<�<fr�����^�m��(�d�����7x�X��߯� dK��w��9��,N��uC�,��>�wc��L�~W�)��{�&�nخ�ై�,O3�����?)��,Oh�����`�����NA�,K�k>�`�b��PY}���qZ�c��ڧ,��Rl9Q,K��z�hr%�bX�g��m9ı,O3�;����%���~�\130��q��k��b��2��Mm9ılOs��v<�������v��ı<�s���,3,��~/ �ڤ�;h��Ej��n���[[pZ釞�h6ʹ�iW�
���.�Զ���%ڔwh:�θdK\yϳٹ��w%#�F�[,�:' =�q����f��y���^0[OD#��֎�^[���H�E=RT4�T�ڒ�,\�=�}����13>��jr�#���y�׫S�RుbX��Y�s�,×g3�7]vG\�Wu�J�;�80\�\��������j}Q,�~�fӐl��=ϻ�D�l<������%��b����fU|{���DqRJJ�q]ۮ:��Zbb�{��� �%����wT9ı,O�ٟv�"j%�b}���mD�,N�W��SeZ�b��r:XU&�ቘ�K�tg{C�CQ,K߾�7 r%�bX��]��r%�bX�ϧ����L�y�}�U����/"��5.	�,K��;�`r%�`X�}���yQ,��n@�ı;�}��LX��g[�u�5p�o	�o�v����"��}�ͧ �%��{�wX�`�'�ѝ�N@������qpXę�����{�����Z�M�"X�%�{�}��r%�b]ߟ���_���d��VZ9��Um�2;Q�y����/DX�%��v}ݧ ��by�����E�_{:}P�[��)7n�ʱz�#3�-abh��MG#�l[Z8hȗ���,b�]R��i�ѧ�UY�&�U$[��÷>����ge
��ڥ��EMY���+�������6K������K�iTJ��c��W�zb�&,b_���n�bX�'���͏ X�%���o]��'�r�b{�L���"j�����2[ksWR�NY"wqp��L��^��sr �ؖ%����k�9 X�%���w�Ȗ�by���ǐ2%�o��[e�s�[i6pWk�Ը,�L�by�g{��`�'~�gv<����,��t��H������$�>�B�1=�m�qi�bτ���}��P,K�߻�D�l߾�7"r�`~Y�?w}���2%����~���*����G�d���&bf&b�{��.������mg%�+N+L�m��[�6�q�z�m.Y6>y�ϻCȚ�bX��_v�9�L��]�v�4�b�&g����l����	^lk��A�4��8WCr8�SRೂL��]���ĸbb�����fǐ,K��=����@�&b���܉p�ŌG�]���l����%�V=Y�&bb�%�oO�Ԫ'��}T(��@�K��7C�,��﷮ڜ�bX6s��ۋ��$���~��v�WOvmU�ժk6�`�'�}�N��L�bX��n}����%��}�siȖ%�b���6�L��;ގ|���ዛI�95��6���%��w�ͧ"X�%��~�7 r%�`��_Mv �Ŀw���r%�a�=��4e���-����՜f&,b_OI��.(�11] �D-��V�V�M��a(�l$P�U[i�p���=�w��K��>����D�l﷽�\Q&gS�}�%v��wg䒷<	��xVF���i�F첒�İl���������<�g��r�X6���u�Ȗ�b{�ݼB\133�g�Wh��[��.s�-�ٗsi�ı/��wi�(5"X������Ȗ�b~Ϧ~�C�511c����qp��L�:.�'��iur'3�����͏ X�%�}��{C�uı=����r&��4�,�� �`��+KIVU6��0�*��:�IHFD�0��"��Đ�)�H�f��!��޻��"X���vgݡȚ�fz|�1�˫�'4�"�5.�abX���u�"X6����wc���/��k�9 X�D����x@��Ō_�}�T��WVp[	����@�K��3���:�bXsS����U!��낥���^v�+R�b�E��{;����ŌI�|��ݩ��`�a���r�X��S�)U��b��卦�E����1�ݮ�lUj\11cf/'�;ڜ�����v}ݧ"j%�b{�{�a�I�L�bX����~�ș�����ilz�b|���y$�R�LV%����6���F9"X�g�;��"j%�b~�F~�C�5ı>���eK�&,b����ݵ�WRk��8�@�K��������,O;��
�b�'���v<�����vg�4�,�L�~G�mNXX]\1l�Ū�)��K��;����N@Ȗ�|�s�NA�%������,Y�fa������l��$��B�R�{:��l�V�q�[[�ͺZ�:g���i��ש:�����zp��½�%����\YӠ�w�0��b[v�^���a]vKg�.�,���[������sƸⰘ�Ӆbc��Y
f����A���Y���P���&M�Bٹ�)ʷ��z����%��o�iȖ%�a��zʁ�L�&]\>�k<+��
H'�u7	��}s�]1S18�a{��r&�X�'��xm9ı��W�O��j�wI5Z����Wad�����I�,t��j\1i����gfw�9P,K�{��C�,����wa�yQ,���k� �0]��~���WNo-��A��r%�`X�Ͼ���~ j&A�?wGm9P,Kﻛ�(r%�`X��l�狂T��󳭯��ٹ�-�_8W5����l;��
�`�'��w���ı<���jr�X�'���6��`X��~��e��vr%�̒o��K�*,f&b~}��	p�L���6��bX�'s��P�K����j�|�ಉ3:�;�,�Kup�&��l*��PXę����]��11c?$�\Ӛ� O��Zp$rƄQ�"������i�]��w�"j%�by���mD�,K�߾���&bf}ߟ�M�75p�%s���� ��;1�qL<C=.0\�U��&b�IŎͮ1mv�=������k3�:�N�RCK�@v(�*��&%��,��,N�nW��AЈ�Q,��Ş	S`}���mA�,K��>�9��,K�{���D�l{��r �ο��[e�W[y��	�,z�N�bw�����@�L�`~��?m9 X�%����x�`�'��ϻU�*bf{��튩��	>]嶊�ͧ �%��}��9ı,O3�>�D�K����]�9ı,Os߾���&bf��Z�p�WVݕ�˻��r&�X���{�n@�Kı>����r%�`X��G{��D�lK�{����df}�>_F�X�������lU�\11cf.�W~՜�&w���p���6�L���A*�A6���s����ı>ϳ��"X6���g{S�T��>���ն�f�����������Ĥu�# ��ڵ�n/��b}�g����K��/���jr�X6��xm9��,N�w6�����־��������ܯ���.D�K��߷�����W�S�ND�K���m9ı,N��;����%��~�7 r*X�3߾�:k2]\1skc\�ld{��&,bL����v<�����o]�9��,Os��u�Ȗ�b_;~�ǐ5���Ӥ�;w8%�y�{wK`j\1&~�H�#�?k����r%�`X���;�� j%�`{��;���bX��s��"Qc~���E+�����[ye��.bX6���6<�`X�6oD�o79�7[���7L��nh՚�n3%��|��m9��,Osٟv�"j�b{�w����,}�;���m���	st\\uQ�U�Whܦ�i!�h�Z2�۴�Kı/�ϻ�D�,K���N���bX�����D�6�ߵ�nӑ,K3�l'��iw8%��Q�q:�.���b_}��x�bX�'��{�ND�,K���n@�K��<Ͼ��DIA&a��mI�n]\19��.h�r%�`X�w���D�lsٟv� �^�Jr�21�}�R+��.Yk�f��H@D� �0�ą��E��R1�1S
@`����
^s0��1$�D!A�d
$�b�N,��]�$5:�1��h����	B,HBX#�k ����P<�4�!<�Fx,�� �$a$JAbK�!b12}�9��,u�l�Uv�]�Nط34[[����75M��Gvm��l#u�)<��݀b"" ����$D��e;#Ev�;h��p�rŇ۷J�W9K��{CMFA��[\���W2�C����j۠�l��6 �WcrAt܈��NVy�Ԇ�:q�5���ٶ�ؕv'&x���$sʡ�]�r�tjq���/��a�u���a��n��FԐ��7�vc��p�@����m��B�p�F�]�6��+�4�\����0݀�ծ����L�,ù盷g1����i%;1m�����V݅��'Gaz[ݹ������h�9�˵��\`�8:���zwm�N���JFsY��nӶ��2Sآ��j=���6�V�kn(�A��ɉ(��!!�.���î�6�-f���N�R��p�:���;\pX97pn��f���[��۶�*�Wq�n-ح��vl�m]��0=���4]cr�YB��0�+yհ�Ԧ`�[#����s���r��V�9 �8�չ���i����ݞ��C�$p�Gb�$���7&�'���n�8pd�r���וی���n�Ak�:*���L�S��ڬp��(�*�`[c�z�[�()�j����*�t��Du;g�B[�f��d��Q:(�<��� ���<T">��U�U]�� O�
)�7����Kϳ~o�,�����ǐ2%��}���lr�pI�r.),�M��eq,N�����Ȗ�b}�w�ڜ��,���v���#�Aȝ�����8bb�/߿*~V��W\��4r�	%�r%�bX���]v"dK�7&M��߃ɵ�* q��f��b�����7<���7�&bf&'}��;C�2%�b{���hr&�X�{��������8:�+P���Y�Z*Ka%��.�����߾�ݏ dK��}�k�9 X�'~�}���ș��;�v~��D���ߜ�Kc.���8�nr�RೂN%��{��9�B9 X�w��lyİl�������,K��w��ቋ��_����-��l��ާ dK��=��Ӑuı/���x�c���>�w���"dK������\133���]�٫�)˼vܺ���Kı>���v�"dKľ�s��Ț�bX�g��m9İ:u�߻�8[�����t�a��֓�)sʉ8Ƹ�ڀ�a+8�;E�j;3κ0��v�u9y�p]��n����/=ԛf#ȯX9M�-v��>5�� p���tt�q/!��Se�śdl���5­O�X��%θdd�cr9���Aد,O������f^��>U��-�㯑鰫Rಉ31}>��Z\11cb7Q���9�Jv:]&����nÐ��X�R�ﺾ՟	C1/g��hr�X�%����,}��q1j��9D��j`��L"r��(��#qpJ���}��Ƨ �%�ߵ�w09��,O��z�����/���cȚ�c����rA�,���6��R౉31{����A�l���]�ș��;��siȖ%�by߳}�9ı���1�S���I��l�qpJ���ľv��ND����ٴ�K�a�r��z�hr%�bX�������Jbfz�;�d����M�p,*��������}s�����%��}3����%��~�@�K��=Ͼ�՜�&g����m���	I��|ݲ]fÐuı<����"X6��{����??A6�ާ�Y����Z�u8Ռ`	������ڳ�T���<�g��r�X�'�}��Ȗ�o{;f�Yu����o�诧�6&!��38�睑��ڈ�H[ ���&z�v���:Ydn�O���u�/M�]����@�l\�*���[��r��A�*�5*���&3�1!.������iB'mF#��$�k/S�%�`w��i�;�bX����eD�l�����ȁ n%13ӧ�ۋ�*bfw���b�@�W[˲I�K3qp��L��^��߄�b�%��{ۮ��L�bX�g~�m9ı,O�ٝ�D5�{��{�\�&�\1;I�#�eԸ,�&bf/z�7ᣑ,���o�c�%�`w������,O��7�C�,���l��z�b�Ѯr+b���T�ŌK����9P,K�{��C�,��>��9"X�����Ӑr��~CV�e��bۼ�{�af��1&b���|�pJ����U��G^
"�wa㑅.�%c,Hg�lv�Bm����;Q,K�N�iȖ%�b}���mD�,|��5sSWO��(�9�	��r��-˨\4k6���%���o�iȖ%�b_>�;������{3������ X�'{�?�P�K�}��s�Y%��6�������11c��n�@�?��� "S�07Q,O�]��P�K��;�v~��%LXľ��}��,�Lξ���n��!&��SRቋ�1w���i�%�`{���Ǒ7ı>���eA�,������MA���ܽȉiupŻ�r��.MK�.���{�{�iȖ%�b{��]�D�,K��n�D��bX�g~��r@����}ej[U��b��8�Q׸�b�&,b_OI��.������>98��KS!n:��n�8��`8��{v�,�����<�bX�'w�� X�%��tgݡȚ�c��ϲ�n��K��.Nr��5�)5��8��r7�(�t�שp�L��OΟ}w"X6��>�ǐ5��=��붿�)<��,K��?p�Ȗ���֩?&�%���Z�R�Z��\11c���]��~EY�D�D�?k����"X6������S�5��<��gw��/�%��j$�n]\1o97�ݙ��l9��,O�h�����`�{ݝ�rC�~uGH�F�dK�����r%�bX���>�C�5ǽ��kV��W\�9G�ВRቘ��"}����r%�bX�g߮�9"X�'�߮��2%�b}���r�"Qc�z}eDuի�)8s��.���D�l=>ާhr@�,9Mo95%M��*q���3V�Q�)j��H�rˬ�K��ɇ����Cؖ�bw��ǐ5��>���v� �;�Ǳ[up�6�\�ldQ��rBX��2���2]�㮎�/LXĜN��?~���`����m9��,O~�;"X6���g�jr�S<�_���s�[y��U�.�b�,O��ݻND�,K��g{C�5ı<��z��șı>����r	��1�P�߿~�sK$�j�Z��yr�aȚ�bX��]���2%�b_;3��"X6���;ݏ j%�D���~m.�0�z�r|�W[y&�w7�E6�`��hdO��t���D�ls���i�9ı>�_k�C�&,f�����#���ܰ��*�,t�uчd9m��s�0�%͸�5�m�[Oc<T��
�̵R������e��v��7$��1n�n�8Ύ�m�v8i�m��.ڳ�8�^̝�0`�����k��U�����\�\PܤZq��XJ:L��� ��f{;��9ڜ���0���k,6���f\��p�NA�%���gyC�lK�sW��n+�(�P"���-��T�Br�s1/�Ą���|gT�A�,~���iș��OΟ}wL���������\1l|���s�Ӈ��p���ev*>�,K��߷�ڜ�bX�'��}�NA�,K��ώ���D��{���b�&g}\?;	%SWO��\���jl9ı,N��ly ?�"dL�b{��z��r@�,N������,K���ݧ"Emﾽ�r\�i�J�I	Vi��y�Ͼk1 O<�}Cp�6�}���@�1.���ͥ�cfy���[lnj�M�9�d�+5.������w狀j%�`}�r@�,N���u�Ȗ�by���;S�2%�{٫�kYr�pJ���,�\Q&bf/���H�L��L\ǭ�A�Ƹ�`��N	q�����lv�%��}����&D�,K�gs]�șĦ.����\133Ͼ_lUH��e۾�ȢHBF"�T�Dk �R�$I,#cxbk2�F�e,��!J�R�p�t�v+�5��Ѝ��'FD�h��y��$:Ġ���)!u�v9���dV��ˣ�`���!��ё�QQG���%���,K��﷮��bX�'���siȖ�by�ϻ��D�l����K��$�;��Z�p�WNټ+��k6�`�'��l�ǐ2%�`w﷮��`X�'}�}���K��.�z_�\��+����_�d+����a9���Ӑr�bw�g�فȖ�by��]�9İl~�}�NA�,K���siȖ%��ݒ�ֵ��W[xM��B��Zbg�J���k�DȖ%��;�ٴ�Kı<��z��șı>��붇"X�>^Ͼ���嚸bs�88��qp�ŌI���};���`ٮ8em0��٨�fUuÉu'Rk����q�,��sΝ��/��I���߯oѥ��`X�{��6<�bX�>>���a����^56C]�v�;���URI`�YS5.�13�����p���'����� j%�`}����rf&b�vw�ቋ��ߜn�n��9]���Yw�����{���\��@�@����6��{v��bX�'�k�w(r%�bX�ϧٮ�pK�,�3�[n��w�$�ֶ���,K߻�~�9��,O{���C�,K��{��"X�%��{ߦ���13;����Բ�jዒ��kf]ٰ�ı;�L��9PlΟo�iȖ%�b}���mD�(��}�S�4�,�L�z)����iup�ͼ��q2�\11cf'�Nϵg����w�b�����,���JZ5KH6)e#�裣Q���=�ޗ�9 X�'��w�D�l߾��VpJ����8O�p��pJJk�"���"�\$���(E7 ��by����"X6��~޻jr�`���{��� ��b{�ٿ��LX����jT��b��ӊ��k2�9ı,N��>�D�K��=�siȖ%�b_>�f��2%�b}�5���SU2?�w�7Mh���W9�	��!wL��L�߾�~ipő,��g�hr���*D`�Ԅ@����Bi$?"TC��D�M�s����K��<���6g���wޣ�*#-[�|8ǭ�a�<�bX�z}��Ȗ�bw�o�c�%�`w�wi�:�bX�g��V�LX���}5��˫�)���yuu6��Ȗ�����Ӑr�a�,^qSȣx�
�C���[$#�������	�"8�%���F�`�'�}�N��L�bX��f|�ip�LL�>>�R5l.����L|TN�{{[;��W��ݛx�%7�"X�%�߻�~�9ı,K���D�K�����m9ı,N���՜f&g�|�L�[%�s�R��s!6��%�|�>��9ʬr@�/��s�ǐ2%�`~�]���r�by��r� �X6�d���h��o9_#�aY��%LXľ��_n��%��}�wX�`�'���v��İ/���i�;�c~~�Q�s�Oy��G��131}�s�(r%�bX��Fw�9Q,K���ۋ��$Ĥ�|�]��B�+L�2�p�SuQ��تSlp:V�қ��u���r�$m9uȲ��Wn�O-���]��lq���S�ӥ���Lyg@��=1m�K��ۮf.��]��n&vl�c\���c��]��])$�(�-MY�����$�\�e�K�(,b���k�A�,��˥w�%�l9"X6���ݧ"X�%���ݿ;���xЃq�-��b�H�D�E�%�����~��jΉ1,K��Ν��:�bX��>�EQc�v�|��=\1>sZG!G���0n���uK(�LKľ��{�ț�bX�{��wX���%�����C�,���;ݏ"T���b��;(ܫs�N�����G ��by��;"�`X�{��v<��,�u��`r@�,O~�׈K�&,b��ߤ���5p��_7u��fӐ7��=�g��r�X�'����C�,+��=Ϧ~�S�5����W鸸b�&g���[c�WWu�̐�jk)��K�K�h���"j%�b_=����MD�,O>�w�ӑ,K���k�9"X�ޝ�3&�\1l�-��tz��I�������ቋ����I�X�+��]E��N9��#�ld���gv>@�K��vgݡ�:�b3}�����1u|ϭu�U��.os�vFb�l�*J�������1��$"��$~ЅĠa�J��4��H$�n0����R����m�ܐ$�;�)�a0�B%X\R�f[%�"A b�RH��A2�$ FFd�����zx�@� �GH	"��DbE�V�H#RJmtE"B$R1XBX�Ida
�0$ �$#	Mm&��@�p�dcB+��@�6��KR@P�@��`@����B!	R`HE�D� �b�,�@� �
V,V��Q�8m�$�b���'9����R�x��%`�+p �*>�V�)�]/}�}.�.�v�)F"�n/m�Xñ�x��[PVQ�����F�.V���`4�r��D��PG�iy$��r�l��ļ��%S�:��j.�kiն����3�z�4˱;n�6����A]%pY�6���*��n-��zڲɺ�����E�$0gT���N��"K1n�mn;d9��6s��Cc�����SWES�.�nH��Gj��=�U=[zۉ�S�ہ]b-zv�l����ҍַGR����.�۱vvK��&Յ�޻	����^3C��>��[�����:���6b(]��㒝�9�u��m����p�rv���/	�����12�Z�3�e345�Vj*�SS3���`�z(� y��<AG���@�L7�d֞;9�!��e�$�.7\GV�;�э��]�{M���.E`fE�<�=ح�OH;9)��GFk�.���%�TQ��Ŋb���`W��$p�:G]W垉S1.����Ӑuı>���9��,N��;ک��`�ϯ��r�X�W�X�:W��.i��ʶ�-K�&,`X��_Mv' dK����`r&D�,O~�xm9ı,N�]^��O�x���߁�m��\1m�6Z�
j\q,K�w��"X�%��{3��Ț�ؖ'���N��uı>���.�����ߥdv�f������u�@�K��}s���@�,O>�gxP�K��<�g{��D�l=�>�\A&g����A���˶�l�փaȖ�bw=���� j%�I�bjqJ�Q���(�r!��m��[rBES{����D��`}���9��,O3��u��&bfu��8�VSWV��Y��U C��M;jE(��b�n�m�m<���%�߿o��r�bX�}�;���6�|��ݯ��MİX��~��\133�O��v���+y[��Uשp��L��^{z_��.,B|�D�8���&w���D�l��㹴�K��=�f}����g{>��\����%��uk5.�K��=�siȖ��>��7�}ߵ�@�}ʇ�ŭ>Q�	Z�*j�J��l@vs] ;��R}��G%��� ��1�ƘܢuLnP<�oV������P�y�u�1��D�Q��(;ۼx^�t��s��ޘ7��Ikf$4���ڒH�3 @��q��ܨ�mPwM� ;8� ׬�b�/���'biZ��(�s����a���=�.s�2�ju%	(/j�\�{��7:�T2 ���;۹$�_�l;���me�ͤ�]t�bĞV�Ԁ�P��5��������R����FK��G%a���(8�����v�닶煮Q��J!<K>��π�ڹ���=��7	������Q�Li(�a���jC@;�z����P>^�t��>�ԟ!�D�2��å�r9&�~��~/w:����h�9Ri�	����X@=�r�G9����~��߄5��cn:&�Pu��}ʁ۳:��﫳Af4����v��諊��mv���d�7]���{!h`x6=pS�t6.:ު�8͢��vM�'&�����m�ua�u=�CP/g�⌺X�m�<m�s�B��1]�΃D�acǖ�$�u��
��	�q�j�p-��m��ȥk%��X�����}�p밒U4ݰڥ��8�;݁�œ/��m4�JV��F���F�R�\s&4��=��8{���;^�Q�,]����8\c.�H�I�x��H&�̉�����㺰�ϹP7vgT{�y��%"��eR8��5n�o�q@�x�>^�N����F��\���9P;^�H��4�b��j��e��իJ�bP�:�?�w\�P���`j��@�l�}���A�e���5`l?=�2�ڛh-#�#�ʫ)mi��� �M�j���{ޯ��zu@ooJgth��+Yk���|�3��[t��G=���v8Z���p�`OТ�b�m͎ؕkj��2��n�f=j��u��E�I.�XH�
��T')sg1f,�ml�B�r�RW �*q[�;86�:�\�7v�2\�d7���#��`�VA�;�8�|�wV-ޓ@���V���c~����#��t�Bi5j�����m���j��M���o��7,q[�B�{˗X�] m����=�D6�75vMX��*�Htou�ǒ��LB.��*E\�u�k*` ������@Ǵԃ�b��.�B�����h.-��^�m�ıI�̊VϹP7vq@=���Y���2B��m�#FP=}�}���~Z�R1��O�OU��j{�*�� Z`��!M��"T8
k�U!CD�T�B���a��c��/E��P{w�kF��.��ے���	��C��\�r�_���Ŀ~y��a���C>������:���ri ٌmX=֡��j��Q�Tkޘ7��;7[��v�:�@[�W;�3� ������Y�m<!�4�!�	2���=�����a��F�W�չ���`ƬS"u�F`�#��F�C�}�4��Pl�6�6�L�%�\Iw�6R��- ��k=jkF��N�>�sq4����)2��ں���=�y�E�,B)U
���"	O�Q��k�rI�ެ���A���a(ՎIa�?�?�}��a k�yPwj5���3u�UڍH�n	$ՆV{_T&K$Y����=�Ѝ����c�(�B�o�/jꃹ�uf{sR|�IkwXӘ�&�F��m�aSf�s����"���j=�G#��_�h9�����+�SH���Pc�bq��9Ȋ��=r�����2�ԍcn:'J�(:���p��9ɜ��z�j=�F������J[f9!@=�ҁ�<�+;���Ğ���;[-CrRJ�e�rqB�k=Ha[���9s�*�IW�흧��s�ٵ�P��T����#K�CgY��ի�ñ�lx���hk{kwhSv�5Ұ��n��@���b�Um���2��ny.��Vk5�Li��d����}��Ϯ.�Ԉne%�Y�Z��r�l��V��kf8-�c���^�H���4�j51�����}�Ն�fuG����nJ�(<i��ҙ{"q)�
5c�W$��/���ӊ�����Y��g6��2�cUaWvJ'�ݖ�n�P�s�·�W(�)ĭ�
(偾ٝPvr[��Cj��#�Gw6T�¹jjƓ�v��+v�(^�t�]՚���"T�+�<������kfmb"u:�IQ@�U�˂v�F�lb��{��罫�Ï���ޮ���l�c�fF�M	#[��u	����9����1�Ou�Z�.��j=��n�`;s��v��ׄ�@D(��m���ٺ�H�q
�ıb�M��oldVF�*j$6݊�ϻ�� ��v��+v��r�{&$�rYfJME�� ��=r� =�h�_��K+��}'�M�v˰�[.]a���ր7hz� �mQ���]�P�L*��!h{�gT^�t��n�:�x�Ѣ0r�c�H'�T���@ٚ�B�Y,$����8�R*F�eR!��eT�*�w��X�ެ�t�ܻ�dmHY\���c��ɣ�gg[�:ޙ���ݦ�7+Y(��jC'��K����]�2���瞪�����5�RЌ`0%FQ(J����
AH�Dc(��B�0#��_U�<�K�g��}��T�������~���Ƙ���aq���z��� ݦ�ֲPk�17��;1�u� ���Xn��{ۓ:�;u�G�� �L���l�I�=�ڻ�>X�`���c����مm���,Fo>;pTw4���=jt͂]6U��>Ř���6�ȶ�%��3��� �����u�D�;������PϷy��RWnZ��HTv�u�P�pԁ�%��r9.5�J�&Idh������\��}m1r	>6�aL�i��\��E"�#�Q6��"i4) �6&�u\�M�Wa����=0b�LP�@�F�H�H��Œ$X�XE�!���imGF��<+	��ǔ �4�*�'�o��R4U�HP"VQ!X���F#	%qc"�禾�R,ѹ���K�[����.u�e+����>Ynfs'%�w<�8;4�ԑQDFh�#�E/e�l� �D0&h���b��8ڞ��q����m�횓�:3��9Ӌ�s�64M���a�f	����9@-���Ѕ����%�ɛ���=TW[�w:ȹ�����uT�6�FM>g�����-�W�`��Aj���c��(I�v�m��˸�n!@�U�힫�ƺq�Wkqq�vwn{8�˳u�	��@�<�ڮx|���m��y�R!lu�<�ɧ���9x��s�$���c{[����W�i�㳌
�����b�G���m��yM�@�{gl+a�@팹4���6���=�u��$�Q������!�q[�Ѷ����6X�k\��E�Kz⤌�a���gҐa������;;��=�:8�:-�[8�n��8źeq��[4PdN�;@`�9[v8�qS
&�֡�c���];�ƪ�v�{6ngP��+lJX`74�Zѹ�,�j��l��[6˲#�ZvWe��s�U��Z�7=�gYg��D=�a!��P��M<�g�Xv�ӽ�V�����n*�7m�{Da��d[9�YcgN���Se�V�{\ҥ[];�S*xy��+�m0��j��&�l�Bq�����QS�/���q�6����� 	��j������">��	��Y�Y�U��?oe�=�;Wu�{�\���	[��X�@����ܙ�n�ꃗo:���)-o��)����v�#�T��EJ≱
�jV�MX��K�y:�cjn�RF0�Au�*���P}عI�WXD$�n�Z�ED���T\��36-�8�H��(�tv*�)�A�=�`w�q@7ػ�|��7tc�6��+Vʻ��� ��jA�c� u�N�n�]��0ne%PyfDZ����}��íy��;��0Y����87P]FĽ*�ч�Ӗ*���.�v�kM ��[���֖lu��l�l���k�X�S�+[����dh�v��pd�����b��jq��5э��Qli+Jq��ڰ��WCoi�9wC� ��y`�����c�w�j�lrF�-�Uc�� �.�`n�&�FޕH��Z�L�G�!U����A���po>�;_�f�9�Rd�7O��y[��aXF�"*�Rʞ���ڠ;�ڠ�ض ��Ru��&��,�:�𢌖��/�?���_�V�~�X{��(g۽"cNe��1W]J�n�p�����j�����ލR%KJ���n���;z�����仫3�;�I�$��{��=��5TxڊkM��jEZ[�٭ �ö��ôlwݯ�y��Pv���XodĜ�ݗt�FbH�ha�����b�FcHȒ1X$d! $F$��BFR���a��$��A�` D���~��ߤs,����l�j�vٺ�v��W+��m9CW�3c/-J�jձF3G����*��ڪ�U��JHWB��1,��K7NT'������)B���Q�g�l�T�[v؀sZ��w�M�$�q��"T/%�Xrެ=��v�(f�r��'
䂩�@�`u�5!��� ��q�I�i��&�)]j�c�P;�;�v��嫺P���3��	�mHX��I��w��@��P��ET��[�{q���p��m���i�������T=��B8J���m�s9a�F��=�UW5s*øˆ�� �r9���wt�������NI-m"cE�r�}���0� ��1�������O}�[��s�u�ܓ��տ,ř~��.�lQI�X��]?J �ε^�DD�y�ǔ���3(Ԫ��q2ͮH=��Ėc�{��`{a��r[TͶ ��e�E���J��J4P9x�����^7�[����н^g;�����px�e�y��n��@>��Y�����+wv�ؓj()���Y-)j���C"r5!Pv���<��}��?���nw�Cs{�PO�L���,m�Ͷ/G#�&�߄�Oz״ע9�ww�܉D�R�ڛ�P~��P���G۴PEP��j�{���;�;�3۩�RW\i%��LV��#�2�=�@f���36؃܈��5Rs{���yD�w$I�̔����ԉ���i�j7l�:���a�`҃�߻�v�;����Wu�;��#N�\�m�Y\(G�����5� �v�t8�Ͻ(���2sI~��m{҃w���I*�.��T�������31(ϟ�|��N�X{^�Q�{��&&�*��⸹-ױpԃݶ Sr�7v��|���)�QcV8�a��r�}�k�'�{����ҐFH�HABX����\8�c����ڂ�k�Բ���XkY]�F��[=�J��%$)�i�h�lt���c�����a8c[����S�s���m�Ӝ��/lZ9�qP�I��u��!eRR[`��'Y��q�x<Ob�YP��
��9m|���b�߽�|������Ғj
��9����:����-}�<K�U�-�sV�Þ)1��� �m�v��}ݓ:���Ƈ:߽N�m��6)GU%J� �y<I�jdTw_T^�uA��r�}�8��n�#M9��F*�q�Pr�v:�M��۳��ޔ3�ٽ�H�%ˉ��A��8�{�yP�}Py{E�ۜ��$�ɻ�UrL��� 1��Rq��r3?�y�~t;���
G$�JX'���ޔ*N
7L�@�I����8Ga-m�� <�G��z��7vq@�>�CǻBbM�m�,@�����6��v�E��>�Yղu��M/�ӄn�Ivz��.�cDt�g68�ͳ��i���pܗ�倆�[�ٮ�w����xH���FE"�T�Ե���<~z>��=:����P=�3�3w�D��m��.��aXvs] 1� c�j��b؃s���D��+�6(�@�<�v��y{E���ꏍָO"jB��V$���fuA���V/o:�g7��B8L���L%��nN)��>V�ndзX"k��th�5�nG�c�%���|�z�7w�����$����h1�rF⌭�d�*���[�瓧T�]7(ݸ~�G9�v�ӧ�
��zʬ�˭��sm�7�{﷦��U������"+���##�ȉ�Ҟ+n-�ݲ���dX�?�J�#�6�h���d�%��#��L�yHg��Ptq��.&��K%J�T�wea���@��� ������7�J��Y�H�����m�k.6�r7.��*�Z�o*V(�l��!�����ޔ/p��s��A<�$���р�B�'�(��b�B���]k��jpn;��@k�X6�.9�$╫)�R�x���MJ����P=�;�3�v)2��IJ�G�<~t��9���.!,^�ǉ�C$"�Tu�~�n�IϽ�f�������(��"L�e���Xv�P�0�j�r#�/Z�J��q>�����G
��@�������v�S�p�⃵(���"���-��5�hԙ����"�_5�7)�㝧�i�?�H!�Lq��ݽr���vV/Ն����7�N!���T;�Csn��P�ͨmP��Q�i��ԃr[!]q�P>קTk�������o��r��o/ʳ��|�b��*�;��V�� ��T�p�Q�r��\YM��	f�F�uܪ����v��-�'O �<M���v�\��3-���"�Xv�G0�ѝX����ѓ�z6���v�6fvR�ŰOl���[a�cK��j��d��мDj�m������b�`�Tڌ� �T��,ř����-x�z9Tu����U��v���̩�G���4֜U9`:�e�KLchE����N�pkӪ�����Ei9���R�Y,Vܭ�� 
�ܣ����.UΚ������������H+�6�E,��k������a�q�(g�898�Q1Z�Wj���jC^�9��Pvp֨փ{"JE$�̈W#Y@>���w���P��ٙ��z~��i���bM˶�T��j�<��Z�j�X�2�F����g�u:�
��{!r`��������Z5!�Z��.jU)�&����	Iz��#B���):5r��M D �A�� , D#<_"�W�H�=G�#E)�솄&�D�vl��&,�.:HH�5*�Č֙B[sR�FB1��Ւf�D�0!4`�H��Fj��.�H<U�����`�� k�:HTH	J��LpH�"VP�`
��	�.������MGJ�0��ص��^3OK�[�S(�[@UJ�Bc �ˀSV�p mn�V���[@��3ŗMIc�wh���NZv:v�����q�sPA���m]*[Y��kQm�.yyi6�ݴlݗ�ۺ}0��&�r�1���[7c����yᔄ��]�+���N����6�S:^Knݫrnͼؘzy���s����R�x��B�su�v���;f�n�RL.Lm�����ص��m������-�ض�Ж�[m۔� �n�W;��c�mX�3�E���[o�s-pӷTx7�	{[\��;v�vplӡHRPz��B�3�r�ԅ�y��mp�q{%J�f�/�6������jcg*F�͕��4�e�����^Q|D� �(uT��⢛D<N���
�� S���V�OGU��7 -�TFٽ���h����^M�O3��&Dti_&�n�'����;���]!���N��5e���JLĳ�b�,şo<��n�V�F��c�Z���=>5��l@�v�ܭ�;�WH�49J半8P=��P�ެ=ۓ���·��\'�5!j�Uq'���r��w�@�xެ7vqCp�]I�L��+�y�zr�7��(�ܨڷ�>��o���L��Q��8���@`�ꑢV:����b�-�e���Q۳3=y�A��B��)��_.&�K����"L��r`�d�Y$sa�������zr�7��(s��U�TǦ��i$�z��Ŝ��1�[9��u��Ȉ�����9�nc����q�?.�àyq�Xn��}��C7ڹ�'��(�mI�藾�a��zPvu�=��#��p�;?w�D�I�Q�Ӫ1���|�6�Ϯ�#���=8��($$D�X��S������:��:���18��!1�@��mB+M�9H���T��ʠ�mB�k��%� ��,P���t�rq@�xެ>�ܨ��]߳bQ�Ͼ��h�dz�n]����M��zir���#1�b�
��JbE����E\���G9�%�b��M��MؗU7WE!Z����E����ޔ�rq@�xެ��c��nBW$i�%@�lά>�#�$�p���:E,R����VV�ML�')*��;����=�{vqC�4;m9��W�Lx6eq[]pn9,dJ��VE*��v{�PP�{Z5 <n�6�����6嶓q������{ʁ�ٝP��v�s��p��n9&G@��b �N�Aݭd�7P�βj�p,��ɑE2�;�ҁ�q8�r�����x�F��O�H+��-Kŉy�=$�NR8[!["ó�ɔ���xA.X0��u��g�a^y��Zԩ���]��TV�\ܜ�zn#]Cl�@�!ͦ.�l��C��km��u��F��\my:w=`�Kt�mLO>�Kg�2�u�l���Hɢ�������k=L G`����zm�2�����.���g9Y�·��O---m�br�]*el�l��Ӏw6؀;��Q����˚����#��s�~|;;l}�=�ڞ��"]]�]Ａ�Z5 <n��-�#�hrq�$�b���$�>�ܨ�Pyo;�=�aڃz$�RK�����@��Pu�d��/}�:g��{:E1��G��cʃ��\�9��@�Cj�sm�#\k.j�*�3M�i�Y���	^���	àtnL��^�W���G@��� �-�ʍb��:wRZ3}����b���$kuvOj�a%qss�t\��tsv���c��+6��N�	!��Lj�n����ET����z-�����n+{��ԠC�J��P/��kH5	��΀�3�@�tԃ�b��Ȉ쇧G���s_��6�,S*�	�`o�qf$�~�Xj�����w\��ڹL�pS,qd�dy+������P7^�P{�T{ݍ�$���\&52e��]Cj�sm�=�s��D�i/ʌ�b��19R��%nBb�ou�du.ɞ�B�v5M{�3��LXɉ���J��[�a��>��9�jY�u�6'���QY$��]�f<
�KI!�<�����@��]Po<��vs�y251�̉�Ґ@�u��9��""���jïZ��[ՙ��Ȏ<�Ʉ��Zz� 2pmW���Dɛ���~ ���A<�$���"�(�;�n����ެ=�՝���O�N�m�����}��>X���r印
������� ��#��j���݇�h;�l@d�AeӒ
���Yܝ�{�[N�8��pw`jaX}���W��y�ua��:�����xԙU�GdI����<�7zq@=�ҁ�y�Vn�>mG�ȵ9\z��{4��wZ��Ā���}�sf�_>�7'>�dx���ɑ����a��:�>��(���÷�8�9sJƱܨ��E�M��Y���u@@�x��ϷC�ʧkY�Z��i��ߏ�ս΀}˺���Q�&���7�rk�Eh�ղ�l@AM�G�~]ߝ���a��;�g�|����P����i�8W*�9$V^�7]�1�k^�nɬ��8�lyQ
�}˺�����-�t�ՙ��m9��0t�pR{��r"g4~�ڏyPu�P��Ȏq|�1o'�o�{��䵩\�*��rM�L���WR�6������v[y8)�u��;Zy۟6ٲug�g�����hT�<��rX����f�wZ���i��0��-7D�lW�9׮��j�c&� �GE�2�ĳ;�3>�J9;��/Ws_H:I��䑖ݳ��+��cl]���n�ls��vX�"ID�ｼ���({x������[m���f,�+v'��Y"�HʪB@Tㅕ���/�����k�e7(#�뺪���E�G 9���}Po>�P>�P<�oVg�s�Sܱ1�1�T��3�[��缨�3�3{7����Sb�;"�V��T�z� ������C���DB!�,��(�@����个�Gj*����$�u���C��Wꪫ�"|���t��3�[��4���yR(a����.�>RֻL@aȽ[�)�e�M�������r�#kCVn�+R�GLV�;]lV�^�퇊3�M �r��-�؉[����s1f&��~ƍquP
�pv��q�Xi���H�:�e7(�jtƹ̂pS,r��L�V�݊��l����@u�k܎Dre뢫�]�]��T()U\Ґ�w����wn�31oV}���0n*W��1��v����Ԇ:n%׶��d\�]D�3
X��`}�ҁ("4��P�:�:d�T60�������������C3m����F>:�st��k���c{��6��|x+INV�0=�>���נs�j�{�j3�W(��d�H��p�@���S�s��9�2pmPs�Pw6.�c]���O$�)\�8�
~}�P3v؀3"u�ʆ�[��/�7sJ��+���z&u���^=
C�Z�/ՙ�k�s�B��K�nN�z�ڬ����#%��&H��6�Q��n����wg3�w8G�eN���̎ݱ�)
��
��
;K��T�jn�R���ꮋ���T��qE@��XyoV{rq@���o4��ә+xҷ"��`n� nD�U�ȇ�9�]�Wr&��0Fᘰ��I[3{��8p	!��+�0��k�Ł! H�1 �a�������!8f �d���	�&2��)��"ĄB@��dO		@ FNF�D!�#�2���	#!��C���x��8}BJ��TIA�Aa	 �D(M�0�K���&��r�Fȶa��L	L�,H���p$X�-�BIp%��ع��r1�H�����D 	,,%X@�2�"�p𘱠�m7Ѕ`.ҩ
R	 ��b@����;���w6�"d�Ɍ��\n�ܶܭ�bK<�[\ac�[����]K��ɷ�����DDDF�E2D^%��h�q�y  �y�\̣��q�,C*9띵�p��E��ɀK�Eja��!+N.��C��YGo>z�9��v{k��,l��Ha��jEɇ48��pp\���vv�oKG7[��nC��،�8�w`��ٶ�Y࣊��6�-��O8��2�v0X{n����+����9x-�����X�;#��#������ӎ	�a1�:ww%spcsʸ�k����ح���2�����E�l���-�ڃ�.Mks���N��=�f���@�.��*[�q���Ɩ�x 
M�Ѽ�ܺ�\7n��
�
FQ�!&M4iBz�v��m�n.�SJ�v� �R�Uwf+uF�U��/�4=�R)фg���9�(��ێqۗ[7���8v��|�q�b��m��׍�����]]��JgW6z�Y1�;r��J�(�\���<��8�0��0и���w�+vy竐�۵;X��gb�.�F�O`닌��6�9n\��udֹ��usk90u�lq�����۵Y5���G�8P˒U��1N�śj�/b�#۪��
:�Vy�y*,��R"3�3�.���}��yW��GO��>E=
�E���&͈A~�Չ.s�_v����;���%�ڦ�����7����w����`}˺���Ițr�r6�
n�.۞l����]ӵ��ǋ����s����(�}�ް7�q@7ط�=���M(�]xd�\x�ZWTQ8��BU�X�����=� ���y��P|�y��F��!\�HEXr�=����gY���Ӝ��Nemƪ�p(�'Z�ܨmPw5�@��w#b�TR�v)ꐓ,�o:�Ӫ�]݇�grb��	 ^As�[�V�n���P�����Z%�oi�� �6�ў��
@��gKd�<f�j�=�H㣲�guо���u9)�m�m�.<��.��a*����T2A��u�OV�u�rDnr��%M��gUC�n��.XG-�Չn,I|�X��Io{���ޝnW]�i+7K+�h��{����ׂ�������=s�9)L�,�1��rd7hʆ��u�t\���%��r�!Ls�"vG\m��n�0π����o=;*�j�����oH�	�Zia�b�Xo�.�{�Br��A��I�YsWc�Jd�(Ҡ{�;�����g�eG�˔��$���b�T�\��֨76.�{�B3j]M(ڐ��%pO
�wfuA�-tj[����n��oK�m�&����.	}��H�Cj����<��Uծ��I(���"�cC����mxn�͞dT" �.|)e�6�7�g����dx�[M�K�[���t��nNb���F$���� ���������8����Y5wWE�?\z�e� �k�����������c�N7b�r��H�u�@fT6�ݦ�6r5��s�9�~����GJ����M;���@����<����ں���2,q�p`MU� ��fű �Z��Cj��s�s�m���;�5{7��iJ�¦�_�k�MN�uUd1�DL�hłO������8�{w�P��GF��d�ynHІ�#�j�d`
����5�}��Xnֹ@9���s��z�� �o�M�Qw��vYe��{��^�$��s,ļ�s����"8�5�ԇgc] Sr��i9�H�j�V5�{vq@���$z"#�ɜ�����1�t\w6*�"���>����g��T����o�,�"eR\�HL�;Ϲ�"�9��F�Ym��AƦH�$� ��1L�
}��|�ӊ���P��g5#N�@��<xG.#��y��J��������Pj��@�w'ݜP�sI�s%i�[�I�|�WT�pꃼ������|ی�b��5qD�v}�w$��}��4!��m毾��9n��oEr&ܪܘ��,(�l@<�r����R{�ȉn�R{O��#J8WV�A�>ݜP/�Ucqې~�^;o'%���m\�H�O �A���@��{��z�yS��(,�k#�A&�C$U�[�:���@�W���(�ܨgn��6�s)$X�M�P�n��׹�׽(n� 3v�߳3^z��Ąv�[�봲��y:�H�l@9�Z���[GY��j�R'G#��'(�ܨ/w:��wX�%��$��Iq>x�y,�	�촗��Ocv�,�j�Ì���ɂ:F�yfDt�k�r��m��g�F�$���1��.Wش���r	�Y�ħ�Q0��nw�;�Lr7Sʯ��kn��rV�7��]�tpX�)�m�z�7-r;�Un��$�ً1d���C�Fiݜ�����l.<2������}�rx9��z5W��\lbsW��G�|^�v���v�↝��nT��k"�$��ҁA�2�G]u4�=�5�l@<�mPvw] �q�������I�*����:�g��vVo��#20����iP;v؀0zՇwa�@=�bfԺ���i�ub�#i�bI�;ߦ��gQ���>:��n���\�A<�eR�VYez;z�T��NAJY���u�kq[�N���4��=�k�7l@=j�ݢ���]U�K���Jfa��S�D��$��z�Lv���L6�ў9�1u����ԛ�x:�'n���tx�q��9�R��o<F�d�X�kfZOW7��ϰ^�<�Ŏ��p�n=�V��{��eCj�����[Rta��Cy#������΁���ˎ�>^�t>��"�$�Kftn�Z��֨@=�bv��Fξ������,z,�O��G����?T-�t��3{��i�������e����a^"<h)��4��u�2������v87�U��û���Nް7w�(nv𠚵[�f�3r�b�r�J(�C$I�םՇ�M��u�r�w��Q�ܜ�Pl���ecQ���7U ��Dj*ls/�ߍ�-;���3�ϡ�(Yb��W�+ݶR�oZ��Cj����Dno�uU��n�ZV�KO�oO����>R[P�챸Tf8���u4�!m�ɴ;�ՠ}�sti�es,�unqѥJ9���]9N;g&�����ߵ���è7��P�y�����|����<V�ٜlJt�A���NGX|�oV���y���uuGv�nA�1Z�ʱ��<�vq˥A��j���-�1��2�I�l��\X:�{z���u~��� ��� �"�����`D�E�@�Wso$羚�n�_"1)��َH�庺��sP���J�DG'գ��\�f�*�'+�j����>�`USot�����Vy�Q��yC���ʢ����u��چ��7rR�w�u����G�>�$�á�Å��T�	f��g�e�!��C=����D��v:���Z�kTu�@����.����r.c4�_������I����|�ެ=��:��{��Ϗvr�dRIR�@��!�ڄ�������\�J'��j&8�1X��	BI���-*�+0"@��U0��h�2��p���5w��]��tld�NE�쎮Ca:]cS8֡�)��ّ�=k��l>ėx{�]\�y�Q �A�n�=��u�!ˮEc�V����0�j�;E�pn=�����=-�M�S��&����dv�=x�u�b��m�u�����}��]�8��{�PI�(��&�V��6�R�R+�8��R(��ʛ�v��`}���缨/ՙ��΍�
��� ��Hp{�ͻhDId���t���ڠ�mB �nm6K��¥�oa۳��?�o�ҁ˹~u��������q���y�-�����P��=���;8� :��p���U��G7Ur�,X�o������ݶ �s�Ȉ�������AH�%�ŉ�V
���\�,����\Z^6�i�GNF� pxG@6��k��x׾���W�g'�zai�Z�~ U�( ���T U� Uh���
�
��� *�� U�E��ET�aP�Q�*1DX����DX�P�T�0U�DYE�DYP�DYE�E�DX!P��E�Q(�`�DXEdUQ AaE�DDXAaE�B$Q DX�@��DX�T"+E�AP��b�BA`�B$D�Ƞ�������� *�� \ U| _�T U�PU�a@W�� _�T U� ��� ���b��L����3�Խ� � ���fO� ��  �  =           �  �
 �                 :�            P(P     �  =%	Q-co�w�uA�(׺J��ZLm�8r���tm��;���.��� �
IQE*���v�6��P3ݪ]�c��z}�i�[��}�y흏
��uUm�Ժ�in�^�f�����{���G����ټ�  x�"JY���G��W��:�t49m�S��{�ًy{���n��Oy���y��Җ�ާzS7{O���� ;�"������<��sU��(�V����w'�+��a����v��n�[�@wnrΕ���OO@���:T타tA#1�z�]<����77�;T2��V���eMx{��3����7i�����x��%P*J��3�{ں3�vݠ%���U��{�8iAtw]z�^=�s�eӡʛ�{ڽ�W[�x  pQ�f5p'^��=( M ��l� �m h ٠ d� �%�S@��`�h��4 3J�TQ
���m��JZ�@ � �� 2hl�RXҀJj` ^� � ���+-� 	 *���R�e ,�y�h=�Q�j@�i=�����2��{[�VuON�md�6�{�;� �!EUA%���PLUm�p.�K�9w2�Vj���er�u�V쬺<�榜��^�P�{����d�J6�  U?*�  ��T�)H�hFF@��JH�Ԫ�����L������� 	4������ 1?��@$?������~����L����cϿ̐�$�}ٽ��I	I&�H�$$	$���	I'�I	I#��C����B�L�R���/�?���R&���%�B��#�Ġ���*��B�㩫s[0�o��O�g�5!�|<����F!��6dK�`%�	p2��؜Lѳ���R2��P`h���d�k|����ypњֳ��)�%��G���^	NY��=K�C� �by��F�ۆ�w�	sف��Xo�Y��H7;xhMxa�a���|���(3Ɇ��g!��ל��(.�n�"�͙�}�<���[��Ĉ�hA���Y`�	���&���D���C�3�rd�y�CF�Ç��H%0�[�g�ݗ\㳟�ɽ�����4�2������k����&�<��o.���@���~ �d�mO<ב,�f� �ڼ+�����HK��y��S�����|��7���Syuw��{�.�%8��p՚�q�j�r��f�A���̹ગ ���0vy��e��7��)0�;��҃"�O�E��Sђ��+ ��Hȁ1`1��X1#�H"0$ D�
H$%IH$�$D	�	�Id��Ob��M��,�ı%R���B�ɢ9<��к�n����'��0=���іL494�h3S`���z۸p�F��q~�o�� ʌ���HV��� 1Y�4��E��%��F�*1� �����Ԍ�`��i��r��f���`�ρ�TJX��Y��,A���M�I8c�XV@����"B�$J�Q��h|=�y�`�QX�+$�qo4�b�z�����\fCY5�k�}2��X2c,-6)B�����A���ɣg�hLQ�����5�z}��4_<sC��	�>�\�Жd��5��I�v���i����|���b0LS�ob�,3Z5�Q�:p�'�$�!P�$�D
A�����=��FE��a�d*B�=�	f%2jS�2�����eo8n���c�����K�ŅL\T��0SV�f�w�9u6xY����j���m\���$A �KL�e��$�BT����}�|$.�,ȅ��RD"�$�.y�fFp�ma�8k��d��T(�0�ʢ�� 	$A����A�+O=۽�n�7�~㬶���6{Ne0i����䙛3D���G���6g&�%R!�h�!�<9�8��(ʹ�|�0� ���FC�4�0ގ���̚�S!�2ja���Jy"D<��rkt�燓K"$�%��F�O<<�Fȗ �]oF�g���D�ke�&G2�w*��{���sG)�3��y�M�ް�Ԋp58G{.���ל�}!&��%�W��9�<=43QX��A(mA%����*Ou�d�{OL��I�#!��i�Q�����y�c��$A< ���%��84ɠY��\@�9w�0�OM�37�7�z9��s<��Z$
R$d�U�_0{ ����'$J`��e�ǚ�Y�g�>�Á�2�ѣ|)���{�<<��K���<�o\|�8�e�j�O<b�8lD8�漉C�Md�b%��%4	D���)�zDģf�M�Y�2�Yc.��!�]�(�iP����0@R$��\��e&�[�l���� [����$�OA�,��g=ӯ0�[&�0˼��&�=��z|z��{���1ˁ��dL�J�29��3P�Pg��z �6a�]�N��!�y璔	�$@بE�1��C�D���0�!H!v�A3"d�7<=�\ѣq& �!H�d�PÜ\o"�K��S��7��~�^�O�"�d�^xf��9����M�̓.��[A�)�5!7=�Iw�g�b��ц���tF�d�oF�<����"��dQY|�����<|�npB��� �#H���\�JyNMϾ�"�� �4� �� dg�������)��83~���<0
�מ��>"�r�X�[�'!��F�&��X$�J��n7�'�^�r	ug�Ot�!��.4��,�M�8lnD���f�Qk���B�r0��Jf@�� r`��fH�����F(�5	���8SC6l�g��,@�A&&�����2�������yG �)�IA�nNxxr�7Y���3ªa��#��Fd���8\����Ta��S	��	�$e�`fjlC���f}%����<<}��E�4�h��jr>x�N�[�ɦ�.O��K��Nˆ�	���hQ�#A��C�rys��cr`��u���Ȟ/�Ё����x��}�J�A��0��y��/���`��D�##\�sxz�E�=A҂1�Td+Ȍ��e��F�,����
H�!��̚������F���a���2�F���2R`���"��L#�1�b�!����(`�)D�#�����~7��P�M%�I��y��$d�)`�$PA�"A"��I=H�R�H�>dg����<�6�LѠ,��A�Jr*f��	d(F����9�(�XX"D�eT�FX2ɣdBɓPeϤ<��XiR4Jo�hX\sw,�\2%4D��2iQ�)FX{s���V{1�
�F��Q�M_S]HjD����M�Y�6"(��z��"z>��F���ė"P1��7�?��7ǽ'�cK�03�pj�>���<�[���ˤ��<3p�X�#L��d�(���I|���Q+1Qa���L��Q%�����J����CX��y��zkg�4�x��Q��a|v��y��<$��j�����%Q-Jdp�+�e2*��a@)R�+��F���e�0L� �d�F�V4Y���%ES�n k��a�>�O��5G���`�`��{r�ߛ�xzxOA��A����D��3A�~5\4q�^��\�r����ɱz'Ѩ0DCJ�p"B�h�rx0a�ѳ�<��ȅ0�7���g�ϵ�*SZs�O|>X0C��f���!���b`� ����3s�OOO�	f�p�>�c�G����fÄ<2w9<B�Ds4\0����{����X!̂Y��h%e����sm��j&<��ٳ[�'	�LL�x|mF��Pi�76�'=<�d0�=eac,��W78�l��\ ���	�A�h�A��F��	�78x&�����)�7Y�p��2$vl�8rc=��3`�43W8���'�wi'{�:�������\F��-��I��y9)+.���5�،e��s����8���+#|���}��'���\7�~��"3��'�o��x�a�g��a�񡱚4n擇��ri�8Xf���<�f���a�Ja�N)�����x@�A�VA���B�T�
���	H��adb�R��d0*�A�@՚���y�{ҊIq�:2{Fć��"��������� �R� Otf�� n�����5O�`'�,�2q���)�"D�D&��B�$�<S4M��ٞᴸ]�6}�X�0�f�%�k�FPe��8`
��g�
�i��&É�!�ͫ;ў��kd��)#,F(1D1,fL��m���(����0�6k�	��h����2=�
p.A1�������h�<s=�U��$`$�i55��i�������)�R�''��ѹ�yS'�&���j7!c78�y7%�"{�o���u�b^N���rDD��i*�Lǣ �^}4ح�eg;��+��-�#�R�;�� ��lè��5I̲�ծ�`�Z7	��};�e�}ۛ�Wo]ȉ�\��(^��6j]�ʣ�aywp���79k�j��$���UW���5M��{2qi�.YL��+EbGhډ���d�{�Y��Ŭ����p��6���^�?Ͷ�^�%h���Q���ʜ#}���͡�[���dEp�`|�{���(��641#���HT8|N��{��o �	$O���]�:U�q5�P��%�\e��ל��� p:whxL�jk^I��n�D���NO��[�B�֗mBB�tjQI[�
#��B�/j%�IE��b፽q+� �lM�&g����V� Y<U�nr�Ts��~�j�I)] ����N��<��F�ţ!2��fjԒ����9.@x 9�p \�pd�M�d���[A�@`  t:�C���t5�$(�#���h�@� a$� jZ$�mC��y��I-�@�t:�C���t:�C���t:�C���t:�C���t:�C���t:��$��$�C���t:�C���t:�C���t:�C���t:�C���t:�C�[D��-�@�t:�C���t:�C���t:�C���t:�s$H$�C���t:�C�����C���C���t:�C���t:�C���t:��$��$�I!�v��F��:�C���t:�C��Qht:�C���t:�C���`t;����t:H4:�C���t%�$�C���t:�K��l:�C���`t:�C���t:a�� t:�C���t:�n�t: ;�$�l�~e�š�%�I�E�B_V�2(C���t:�C����C���t:�C���t:�C���t:�C���t:�C���t:	$�C�[D��-�@��t:��t:�C���t:�C���t:�C���t:�C���t:�mImC���t:�C���t:�C���t:�C���t:�C���t:�C����$�� t:�C����C���t:�C���t:�C���I$����t:�C���t:�C���t:�C���t;$�=7�]��p�!$�$H$� ��2{Z4*�t:|ޜ�E�I'Ly�Fc��I40S\�ݼ��:�=�-7h]�8NT('+]��"��x�*��9%˿E(�M�&I���S<C���,􍷋ӳ�{�-�0�g�(t-�i�L7�(Hw�U+{��s�W6�WO���L�Z�
��/n�K�ӎ��?T,8�Sju^���7 t:jo=�+��"�`(�n�<=���1�`�t��^�\,��e�q��e,>]� �Z�*)����gLO�G��<k����n�1U�,�< r�A!����,9�B@t�Qȯwp<,'M�OzH l^V�����wt���[W$R���N��_6�BD((P�$/*�$ԃ�Дl%-��+�Y<��������tǤFI�-�D�)�o*�����$^|D|�a��{��4L�&
a�jBt;�z�zR8{{���R�2�ڈ����a��IU�� yS��w�,���D*�:6�t��T8��O���T�]մ�wGT��:N����x]�$�5��o�H ���[��'Z�����|kv�\͜Et!����۳S�;R�컻�o����/(�<'8��5��.��b'� ����>9b���f�������[�tI��&�|ql̜l\2�IRI(:!ŃYs6қܽ��=��Z�l z{���C��Y�T��:f�0<�~м��-��9��DZ��g_ �����V�̜�g6�~7�hP��O;�n<݊{N��|HO�å;������ ��p�O�2����J�����`�C���z�����\\��q�8u㙩tOS��J��.�d��t:P(P��2NM�{��ߌ�u!,�J�!�?e�2v�0O\���J��u�Z K	4x�ʸ�ط�{ =%�&��aq�K�`�Q"��˧7�ى.�PV����&��ƒ�T�̾��I�x ����[���nDC�m�wڟa�ٚ��2��z�x#!%���s-��O�w6�m�N��i<�J��/|9��T�ޣ}_{�<�e�i���'�$�;��p�%{��Ko�'�[����;�����ݐ�a=�n6H�<��po
7$nw�s�(�@�t~��c;.���z�������M��"!�/L��.̘��F��ޓ���V$�� ç���s>�y�š������`ٕ�f.�E�tlO�NͪT|�[���t(jp���f`D�I$�<p�C⠞a���t� � �h����y$&�� ��� �v��Ha=�%�~�k�c���Y�Y��(W��$ e�ݸ��<�����ܯqŨ���sC���¡�u�ج���I�N�6��������C�}�$��eIޑ��RD2)|�����~\u&�&yrA�����  ��	k�kBa��n��}t�<�ni�``y��[d��"wI���ۃ�%�WAҹ�#�ZAQܐ���%�層[�m��* ������t'^��qFh��kV�C<�&���-����j�E����<M0�䔋�8d����7wv3��8z'qD�S�nqk3�	/<��cN����?�$XH�n�4��}&�M]�Q Y���� ���5��S�ȍ�WP�32oofb竅��b�C���:6����{S���鄽�"5�yS�a{�݁���zf�� E�5�Own���wt�faYRS��ƛH��]�6ؘ��@[��onx��w�Q$�0,bHk'%�*��x#ٶ�e�V�"�� �w�(æn��⼐���B�A$�΀ܭ�Q!�������=��\����{�;��2[�pz>������i{i�E��^��}T�zG>owuxݐ%�����}��͒��q<�67u������4@ ���P9� ̰Pgn�$�,���I�����X�a:��@yܵk�¤��I�9{�<�u����$�,U"�� CK�L}#cqY�;��Z�Ą�����CS��`�V��a��&�C��ߞ�8�%D��^K2(IW��aԖH�0>ҷ�{�q��wm%���s<������}	=�޽��?���J7.Q܀��� ����,F:n��u��)�;�ztAϮ#��}�v{9>�l�a��37w�ޖ��wJ5Z�P90�bԓ��b�7�.As��Bî�Q{�� � �l�:,�m �#b�j�A[$��s	y�BŠ@X��iN�]w m�\��t�f��9���(8yj��f��H%�JȞ�ql$�� wzFhx�v��M��ۼ�),CV;/]�Ez-d�����	�Ep��d.qn�.�w	ͩ�c�q)Zm���@#�o����|�TN]�T;/w�� �n�nX��F��3������n� w���V�"�zd>�	���Qώ�E��Ƞ���65�=ܜr���t۞�|J��g==kX1���[Gçӹ�e�6�򑴯F%�d�n�6On�٠�8	֋X��<��sU���Y���1�<�o[��?�K�n5�<�	k�RR��Hϖ��L���0i����^#��o����.X�Y�|� �A[�qw���O�!���߄'۾sd]���מ"�&�/�6��mK,�X�Q���Q�0vg��"ܠ�C2C^����� 3��5�p�^WñhBIWRH:$Č���r�ѽ��zuȱ��O:�a)b2�K��w��
��wr���:�x/8�i�ֱv��@
x8�Ͷ��ݒ 5�v�hP:	.��d���dp$  r\N��R�?szbI�6�y꺨Fd��P��Z=���Λ�$�7-�2snw�)�*�V�p���1���E���o>��݆�%�'�|/��!�LT��Ē�EN�rGf�zAzJ�m�7��D���ͦ���{-d�n�`��ļ�ح (9�� K~�8�w�ʔM�3}a�>�4R��3���{ԈC���wRy�3�` n��I��|��&�zoQ�];}}qf_R������iY�~d���~�Ϯ*Hl8��I y���C��뤒��q�M���Z�̑,0�����^�Ƈ���I$� t>l6X}��ñ[z��t;����������Ġ�	��ؖĻ�[�&$����rA;�����Htl�S��ow[�E��1����8��f�4grkZH%9��c������C��`&%���m��C��Ƅ6bI#A�J3Î�}ۚ�n@���}����6ۘ'n��I�G$�Ak�m� iѧ�Bl�o�=�5�Hѝbm�C��6�a��t�I"�� t�C���C���*�瀜n�<�#��:��HZ��$t�6�BB�d�(��U
�  6��á��t:���6���56�&� yne��ww�t�<�����nx�U
�s�v�]��Ѷ:���f��ty� ���&I�0��l9���u� p.�y~�׻��`C9�czC�8�w���oTP�����GdH'#�@��� ��d����HI][rQ t ��TZ���C��]��F�S��	$��a�-��$���$�����0L����Tݔm�E���K� &�&d$��Ѻ�N���C�I����D�B��PV2)���3T
(4�#{c<#g���審�x[�N�;�����bҲi<;�c��s0�KI{��
J�� ^�e�U�I5Ѷ�͒����P�:��,��C���2�&ap�����6��!$��C���ڡK-�I-�@�t:�C����t:�2(G%�$�C���t:���a��wK�BbP�t:�a�ò	$A�@`��I�I(�m�I-�@�$�H��C���t:�$�H�C���t:�C���{�C��Ht;uZ��:� �C�C�
�֒J�/68�Ge��C��֤�T:(t�{qN��E�[�o����
�xw;�t���X�Mܙ������\��?�s��ewqPi�1P�wN� �tHdӜOr8,�ǸNY��oGv�8`���I��@�^@  Py��O�ˠ�C	&��ۼ�vv{}��dI��<"��oWT¨������f���o���3K$,�F��Ia�bI΅&����λ�Q�N�|;0t���x�;>���u9=6Gv�K�}�ٯcVf%���{�k�e�9��OB�yMI����^D�hLi�|A�5m혈���YѨ����k|��p����e܂�4��}���,t�ᅮ��"qAC`��{1wE"��X��$�ۼR����f��L�)����ϢA��R��ۨ($ÇϦ�"|c�L�`�zM�.q�a�p�ś�@K&rE��v��gu�Q&��n�,L[WU'ق0;�4;uŃ��q�~�F�}������ۼ�{��Z�'�hh����\\��4�]�M]U������a)��2�>���$��"Z��
����<�ݙϵ������
���|%(���H+��+�0lj�D��P�葰%�l�D����	�Hڢ�h��t:c��
��=m* 
[�����$��תo �n�R�p|��h[��F�h�AY�^w�+�sﻈ���wBZ��$$y���`�^H��L
���pr\w�ݼx��c�8W���wQlm�lw4�a����������6l0 "0WS����j$��*���r�n�'�f���Zv�JI$�>$�� `�7t6�{�\��{[�@�� �ce����x	rP�S�+�m����H/���'b�N�>�������F��y�ƕ�B���7&<E�b5�S�K��ܲ��'�B	s�"��/���>� ��!,��K]N�(D2z	��ڼ�@0� ��K3�Q�_o�#�����!Ӱ�뭯*�ˢ���9�ۅ���h� t?f�Od]w�>㻨��|�a���l�r�F�#�k��#��������(���Kú`js�P�B�e�����I����a1a��*Xc��p:4�f��d���g��C�s�P��3�{H�.�%x��t;����n��y6�MJl�rO�����_*.�����={�?3�ށ�U���ϵr������bZ��:�Ug�m��:���[��i���2/� >��};y.CY#��:�vo6�J�o�b��,�܊R&�:���K3�; &Dh��R��w�]�J53y�jǈ�
��7�� ��mפ�[���СY������mm�m��=�m���t��#��&!ܐT: ��6{��䦶� �����Pj�h����Z(�$��3L笘�b7 }�̒��£��rK��GJcݓFne���4��	�wrCwe�a���*%wht:�]Te�ř���n�qc��Aڐ M�Չ�Ʊd#qo��<&|�I({����E(l:�:Ԓ	$ܳӓg�ocBm�ͭI/q��~t�.K���� V�~��Y�N���2sA�}ΒY��x^��i�\V	�Vd���$U7 #���-g<W��f<�>��c�N�11ջ���mn9�I���~�}Gw.��ɣ����H;��s�����٭�Ht5���H��:��$$��2@����!@��$���I��>�$��8I'��I ���d�� �� ���5� �!�А����O$��!���5	 0�&�pH�A��D $���!�I>0�����
O$�
���$� ,$�	��X{!$� ��H} I��B�@I�$� n'$�R� M�=��Dc#�D��AU�Db21� 0� H���؈ �dD�F�	����� ��0d>�!�I!�����I#�c"0X���	��!�M�!�E�� �2aO�I�A�b "FF"#�d($ ,	&�p $a" O$ I �$�đ"�`F �	� @	�'��aIH$�BH�$�� ��7 �H@�'�@�a HHC�BH}$"HBId ��@��$�@�2 ��jI�I	I'`{$$�e~�kN��f\u���̜�J�q��CK�*�m!f�J���U*�gl�Gm �`�Zj	pm�Sg*
���۶��V�D�`�m\�����*��X����HK�p�GWTq�*�m�%Z]�H]l��F�:Sr�80ʹ-x�J.ɰp�Cmv�-Ѷ6�q�ml� �.5�f �]��Tک-�� n��8�&��(\�%١WX�W�2�xJ2ܦ�5�1��0Ү`!,���%�6�ت�m�M����*�b��LB���i���L��UW�.C k-�L�&.��5��#E��W��	MJME�kj�L&n���b�A�D�m�J�&����b���ir]�@�K�P�,j���4�0�vfg9�s��9>�� $�HR�� t	 BY'8rO=��!A&s���Q�2�j�X͡D\�k��:�s-�Ӗ#VJ�IJ�5�3��9�j�J� 7uXeѬ�q�fkGX����ӫ�	H� #V����|�ߧ�}`�C��Έz��+Li6kSwZ݉�ID��z� ��١}�,G�[�RK^Bl7f� {�lA{����vˋf�=qb��I�����@{ָ/Uby�����U���ԜO6B��^���wh�,t4J(5�n!�\��4%��6�Z��~���ܭ��́��*�$��k6n���aj���%�]�,2נ{x�hw��z� ��+��n�bGƇwY�ۗeڼ���o	���d�A�y�!��[l9��v��Y*�ɱ'��7R�/u� ��vˋf��<�\]��Z�FM�cN��V �l�˺� �+f����z��7��(���T73p�CƖ4
�k�qf���J�1�
� �f�Oy[4=m� ��v(�s�v���Itw
]�13tZ�x'������k�y{��/[2��e�f�M��X�=��\�����l�;ָ��Ǻ�M�������<��hU�vf~����߳v�yb�[4���x�Rl��u��l6!C���X{�m��fU���V"ەk�1�q��"Kq�� �Z�YB�,�k���� ����f�ڍb{�6�{ײ���hUz�u[Fbx1ǮD��wqn�����{��B���9_(��������f@>^�b8�]�t����S�Ӏ_W� ��-�z� �����4���cQ�=[3RrW��3����
l�^��u�6l8y�BwRnn����ܬ@}�\�����s���
��٫j�8�٪�P�Z�V��vʣ�:+x]�K]�X+B�P�k5�Q��R�Q��j\�մn�Xkb@5��� ���*Lb�[��Tn�V�3ylbMh�&���U�m	fv׍�r���er�2SFěf��~�[4�������tb2���Y�hM��չ5�jƓE���͢��7
0E4�l�}�la�z������{���wѰnq����FhM͔�0m%�C��v�l��ܬ@[���um=�ڋdP�օ� �ܶh�\��H�[c=�RKwr��s�͚l����+f�����f@�˴@-��Q=��h�؃�ΐ��f�޵���u�&�q,����D�%����0E�	�\GZ�,R� Otח�u�ut��i�v�0m\u[e�#�s
��aiZ���es*��0.�I��鴴ڿ��C=�Xgc���`�.Z��錷9��P��Pj���Z\��K1����rN����Πh%:�j��y��-^����d��X�����f@��ĵ�&�7f�w+f���H�[c��4��+�bNRœH ��Y���Y���2��V"���6��N-oV���2h_u� ��:��[4>�:@��V$����y���~���S�˫53�b�(�j�T��01K���,^u�O�/.�C�ųO\\h��<!��ve�p�h]2��!�*����yl������Z�D/�oefܙ�\�UC��n�U�#���������)"��H$%�$Q��'$�B��ǟo��﷡mt��b����4��5�ԁ��١��2��V �{���/��ٲLP�� ���4���{� ^-�|T�e7u�["hS��Bߟ��,����D������X��:�f�����&�2������<��hw���Ĳ��{�rl�n,2�8�D�s3]�+�o�ܬA��d�z�y[4���ch�z���m��n��v��V ���}����ƒ�a6n�F' w����v33�fg������ {�]���ܛ2D��y���l����<�n�>]U����14��sT�r��}�ߞ��a�u���k�9%+;TDc�kY�s����{� ^�`x�K���`����'t���e��.&����լ�=z̀}w��������{��Dz�3�m�蔋q)3R6��A�ِ���yx�i�������Z���yz݀r�4=z̀}w���U��ת'�E���H~���km�_sf���[.j�T�כ�ZήSgm�,�v��\ma���h�eV]�&�\@��mk3�$vq��e��+K�!�`d�%���K�F�4m�5� !�Qj��ʍ�0c���V��5��lrፔk�EDq
��<��ئpॅ�s�'9����a�Y�M4�M�Ҳ�*�r�>_}�kc�ԡ��Z�QGi��
�$.�Z�M��g߽���>W�����:��3[Swd��Ē�r\��	Y�V�:��P�u�{�X����u�v�lN0��l� �ِ�[4<�[4;���.�	-�����݀{��{�� ���4z��j�ri��f�EJv�DD$�=7nC�7f��̵a�BP��N�3^N��SSs,��(�m�>����W)�iHd[\BV����k-F�͸9ԍ�{�n�}��=�t�Kn!	n���9$�3�be��3���QKR��VcV-n�����лG�b;&�xli�*�i��ͬJ\�ZR��NS]ŕ��q����rL��Dn�Y[���
��V[��@-��{�X��ųC���늕ᚒpz�lթ���?�g��E]�ֿ���٥���M����^�٦�=�t�w�:�ޮ����0yCl�WUcwe)��vlD$�9�6���� -����[�����{z֩����ﻃ3�ۜ;WM6�������M�����k7r}�_��γO����u{״��mJ����^�-x��l�s�yx�h|�݀[l�{�pZ���"պ���{��D(S	)����`u�̹��U��Z�������������4^������٧�IvQn���9��vh[l���lA�T�Y�>�J�����#���.�C2p��YX�4*<A�
�b��޶�	-z�g������4WY�{)t�Ѻ�M��HţA���V�l�m2�l���}�py~-��2 }�"ۗOJ5���n�� r�vW�f��.�C��2(o��fiT����,s2�'Urͺ<�_;xrp�,���Gpfsip�C9��Қ�#���R�Dh%��4i��ӽS �5#!���ė�!�,��p`�	�2�XPL*&2DB���`�	K�����Ƃ1��d��f2��G�����v! ��3 l�܉r��d�#m��H�H�#�Q�DA#["G���35$3SP  Q,�2��a7LV$T�X,&f��b)���m,$߅�F�����E"�LG+�H�5b�R�a����*�$X��!BHs�'���%�����M2�ʹԲ��nx:R��ge�\��e��o4æ���M1��8�1��c�01�c91�c�hlcƺ�Tp&�#��av�jֵ�kq�V��kZ�1�c9��rc�2��mY�mU�e��ٷ	���!j�lcZ�m�2����8]��-���ݪ@!6Jf�uѪS\���Y�vq42�݈h͍M�l�4�ĎNj
D��6k]FŖ� �gm]X̨����4�Cq���������a�&(e�`-�$�!�n��u6lk.��9�җQ�4EJXbf����k願�\QWXcJ�4�e�f`xi��J�RU�QV�F��y�ƪ�X����7��{N����17(:K-.�4����&C+��� ��jK�f��4ږ�Һ`©P�\]�uu&���F�c����j�V�[h�5��ˬ��5Z...�+��l3a�m
jP��m���0���Pդ�(�T��1�Wc�6�	��e6n61����3�pkm)�VX�И����3#�HX�k���fl��3��L�3[cR颋�[ilX���3e�[�\��%h��UX�mh]�h�P�R�DéH�+n(q�\fׅ�M��B�m�-��gK���J�ڋ0��minS�[Aƣ�����֠2��[�Kn�u3V�ź�5����,�d�=�$!��BC�����	Id��I'`r&�'����}~�x�_���?{ڊF���h=M� ��lA��+r�vW��OIvSO	݈�^�|�����\n/R*a�-��s�f	���T�[��1b��u�@���:@��ebz% ދڇh.@���al�כ���f��:@>^����g��C˪���_�nRCr=sS��p������Y��<�����i���nF4���s��ųC��Y���Hi[X�69�Q��Ԣ��X���`޻b���ٍH)�CuK��1̷\敹�<�&V���M����6v��Dh�� �6mWa�ΪP��[�05�bˈ�El��	�j3l�f.�b`�[��P���P��6�A��vj���q ����0��M��53��F�K��(�6�jrr}���}ܝ�}ź�3[P��F�@;޿���e�$me@��ˌ?�{�oi�Tm���m
��?�����: �x揻��n�lOG��Ŧ[
��n<e��&�!li����t�z� >�m�9^V#�w$"���r~#Ǧ� ��Y����;�� >�٧z��wJ��-ֈ�{� /Z�*u��yb�] g޹u�l֢��n��r��@}�\����m%��/�jX[qKXB9����.� y��y���'/ϗπ)X[��Gb%�,��l��虧O3wC���9�_|�c���T׿K��	���u�9��v&�j�Y����B��-���a]`ՠ�4�NUeM[R&�v^)��ͥ�40~;�=�#���f���X1��B�$�9ɐ��e陔�%����2醭p�����S��ϯ�x��j�I/�k�����m5�6��nK�m��k>�Т�Yܭ*�m�k��ݒ��wu��G��8o�	f%�� ��m%}�/�jKݮ�$�_y[��/sLH���qMi�TԒ^���I{Qlm%��/�jH�:8��=M�}���<��y�~��t ���;�� �5��섵�U���f�:����=��K���]�~�R뛿�$��[_��­�hr�l�eڎ�tw@��߾b\�S"HK޵ϒI{s��\wV���߾�E���h��y\y�$�F�����9ܛV���U�����R�g��oV���uA��Y����kʡ�K�Z��	r�L�/\K�����Y�o��y�7�����G���Z�ܽ/�6s����7�fW�6�5-�݄sf'���J���I~<g��H|�.ف5΋i7*na��UJa$�U.~�n�|�o��Y����f���y��a��y��zy-��Z������j� �4������n�δq���i���˾��Órl���X�lZ�_[_�$��vd[���ڗn�l����'n\�����&q�>��z y�}���s�BI���h�I$,�[)D"�$H��@I��������TϞ���J؞۴��G��m���]����lͩ=n[o�̯�m���	'��s���ݷ���?�f��r��n�y��<�
}�� ^ɛ#{L�qm�Jm�ŹQ�֢Lژf�0&�e��eԗ�XX�%����䗲�͠�v�&��l���K)iCF�Vng_�/m@>���� �����̼6#����m�^���c�����?�������n�����.���/�Uv߳����e��?k7mo����s����7�������Ӹs���o���m�����G���=k�􍽗�M��aTEUS���ē�*����ʫ7�=nX�o��ϒIwY�	�74[���bǋU�s�v!�v3��.t�d�ՠM2m��4SacX0�ێ��u]���I��S�,*�ܤ K���cJ�cځxW4K�X:�������E�LU����m�T�j��*ۃ�2L^S-kX7P���Uа���A�{����?�~��dlݹN�j(=_}��yK_;�1tfj�M��l�"N�M�T�m�JuU4��f�g�����˰���M��9>��͂��vZ1p�8�2������.��y/vl�?����l�jLߦ�o��~����Fگ�[{���0�z >z�皕L����̶�r�����M^��WZg��f�c���d)����� 9��Ͼ��!B���l?~�wm����|�Gs�)+��������?I�m��?~��6�}t[m��d��K~K�S����Z�����47�y�����/� |�����]���2պ6"6�X�Z��)�r�-ӕ����=M�N׵D�^�L�}�g��cm5�h4��@�Y��6��h��*�1	���,���t�-*ܪ�� v�S6X�IV�ې#]���m[,xq��-R:��,7$��ӆ�e�nE��͎]v��'?y����{�=��|�g2��r�c��(^B�]�ͷ����}���m&n�y�爾]3���9~J�.��o��o=4�-�Oϼ�'�9���O6��cg���ޝ��Ceݶ߾����[m_��{��~$B@`"���~>����I�r�Y�L�3N~����<˧.]s���B�!�}��iݶ�����s-���o2�~� �"BQ*����~�:�����������ށ��}��ji;�C"�u5Vl�`�0eΊ��K�B%�{�b D����~mo~����u�E�ukq�ݟG��]Z%�r����f\�~��BX�_R��m�5׋%���̿�m�-y/$�(�������~��uU.m��7%*�m���U��Q��%�Wv���Z���p�����X^ǡ P��}���.f�0ַ�o\[�/8���]�o�v�}���%
����V�����y�紾��k�N�2n�{HP�Vg���Ͷd��\�m�vs�އ�2�s�ݷ�ߏ�]-�s��;>P�΁����T���z[�+3b��
n05m�������R䈈P�=�7Ͷl�����ٖ���>}g��ɷz�W�Lj��6����~����'Y�ŞA�6���/���̩�d���ϖ�(�Q����~��V~�������Č�s|��}�{]� ��	,$�����s����گ��[|��<�I?0�$D��m��X��6��h[N��z���?s�m�{��wn�Bz I�'�HD%�q�|���g����|�H��)T���k���ц�r�� ~d��`�H���/�2�~����Ko���[oTB��0BH,$��!�}��߹�7���f	$7��4͓R^��|�?Ӓsw��~+���ay[��p�m���,t9\�D��'?�99�0$b@"�� �v����V߿z׾�[fv��m��<�"��O�鱿�¡�euA,ƅ���'$�����L�8sN�=����n��̶��~ϾI#ں�I[��}��J�@�W[�֌˛�fGm��<~���$�0$�HĀ�^޺?o2����[m�>��� � 2HL�~~u�Ӭ���[$��U7���^�%���⯾z�?A 	�$֟�t~�eo�~��|�����r���jKN�۽����I�H�����u~�~�v��Ͼͭ4FA����%	Ia�IIK!d���o0˛��nKj�q��m�kWlZ+r&6v���b��uh��T�..�L�ie��{=�s�M�G&��b�^<8������P �٭!#TU��M�Y�Z��v,��\�R���b�\aY�[\ne��&�k�:.�uk��'�$�Y99y,�C�������,��?9[�������O�}{mf݄��XM�p�C0��9
��ѵX�H~��(�'����گ�w���Ͼ�����zKw�Y�U�:�nU�5��k�Y��k��I  �#�W���|a���`s�V��9��� "I ��$d��K���������4���`��7`w�K/W�I@FI���#$����4~�^߻�6�ϽϷ�� �$FB0	BMa��]������ ����>�ybz�����,�xe!H�]ʷSjd���6�(!�D
 L�~���U������h�u�ЈA� B3����2���16=ٻ&����V��s�����Pjfmi�����ٖ��f�Z����?�Y��PDB��}?���{ʬ��Yl�:<�Ku];�o~�hB����N\=�<���`7	Lyְ�S$9��X��X%(Q��4a���s�<�i.$�R8	��Ķ�A��P�*� ��
ae�DFH�ϩ57�a�̌H�,#,�D��d��7��>� � ��Ĳ%��C[��D�9&oZ#˄L0�<��� �_<�a���n�jh�Pդ �!�$�2� @bɭ�I����"Q2KS߇D�A�`� � Č`,EP`	#*(�H��J�"X���c��=� ��Jn�{"E�#���1FT�Y����`j,V2 ��dQ�N|�a�O& X!��[ ���&��&� �L5"�	��7,#"  ������o�h-�nVX1-\8إ�%.m���l����
��*�m��am�mmܴ2��/iު�EUP�;;ef�`�6mAF*8ˍ�m)MfD�*)+��1tЖ�ˎk��CR��u���8ō�n	p�*�k�u�B�6��6�2�ԅ��p��q�c��1)��fˬ#3Wr��͕j�j:�	cjd��m��5,�RR��c��[�	�ԉ�sU��6R�GPB�\�Dͬ�q�m��]v�!��W�-�6HMr��R�3D,n��֪�]��V[u5��KƖ�iu��yC,kLUohז �����u�	)R�fK�2T�5l��UV�f�-��cij�e���\�D5KB�*c2��ٝ�5֜��@���C@�	� !IrH|<��@ �$��	쇲I�I����kZƮ	A�ԃ2c+&���ɂT-6�X*,�
l0��	�+q�i���'u�e�a��X�ŃvA�����t`X5��ͬ-�J5g������rO���Q=`{���<ː>�NlB�$<ҽ�������ff淼m��ul9ުYz�/ "!T��������@w�lG����sS[#�6I���;K-�9��ި�$B�2w��X�듙Օ���M\�S*j�3l؈O'��`gv��w��[5$�DL�o���������p��-�~}}�j�;ܶ�u��A��3����Q�sCh�USsOTD}��U��Km�r�@�[�_�6�lNI��c���3R�Y7([�h���$�gzgx�����}���yu���݋���oz㲗�1�����Fnr_�.���䁣��L0�B���A�1�C[18Kc"#��1c�7 �S4�Ce.Hf ��� �!``��FFXBB$��y����w�;l�'�
"���O��4�ɺ�I�Ԗ�Խl��.u%�(��MY�U���/[>�,C)T���˦�6K�6z�����,��l��.MQ�=���;�lς������h��I����Ӵ)�ޒ�v5�Wg�431�GX4��l]��Ǟ�Ԡz��U�i������i:�(���nm&�+�I?�(����h�f��;���`|w�t�e���O� 0@�=���Ώ�����_�5t���wq�f��^}���I!�D�c#$�� ���}�u���~����k�z�m���ƈ��U����⾞}���rd� !��H���2@d$IHd$@�$�A H�AH@!" 0@ ��e�������Gq0Cmӫ�v�kk� ��$�	$A	�`�#$�I �k��|?�U�����+�>�[^!'�0B"�B"�B$`���w���z����9�owz�D��~� F19��ۥ��'
8!V,3%i�f��sV�4��O�0HI,�����~7� us2�>0����[s�q��F2U3�".��u5R���r�;���c���Q�y�&�.���wNPZ�U36ݞ�{�"Xw�:����Ձ��Z�Q�B�S8c��.�����ˤM���������BlᙷA�ݵa�#�Rʺ�aN�i̖�(��{�;�}r{���;٧z��*m,-gW-W<D�A�\�ٵY��3b��Z@tur�[sVa�]L,ֹ\���KJXp�# l"lhˋ1�;m�*M��csmj����Em)V�DmgS)�֘е��4f��j������؅�����fWY�j'�:O�HC�����l�����u(�����d�!��Z�o�������6 ���ĺ����,��A-���N���3O~���}rs+;��
�UM�vl+k��4�snɓ,�hޤ���� ��:@����?f|��^�ȷ�k sAsvʺ��,���z��̝���V���D%MgS�iJ��V�m9SUWa��i`���� ���=����Ǳ@�SUWF�(M�v�9�ZX9��٪^"&s�>�x�'��U%\�nKT.�|>_���=)��bf%ɀ� &̕B��j�	e�m�������-~�$3=^,>˓�&X3K�w���9�e��Xj싚��F��B�� ��v� �^emH4h�����vn�d�P�F�����l�j�t�n�35&e�h���2]�5���7+ԝG������o��^,�}ː������BIrû��þ=1+�]L�n�mPU+�9���J#�L��Ձ׆��,y�&w�**e��#������Y���X�石��
?�*�o��~�rp�KĜ�W.�n��k���$?!d3�������O�گ�{�n��'�$B$��w�������n�����VR�&���Ǚr�4�J�ks(:���u!���P��k6	��~�{m��������ˍ�F7#�`��$b�FKpҚ��[��nvH�0�""!M�"N077�`|�w.C��,���#@�i_���[_��K�NfU]Mԫ�N�݇�ܵ|I(��IL�yy6Տ�rs)eꈅ�DBU=�/!��'N�lub&�מ~�����脗�(J����X������
����ڍ=��@{ݕ��h}ź������=����o�Aw{���/{o��gݠ�[�v:��鈹ֻYjU��R�[uh�_�'?ÐDG37ՠu短�s�a��T��N��oE�!z�]i[�nFu2:�rU���rw����VV�(�\�Ǉ�rn7�̍�M]�h�3[U����I~��� �K�����/��K��9��Xubo0D���Ӛ�ݢ�wW�>~ٵ_���m�I,����I��=���/[�^d�5E;��t��
j��DC��ݹnm� ��ʰ,yf��zӍkջ7u�D���'W��ZWV�
\!�b�af5]5�B���$���~��P��mXyܫ�'*f*���?�;��ɧE\.�.�hF9�$��;�7w|<�D^.Y���١��#Ǖ.�oF��Ԉ�� =��?���M��R�`w�6��2����L���Բ�j��c��6�l��u��6�yb/�iܳ��V���I���6�|ܵ���<ې8�2�-/��#��o���浚�p�W;�׭�u�""�\mm�-(�h<1�5�ce٘�^2�A�!��K���$��Z[+eȴE������&���;��h�&�a�m�++�nkpb�ĥV�L�(���p@��WV��[30Z��q3q�c��rI#�J#��_��u=�mN�[���u7����=��v�B�6 ��0�+�c���b��"m~��������/[�3��o	fb�
6;�-�����I!���榾a��܇_;�`}�����9��M2�*<07�������W��B��K��܁�ݫ9�Z��	yB�2��
�GJ���ͅ*�������=y���,���]�N���5j�˚w4R��j���ͺ�7j���K-�	���ܚwI�˕H�5nmδ�}K2 �F�x!�X�$$n�6�A�����c�����ң�ܝ���3&��v�[8�&1L�ɷz|�i����=�s��̱��m��,��j:�\YE��К].���*�C�F�1-9�!/�ָ+r͝��t�Q��6�CcT��x�s��.�$ym�s[3K�")T�.��^f́�v�[����[\{+��SQ�G���[��_�P�
��}V�ǭX����G�*�3��d��V�S�RM�g���|��f�����ΐ3�u+�&ܹ�D�*mIWF���gn�������2���(��{羹=�l�)�**��J�6a�@<���h$͵�q�H�*�pF.s��Ҥ�Z`��F�����>�f@>^;,��_�F�m�7m�t#�6�bĉ��òB�Bo��y��k����^>}�����c��@�vSRxؚ��!	�w�y����! P��A"F�
XT�Ia@$B��B�al�p� �}l>|���B��"D*�c[3੩*�U���J���W�CL˟�
7����9כr|��̡��M޲ԣ�v۽?ā?�����j�����W�u����>�櫬L�޽Dٻ������;�JLN�iU��̐P��h��4a������	fn��:��W!��ܹ;��Tܧ=sG��i���!��aՔ:��UC,�>��q�ǗA�r�؈��`g^�ɋS{�%��ꩦ�5SrΪ��"!x�!������~���V㕺~�Ƥn-Jf�z����C׵�Q�b"0H�AP�����k K-�,3QF,b܌-��0�A���b =Xl!�ɚ��5���F�p�0E.�M�HA(�r	���nH� �PVdh ��R)`$dF1R��	���1F`K ()%�L�U# �`�� 2$�L�A�&"�i&1�t�1 ��4�2��>vՎ�����$\;9B�l9[�c(c&��5a�Ζ��Yf�v�W\�p��q.��Zֵ�m��kZִ�cɌc�01�c�U�F��Ÿî���SU�1��&1�c�1�6����W:��lc#���M�!��Xj4�FL]e����K�5�hff��h݅+E�.�&R��h��f�M
%V�e�y��1��nm �Y�B�0�tHjM-1�EsMWE��3Lifs�JEřr���j�B!�V��5���S,�[�v���,��E�i�1�5��i]0��jl�h�XRc](� l9-Ͱ�L���s��R�
�9�dV�dR�Jك$�C#f��jb鱌l�1\���ͳ82]f��7M1N!�F.��\��ͥ�۪� Ap�54E��u�j�cL�Wc���UyXL�D��SmnF�k�j4�؆�;q�Z5�&1��Z�`�7j�Qn�.�\kX���la �3�.	k�WUؐЉ��+�;��ɢ5ˇ%v0�65��v%VZ���ؒ�QJ���<��l�̡+4.���j�Z(YmIc+�D�F��#��q�mj.��ĕ�Q�K�X��+�Lr��u�ZJ�(�<e�#�F�s���k�%n2��9H��s �[�T1k�N6���2�0��P5��!5�ͭ��k��&+
��f�V��H@	���H� `@z&� �	$(NI �HvBO̓z{�������oO���
iU[r�w$�HX~����Հs�v�9�T���|�͹1w'eȪ���-,������ 
,�F4���k�����i�5�p�Z]��f�}��o��ųCמX�]R�ܥסmu�u-��Vhڬ�؅�wjf�_q��)e�9���(��(\�;羹;g��u2U�J�4�Z��up
�+w�� �wU7��Z�e�Ћ���I�4������^�T������]�\mͺ�D\�n��l$��ې�b�����~���Q�C RW%�0%)BZG`�!��r5(H�bJ	+D�,��e�VI��&�#�ffKlKm� 6 YF�e#d�B�d�!d������m��ѹ1B�5W�)�m0+6\�`Pvq���S��q.Y����5���$e�E�1�&�vG��L��P-]s��K^!8ԳUʉ���[�:\Fm�aBn.4,]�,����ٷ*6���(���̻�S55QT�&�!BN"!O��[s�*î{�na���_}�nŴ����$�f�KU�*-���iʔMU&��.�Lݐ�e-�_������|Æ�^�㶋6*�j�T�0�fO�r]�h�k~{��� �� ���Cױ��������M7&�� �ų�3�	����@*����f��.�Q�S!5���B�|�ܛ��x�uC|��V�ݫ9Lҭ�q��n�܁������V>�&��+]ف�[�v�mN�t/��wX�;�Gj:m�v�CP-�ra�����-G�vX��z��u6�F�{���5��!�	2�"ɀR+$@��Hk2S��sWZ�֭�KK�u�ɝ-Z� E��4�l�\��nH��,Ġb��X�V��j�3S`,�U��t�i�CDj���[��m8X�Pח&/���m�6��ڰ��\�3���(���ͫ��l9��]��,�i���3-_�6k�z�C�3f��{K/a/�R�|y�-oVǻ�-�?5 �]��
��d ��l@}z��w.k��n(�dx7a�
&{�}r�}6������^;����ѭq=�Oq8��X�2v���0F�.6��%�3	�\�I-�橴z"<���{d=�����2��������=61����1H�c�J�.I��ܫ��V�s�	/(�\���z`S����m�lٺD�^�r�<�0@�	 IiH$d �"A�AA�FE!��D$�2@�?_��mN��|�w/�D��VzY�MT�WhR�t9�;��V�vr��6wsj��ꥶϻ��95JUuTl�տ�_�D+���:=��X��t�����8��bxlz�,݃�b���m�rH�ɪ���GJV6��m�u*�3L�� �SST'M�Q���~����L��m�츭0X����e��]�؛ U�B�.��\���1R�`}�2�1�2}��!�mx������Rlj8�Ԧ��<�� �v��>|;�!���w���v�jiU[v�M�5����^�Y��b_u,��]f������P�yC�q�����+{���<̛��aaÏ�ܭ��lq�&-y� U�4X����FLX��+n�Ks5��PI���] ������]=����:�E
wl:�gZ;�-z��M�����
�u�gr��Ù��[9ִٙ%�H]Y6�f-{ {����-�x�M�����vu���n�nlŚ47{����>��v�Y�W�f�����Ql(&eӕa��3/J���t�k
�I ǩ�mP��m�W5s��CE�ö˗h��ʖ:�yjU���ͭ�p���\�f���/*X�ɩQؖ�Ѻ�49���]���&�ܵIi5%�A0ZUm �6�˫jXq�ka��lQ�M.pd)�Z��ԙ&`ܪuL��G"!)��̹�y���UF��-�c#���nȒ�F��mr��:[����+˫�n��^=�����K}�U���ƬwN�gx�\�Y��Ûf?ɚ�D���0�ųC��d��������є����Zjd&�lF� �ۖ���Rh}�� =��?�g���ۺ�{5��������m,@_+f��l�������MM�P�j&(N�0����n[4/�:�N���k׻�-�a =��M�6�6լ +40��X�4��UEUM5-���u4��;���w)�l9���K���Z���Ǣ֞5ql�H1��ޱrj4ef���F�ˮ� ���ي�h@�e��i*n\4�eiu�m�؀��Ͷ�l@P& �\�mv��l�ua�%��cn44�hz�L�}yY��la�s����Ğ�MZ4�f
}�Ԛgie��;XXrp��Ʊ9�U{�# �Ĝ�ݿ�� {�١�WH��f@�y.����oV)�������w�����r
$��km��ZJz6=Q�M
3B��� �zM�[�-VP�Tw��`n8�VcL���Bu-K�����fNk����>>>�*=�ݗM�oy����U1���7���O�qf@��܇��Y���������5S�U7w.�Gx�����n@�2H��+�P��+�����2�cΏ/�|�Ss�k�b�Ʉ54� ^_��C��K6"��{�i`כr|���eP��qb����@��ɡ�s�{��e��AbZ�s��ֶhUz���nmac�bnnnj���M<B��F�1��g��� u]f�z�@�ֽX��`�i���l�9hl1�q�si
�̧@=�}�@�ݱ{mP�n8��񸔛zkz�z���ܶhUxV ��j�sݴ�Lm��y4�OZ�w��ױ��,2����K�8�v�|wm7w[4rc&-y� [q�>����yb��T�~�5��D�{[�<��>�
�ev��ƈ�,�:�*;l��T%��\����_������yb>��(A���z�@�\ڭ��Y��o7l׮ }{lA}�X��ێ��#=��b�5�F���ǏA������4>����W>�\C׊nǩl�wS[ �v<�}k�^�w����ڋ��r(9����Y�?�%��wu}��;���=��@#qtcr��K�\�gj�x���l.�vuS<�@H1ղ�ц�Wj�i�Z�yT��75�B�i�KnhCU���,2��1j(�t
���K�I��J�\LJ1��
9�EU،Ў]�p���k���q��d�yM4x�к�~�?~���i���c�SǳT���֦���~z:w�G-�4�mHk[���b��&�+�������yb����b���jj�IM`�[�]b�f�V�h�2�dA��,@}��{��=���S������T�bר���C�W� /��z�@�������!��""����� �o ��D^��ͺ=[��L݌dA}^X��T ��� ����e�ņ��5�]l]�}��m^����X�.j���+���.3d�kuЦ�jG\����V����ϯ��Z˽\ےjBCHI�2ȒX�
�&�K,}�	�)d���Xd,�� @�ad $,�!�d$��"PK	 ��A�� �J<<Y�sm����Qc�+�+�]a4��@!��Tr�����U��UEr����������
�����۔��#1`�\pҶ�U[j	��+[q(#�D�ҹ�m(�g����$!�ġCkv�v��8P3q��)e͖�-v�5DѴ�p;nXU)w+�@Ʈ�DBm���S�w0�QyZ�X\�SG �2�vn�W]ªmA��X�-�r�B1.׎D\Y��(I�o2�XX�GU�(L���Q� V� �14�#����(L�Yp�5�e���;&�CP(��[��v�f)�4��jR,�t����lf��j�-5U����T24p���ؙk]fci�B[�����ee�ha̤ 9k������R��	p7L�H� O�Ё64��}!! � x_K�GXZf�J�Xj�Cb�Qr;[s-�	r���!5e�a�ԉ��B9�`�f��mvuZ�lA�s@�K���5s6L5c��GGp��L��r������Z�D�� ��,A��:�/%���\c��LPp�^X��>��w���w��^�����cj�9�������$����;�ň;�K�{�a�Մ����wW5#n�e�TDF/s��4<�/��>�yb�����x��z���Y ��yb	0R�����h�hዉ4��-I�����Oyu��k�w�����aÞרwl]��\��y����4�7[X�z5�0�o��;���{s��>���8Y�bm�p!�W3u^?{���(�##cE��D�����"!R�(�3d�rՁ�꥖��r��r3����m5o�;�ň=�yr �� ��,Ge�o�w7u���ǋZsC��n�>�yb���;�́O.E5�ԑ�И�ů yu��hސM
K���eM�ҁ�L{�6�{�Z͟r��]��=y�ȏ�P����Mh���x���kZ8��l8�/@��~��v�B��١���g�n�kj:)]�WA�r��(P����mX���}�l��h�[ո8�xLZ�\Ͻ���{�n�B{D��A�A�	D�ADD�E$9��/-X����#0y53%YV�HwB��RI'���`�ݹ������́��R�[�В53V�^��_}���	�h�ic��G�"�&��6��]�}�߾����R�lw��Ŝ�2Ju$ܹ��	�2�	�3�bBx��k���{�/�Ъ��h}�� =�l�>�m�b�cKf	�k`�Y��[4���� g��q_ێD�(��=2h��{�̀}�γB��٦\��u��	�n���+f��]:�{>��s�NC��݋�M���`�q��Ĳ�8٪jr̬��B�q�:�^m��h�5�H8��J� 6���X]���]V�S 7<�h	S�SI�f��aM�\�2э����c��롕4cǋ���V�L.µ#�� 4&�O�D��^�=�U�i�غ�{�jj�&��dо�2��[��s�K�������`�՛�75��=�e�t��z�����hz��;VNrD�)��.��J�֊�n���k�e���o���޵�>��g-�aspd�0�D� >���>�١}�d��q@�����=[$ot��d���d�ު{B١���ꪸ�m�PM�6b6�m,Aױ� }z����L��+�$��c��[��@>���c:v*�#��l;+.���gUK�Z;J�-�6{�߯���� {z��J���֋��g�M��kj+�9�*�q�SiIey*V��YKm+;&��3&q�s*�hے�fD]A�)�����)���x�!��46�kC��r3��K;ŶM���Y�[�8ъ�C�޳��>�W ��� ����}��S�'�q��<oP��]f�{� {z� {ˬӯ~�=��9�OZP�z����m��/v�h�k��v����Zشՠ���ِ�����4���?D=�^��\�U2f����D�N��/χ�z��;��
���b��v��ǋm�.��9�������{���R�4�8Y�f��m�١��71��Ɉ6#f��v���p��,A�u� ׫����[�l�t;R���v�^Dw��%tu�e�ܺ����ˊ��w7u� 8ִ�د]�}�������v�q�SY����1`�<n w�p��מX����<R�C[&�gmfu��=��v�#�wR��;e�M���˚�F�6�P&�55�}N���]�`z��z�գiw^��I8c_	o�mΖ`e��;cz��&?�_�� ��f@��wW�TM�����5�ů�>|:��!*a�ݫ;���|�w.NA�T�z�rd�x(�l�W� >�y�'��Fb5�U���#� 0	$dd� �Bh���C)��F4�IR2#�H��DDcdc�(	ƐH�		���!$�:Ϲ���_�ٵ�����u!v���sD�٭�3j���[l>|:�h�W�/�]y��d���|}�}�h��B�EV2���`��Af��Yv����������s�yu�g�M�bm��o���fVPt6�Y�L���r[�Y�����`}���_0��[l\깨���� "-5Fa4{��w��>Y�cb�.u�U��צ�Q�D@}��hu�޵L��#�b�Q�p[���<���~;���ߞ������O;�6�9�Ƴp�Z]\�.iR�B���Vp��2���%Z9��t���u�#aI6�ZY�-��B9#B:��<���	�@���ѳ��LU%�u�6�8�qv��%�N3Y�4e���ͫy���������.�3���''o�ߎ����,WRf��M�i�0������8v��e���l�jB����m_�zf��ײ��h^��~�{w}4�n��#�-�qu\i�΅���?}������v�؅����ɸ�AK�R�I�b606�ΐ�wX��\�a�����q`�X����F�D`}WY�}j� >������+�$��cnx=Y ��Ԛ�V��t�|���\�q�6�1dl7{�����@��
���	t�f"@���P!���ie�ͩ{��٠Z��^Vd{�^�-l�I�{�+Vl; �4h�J�r�c��1
]Q�1Jm�H(İ�R.���e.s�l$� a��iq�ˌCn�rjiG�䜟�:�6��&�4a֨�-�C_:���v�[f@=�Τ�>��i}�F�=��D������Y�{�+}�� }�٧�����M�5����+2 }��ݶ �d�[�ƍ�s�ѽ��u��� �x�4˕��<,���zb���׫Q �}=����bu1��B 7e�ė^ab�A�,t����h}�Vd ��lGa��e׉�nnlXچtÆ�,�mK�VwC�ِy�٠}ˬ��s�x���&Suwr+wNh��3��/�N��g�߳>��� =ָ�]f�z�T5�5��CMɎ }��h�lA޶d����Nͨ�ɺ�Qn��!��yb�����,����y]U��ܒ	�z@��41I���pb��m#B+������b�I�z��I7�{���@�\ ��_}��}X4�ۻ�9�+�)��x�5�4���lpw;� uV�w<���v�B�n�8�ķC�,@}mp���'H�L�j�=	���� ����6�%��r#��(j(1
S	�Lc���A�A�$>�R�a�¢5� R��-��F	$i(4��s@�k%��;)AD2Dz3�
e�.dll0�#xH$50�F&a 5���]�d�Ǝfh�F�!��*Cv�fo0K2�j!@`�""1s ��P�'4����`̷�1a41SC��, t.\�-���p����ur�q�S)E��ȻT�1�c�1�`cð��1�`5�c�665Qʋ�ZcD����T�1�a�	�c� �5kZփ\�V��e-�ĩ�v��	u��D�`�Xf#�)s%�ʶ�(�j4n3o 1�L�n��a��)5#5�9�v���-SSU��4������d��+�Lf��U���ZL&"�:jm�V�,b���.��s]R$IV2��m�V�	j87�E��,1��[��L,�Z�LL.aj�p5!e�,lMM��[M@�@H�M)���l��Kk��ui�W\�*���kź)%\:�P��j�Dj�1uE�Z���`�&���SZ��J�W�`ѕwb,1\��k�5uAҷdSFE��%f�1r$��GE���F������&FYj��+s��2�x�)�n��m��Z�#-[.7D4`�X-��L7
mv5�kZ�
���ɪ�՛A9i�U"L�ٛ-�16��Sj�R����6�k���15���5r���n�[���,�(�p��\Сt��E"�]bj6������%����&v�U�ÏRS�N$L��%�A+@v�XnZ�6��̫t�����ba�T�4�#�G���;:�(�lsU�.��[����I�Ia$��=l�C!� $�	<�7$`�䄢"1Gy�U[v�y�'Nx�ҙ���M<Q��v�U4>�f@[\���LM��Z��[dо��{m��t��\*r�X�E&�[�KMX&�o|������f�zِ3ܺ���Q�?/��wX���6��8͘a��=�f���X��� �^UM2妬c,swET��n�9��~I(l9�6�7��� >�W���@�jjh{�5=�ýl��uN }ˬ���"�����֥�M�h(��8�l�������om%�n�7Q��sW9�Bh�m[�����v�]UK��pK\ba�D�����@ͧ2%��ơ�<f!�fu�@��	��[,�k�Vc(�� �	V6�ͱlo)�f�8�I�P[�v+�j��Q�뵭������sD���D(W�1�ܜ��)�=�:Cv���y�ߞ�s��6����r�iS77A��u�Sfnn	k�'����] ��vi�z}�o�ӽsׁJ֔���JF�������bm���yb���@��8�l��\�7�s`�n���F׫�wp���]f����g�뚴ě�M��S����h�\ޯ,A���i�qn�Q�kV��u�>�f@�v�׫�u���b�Zm�Ș���� �up��������[�(�B�
���@�u��Z���b��������וM��콚�]��G�~?~�� a'�@�<+T�X�i�Z��,6�837m�F�-tL7����pH�mf΀�KKt��\�\����uYHV�]Aܡa��A֑G���N{�JvcK��ڈ�@���˪��_0��ܹ�;��w2��%����f�ݠ���]��m�!�.���� >�h�\�ΐ-�Z���&�~��m��z�����/f���6��r�ֽ�FۈF�[ =� ����:@��4�b��*��TCx���H���A=-�!sHP6a4\�#q����g�vUt�W ��H_a�d6���q���4�!-9x��?�ǂ�ֱ��-ɡ�[2 s�9�
�C���a�3UK��f��R����ѵ^}}�}��0$Bw�6��ܚ���{�]�q�W��M֚��{�r�:@>^-�*[�C�d�jm�m��� ��D^��w���]f��V�-�ۯtI9�r�g@���}��w��M�͆irl�q�B�ۍ�z�jQ6cS%Rl�M���9�����rq �1L������e�U��h�Qaƪ(*hB���j�9��[>c�D(K��ǳa��"d*B��-\�M`w�2�E3�͵`w�I��w2��d`����Y3rb .-�.:��������s� ��،����6�ȵ��1&� �N� >�٠{�١���=˪y�Ĉ֒ca��qN�0�N���k-2i��D-�n�kMn��3qb��jBϻ��T�4>T�&�p��Ǫ%2%��ޅؼunm�cF���@?~�b����u���؊\]RǣSSC܏D͌>�f@=� :����,G�L�J��S7H�#�:�B�� �k�|���}�Ks\xc��D��c&���p�]f��_�����$�{m����ưµ\�g1�Pq���xV;V
%�kv����
ٲ�4ŻeJb�50+b��C@�e!l8;F�.ZZ��W��ruU�Cb��&#�]�gh�Z��c��TbI�!��Ʀu�R:Q%�v�.��2�j�3F�1�X�{�2H����k��D�T!�u�מX�?��	��,3�E����#5��f�LX����n�ˋI���#�v�"�M���y4u�ypr�`��-���t�|����\�@}�_����޽ۑs3djQ5Lw7T7h���>�'H�+f�מX���g߿%p��oԍI�iEzϻC���?�$���/��X����Dzڇ����5N {ˬ������� }WY�vr�\{�jM���
�݀~}�Ż���2�㨍��%����HI��}���hw��}��������]kN��c� 20!�e���2H Ą
��
�"�IA�"%e�� ���|��êm����4Qp6D�n�k+���e���4�˔���J͑�@B�ř��Tv�˶�j�\M	]JG�]`WZ��rU�h�`��6ː����SG��ʫ� >�� {ˬ����z�bǮkk dŸ� �u���1�2l�y��*|�	Z!�KN��5����@>T�hUWm��k�ާ�CX�e]K�U2l5C�m�`w�����]f��v؏x������v���>����M��Q��ZiCYYlҬ0�M����J6�ƞ��v^Ao<���v���Y����t�j��A�].Z�{��i��a z����WH����<v*��l{�5
 (�{9w
!.DBV���Fe��p���e��V�o^����x��D/u�G��@��l@wup.uͭ=q(ѿ��f���^� }ݶ �ܬG��F��{�4�0��>�f��v��05#�+��b�M,\M.э���gߨ|�݀r<��/]�L�xH��Ň��㗯+����Yx�4.]:��\�] w'� >�\2�����{�Mɏ�*�+u��{��9̥�����=�buT����H�UMڿW��w��ϳ��qY#�	5,
Y ���Q��K3��ɖߜ�:@�rꞛ�B	�1��@}z���lAW�X���������4�R-�z��;���wPR�H1� h�6U����[.�Ԧ.��<����<��|�>�yb>���Cѩ����F%Z��KC�dq2/4�jn��?����׫�����_�I�FL�P��fN+�
�s+K;���|�u�{���x�l&�1���^X��]f��l�����;.o�f�5B�^ ��ܬ@}n�:\i�T^j7�l�3U�֠�5Kqhk���x�h��%K��%����3)M	�M�Ͷ�f�c��́� f�)ZMa��15&.D�%e���TqsH���\�u0���0hĂ��v�ƚ!x���KRiqPα��&[�L����{�,9̓SMM��	�,۴<��~�wts�kc �M�ݢ��Z��\�%q��k^����s�=�2��B�/wP��D4ܮ�S68�i�w��w Z�X����@���^�b.��UlZM�7I�&�@=�\מX��������zچn,�m(��F�����}�̀}�X����K�$-�����k\�r�}�r =�\�<����F�����4<��pG�O`Ƃ��i�lSi^#�l��Y�����߽{-@x�c�ِ/�}sF����Z��܋b1H�VA��0A���H��`Yo�2�Ȉ�bh�A�� �3Q��,��̉I"���$`�PI ��1FaB�d�1� �HD��0�` ��HH$�#�+#,�,	#$�1������>�)�`��MI�CFj�]͖D�	5�#I�p@��$A��j"nM��7H �#X�Yaaad''L.��h��H1�IH�A�(F�B�($���`�K%" �2�#)����K,�i�g	Gp�ov���6�`kpM��X�R#H�%#A� ��0AE�X!��ѰJd�Pe��L Č�ɭ���DA�D�ol!��I�F�LJdPk�Y,��L����p��vU��QMv�p��(sVhR0�Pr*����*�l������ ��UVЪ�����fݶT\D)Wfh*@m�V�Q���ki���@a�@�Bj��x9�&�f�Ρu��Њ�`i0昮�sf��xVZ�䔕�%Ȯ7\�R�yfx�	M[W`BR����nnQ���$����M.y����`[](X��
B���ret�\cjf�b�$��p:�s�j0Sjْ�Uamrejm�B!q)���x��V�3]���Պ
�T�U�m�.q�B�hVؠ��%6�35͋�4�6��جU�9Jkk�,�b�U�s-�&��)L<��
�e��j0��񁙓b�ͭ�iD*at���.���Hr'�O��C	� M�$>	 B@��U�kW�-2;�aA�h.Ғ�8Q�*Yr��śQ�M��� `Ku�D��ˊ�^j��ȎA��J�lT����ˣ0亇��p��u�G��mp�K�w,��	��/�}������U�V =�"-�7)�6�)px67 �� *[4<��p�^X��t�H���CD�(��d��� }WY�}�l��*�����⍽a ���"���/[2���i�Wn�ڇ�95��7a�@��ӠK�v��L�[����gZm�B,�͝��ߺ����m^y��������WZћ���)�G�q׀Fqq3Nl�;[P$u�܆s����'Z�/��N�/*���njl0Ќ� �x�ng�腑�(�D:�y�!�{XX�y��ιu�qMf��� uN�?�0�v�ݓ�i�IP�{s���M!XV���ZaRT�����t�[8�Z��q�sI�q0�*��u$�+
������T�
���ϻa�4¡�H&!����8�HV~��O�8f:�au�i�oY���
��X_=��l8��T�s{�M[�L�pt�Z�0]F��6)��)4���w�u�<IP�+>�����aX_;s���0���oW4���'wD|�o]m����æ��Z0ѫva��a�~�]Ì+
°��|�a�+
���ٮ��°�>���8¤����uiu�\���<洖�X�CL*J���s���M!XV{��ZaRT+���CL*J��wz�ĕ
��ߞ�kg]���C��һ0�*��>��
��|����i?I 䄦�i�ﻛ���
��X}�g���q
³���Km�:�s�oZ�\�evN!��	"ÿ~��q%B��=Ϝ���i%B���}�a�%C�{���V���&gZ�]�a��7��fo5��V�a|�����°�lo�XX�d�qb�v��P�1�a�v!�
'y������N0ĕ
���w[�V%B��ϻC�4³�~�L��k�gk��g{���۰���%��ҹ���<��
°��|v�aXV���f��c
����w�P�J�aXy����T�>��A�t��q����1�xk.��6¤�y�w��8��$�iaX_~���T�
�����d�¤�y�n��I�Vx|t��sW6q�7���Y�ֶaRT+�>��
����l��Ę��&0�����08¤�V��5�0����=4�T͜a����n�ۛ0�+
��������aXy��>�0�
°���Ohq�0�y���9���e.)�T�̙ha�sJݦ�	��\�@(Ptҟ������T�6!M1��j�ㄴ���cA��8��Wb��IG<nm&��@8�69�g@�MeFl�늖!v7.n
a��V�l�`��¼h+�X��W�Y���8���rNO��9�'�����5�q�aY�~�kQ��n�0���3fl�Cl*J��v��P�J�aI��9�r<�yN���`Յ�̮e����)��bnfByϟ�߷��%B����vN!�%C���=�Ę�c�o����u��9��x���3�A�bkf�U��q�n�T�
�����'�
����w��ĕ
°�>��XaRT+q��ݰ�aY�{ۻ���k.���+\浬�8��+��w���aX_>�k�q�0�+>��6���aX_;�u�q�aYߏ�u��n7gf�sy��k36a��a�~ޞ��aXV{����V�a~��ݓ�i�IP�߻ͨq%B��}�ꎴ�������mmѫ��
��X{����CL*J���z{C�1
°�{�wxaRV~a���k�!�+?w��4�f�8�kn�U��tkp�J�aX_;�wl�^B�B����<��f#0:1iYRf7r؈�8����w�>��i�IP��l����aXy�ĕ
����[nk������U
3�;�VQ��#3�m�J�١��n��h�Xi.�ҷ��.2���\㍀���[h��ukXsk4������''9��Ţ[�4��v��E�8���<aĕ
��{�=��¤�y��sp�
°�>���w���aXy߷��CVt�;C1�͜ay��u�p���V�{��8�T����mC�+
°���wt8°�+�w['�@!��߻m�v��7[8Ú�5o5�f�a�°�=�Ft�C�4�aX^��wxaRT+=���CT�3�;�I�+;�w3�7Y��]�aͺ�����Ì*J�a�~�ݓ�c
��|����i
°�{�wt8¤�Vw��ÈV�����֌�����ܶ�MÉ4�aX_>��u���Y��X�y�W��8�l͕�<m��*F5vZP�6�7;��i���a��:wp�0�+��w[�V�}�[�5�]kg]���ɑˍX���e���6�tkIva�+
������i�aX_���naXV���z{C�1�aX_=��hq&���ޝ��V���޹��K�:�Ì*J�a�~;�d��X~���/�ta��Ͻ�$�IĹ	�!�"d���4Mj���`B��Og�<IP���׈q&!XV�s����%B�������1�g��>���5��5���p�kp�M�XV�s���*J�a�oOl8�3��&$�=ÿ�nI�+
�����o�*J����q�eѳ�35�fq���Èc
°�{s���0�+�~�0�+
���w�P�
°�/��5�8�Vv�N���F���\F�4��V�a��ޞ���p��t�� JD���j�Lw*�(�Ѷ�v՝��ޛ��aԚB��/~��xaRT+;���CV{}�;�Eֵss�s��º�wZ��	nV��hl�	�<I�+
���;��q�IP�<��;�qaRT/���p�M!XV�s���*J�ݿ=�)��a���o5�����8�aRT/��;�q&!XV��]�$�*���z{C�1%B��:��hq��V}z?u��c�w8������Ì+
°������
°�<����8�؁� 2d�H���H} �Ѷas��w$��a���Ì1�g��]^�I�uw8��˛�k-�ka�a_�C{���`q�aXV�w��d��aX_=�k�q&!XV��u0����-��j�q���s���%B��:�׳�'%'(�y�WVjg0֓eT�e]fT�{½l�Yt%�)���n~�CĚB��<�پ�8¤�Vg����6³��*������.s�)׳0"͊XJU�qL�f��]l8��V���7ևT�
�����Èi�IP��}݇�� ��hV�~���aRT�����\�8�y�f�v�[4�nC�*J��ﳻ��!!CL�{�چ�
C����h�,<�����³�c�G.�ӭ�a��MWZsN���aXy����6°�/~���m��1�0��s�aRT+�o��'�
Ξ���n�[��5�g9�c��l8��V�������
��X_=�wd�¤�_>�5�8��vHf�<s�y5���n�Z��V�[��W9L�\f�*͂k�/3qiV��`�f3��$Eɡ�撄�C)-`G<�J5���Ȑ5�kh�qp\�X-ܧ.6�nUuȪ#��\C��
CjD�5���9Ÿ����؍[7�j$����y�9��0���!�%G���˝պu��7�\�|wu��8�T��o��8�$�%'h����0�їe��x��mZ�&��&�U���o����IP�/�\�l8��T�����a��w���
\ֲ��ޝ�I�%��nűf�6�L�p���
°�/�\�hq��V���v�i�aX}����aXV��޻����o!y���5T��N�/"��g5�aĜB��=���aRT+������4¤�_{s���M!XV���ZaRT��w�z��8�y��n.��4¤�^��wp�M�XV�پ�8¤�V�nw�CL*J����w$����sx��kgkZ����/.É+
�a|�������X_;����¤�{���q�aXVϾ�sXaXV}�S]W5�vq����̚���Èq�aX{��;�xNbJrRy��DƸ�9�"J�W��E(�u��
w�|�s���$�V�{u{C�4°�>����8°���v�c�6q��#�(҇i�2SJ���F����-�r���-Xk-�,KWihV75����`��]�ܵ���Iv�K�ҡXm7@eA���At�t�l8J]�4��f]�s�%9+
��۝�C�4�aXy��z���aX_=���8°�+��gvN!�+;�׹�̸\���7�n��z�$�V�s���T�
����vN!�%C߾ޞ��LB��/����I���rr$�g�����3���/#���.�m�Èq�IP�߶~�8��+�����*J�a|��ݰ�aRT<�뾻�T+>/����Z�gk��zշ�fl8°�+��f��c
°�w�P�
°�;�}ۛ�V�a}��ݡ�aY�s�޺�Z��z���.Ì1�aX_=���8�Y��Y�琳����q5E&5]P٭���b�3�������aRT;����I�V�����*J�>�W7uZ�goz��n�l�6K�ҹ�XD2M�[�q0�*}�޻hq%B��/����T�
���ϻa�4¤�}���q%B�߲߰�s��gg9�sfh�usa�%B���s��q� 8�!
�2B�c"F� B�D�" (D��d@i ��A��2��,bH�Ĥ$!$����J�����I�V���0�+
���n���Ñ9)��~���q��ɺ����:͇V�a{�{�Ì+
°�v�{C�4°�<��z���aX_=���8¤��q:ޮi��7�Uy�e�8��T����ڇT+
�������
��X_~�wd�aRT<����$�+=���3K�j��0��<�w��ka�%B��>��vÈk�Y����'>|��|֡L��6�Z!���R���_'~���u%B��/{�wxaRT+��>��J���ץ]`�q۾~��l���Q��C(&�.�5�Z���*%B��kp�
°�/��{�0�+
�Ͼ�6���aXw�|��I�+=�z�u�un�0�r�s���.Ì6��Xy����a�+
���}��q�aXVg�{�'�+
��{�mC�?I ��t�������{�ݧ�:��Ó�r�V����0�+
�οo]�8±�N�і�)�{$`ă3�y���,"f��(%��A��,�P� ���L#,u��l��IL"R4ig�l8G�#�FX�Q�@b��A0�ܘ��#2"CԬ�$ ��!.̉�a`d�A$A �{s���4`aac�u���h$�iF��:]�q*�\bmq�5X-+���C&������n���c�01�cG&1�c���1�k���ҵuS)�v�V��kZ���1��c�0�q��ֵ��Ae�f���h��&�f�Gf��\��6Vb̙[v���躑,��F��M�JU 6�6bsL�H�l2�cWD-r�m.afP*��e�F�b�5&i��5u-��qjf-pXYB�G����Q0�f�58�D�nlkEtjJZ���l�3�8/
�3t�d�գ�� ����U�F�NP��&��W!��c\�th&ˣW7:�M+YCaIn��ln��S"ۑ�XNjbW�x�T&RbT��L�M4	p��ܮ�^ ̬��7!�!��!�k]����"��S�F�K�K� iv�qai��Qv�5�.�rFaGI�c��ᘖ]�gP�-\V����k*h�ER�V��Z�pʣ�`�;J�54 lvn,]m�7#E�jٲ��Z�ip�\+�붫��nȨ�v�8���K;R�����L�%x�!�-6�l�.kRb���a�F�6j��vCjak�Tڑۘ�bZ��B[4�jU�պ<��f�u`�@n� fˢ�b(�S%������KYc(gX��P�%�����2�Ի.�LM
�ˣ��ka0f��
�|�9�?���r�B OhCd섒{	&�n�� 2`f���I�ěB��s�I�+
�������
��~�Ku�-\��0���f���vN!�*J�~�γ�8�HV������*J�a�l���1�IP�{{�É4�g}0�Q�U��0��5�˭��ka�%B�����Xq
¤/|���fb\��h7dҲ�mQ�l1V2錕������y?�
°�}�wxaRT+�~޻hq�aY�ޮ�k��0�r��st֌�nG��v`�c2��QbT��0�+�w[�V�a�ޞ��aXV�_:���0�+�{�ny)�N}����G�Ñ�{���S=��aRT/����8�HV���u{�0�*����6N!XT�߾�u$�+;}�^�7Y�sg]s7��w��l8¤�V|���'�*J����w$��a|�>��8¤�V{������~�ou[�[�B���uu�p�N!XV��{�0�*���z{C�1�aX_=��hq��VO�����>P`���3���g3V�]V�j��E��k��5�<VU��ek�� 8��������&�j�u�O�n,��la��8<�5��؄-q�J�X9	Mj��Z*d�;�+vCQ��	]B
2�L�K�����Kq���嫝�!�a����70�+=����B͖��M��:��U���
���]C�1�aQ�i��%.�
ij�0x���n3�����գ��>���>aXV��=�]��V%B�۟v�i
��{�3/Md���:�xv�`��Z0��)�S.a��ֱ��q�IP�<��;�qaRT;��ӝ��M!XV��{�0�*����=��³�}�Gz5u�78�f��f���I�+
�������HFbLB���߹���*J�����É1
��}��wt8°��׻��f�q���9�Zk�h�q�aXV���l8��V���8�HV���z{C�1%B���oNw�4³��5�sU��C|�ܙyuG[�V�a�o���+
°�{s���M!XVg\�Za��
����V��L��E��!y��Ѫ��m�aX_��5�8�V9�q�"�����f�lu�6������4kE�����J0�*�����CL*J��۟v�i
����s0˚���g��c#"�BT�2�ed����@@���1"D�F#�	H1Y��  �D�Z���� �A"p���&�j+1�ͫ/�ܵ���`˱�����0��IcX���َ���c, R���IQ�a0�д����K�;$�I��''o{څ�vyDv\��]s�鯡�
��Xw�=�8��T��~�p8�hV�����C�*J�a|��ݰ�aY�s�;�u������3uᦻ�q
°���\�
��X_��5�CT���gw0��a��~�naXVt�_����vq����y�o͇m�aX_=��hq��V������V�a�~ޛ�0�
°�o��m
����r�:��0��Jl�%vaRT+�׽�8��T�3�;҇i
°���\�
��X^��wd�³�=�p�j��={n��C�����������l�^B�B�祾qc���՘Q��e��
�Z��Z��<��ݰ�0�*ϯ{�q&��+=�o�0�*y�|ff[�6q�k�������n��Ŧ��S%"a��Èc
°�o��m�aXy���q�aXVϮw�~B>0�
°�?9��0�
��w_�s�vq�o{��9��aXV��f���`$$��@B2B0���}$��q%C��\C�1
°��?k���%B��{~���?H7a���1���7s�o��o.��YvI�+
�߿f�48¤�V{�'�%B����8�hV�����C�*J�W����֮l��\�sf]�[��
� I�����q&��*����0�*��k����aX{�}u�CVv�~�5n�go\xsC�e֮�ĕ
°�}󿬞^F�B˷|AJ�ʵ5j\Ҕ���s.p�x����˹�=������T�����8°�+���C�+
ϯ��k]f][��'|-�K/��pG0��ܬ���Z˚͇q
°�߷��8�T+���0�*J���>�g� |a��a߻�?�q�0���u���K�Wgo\�xfj�q�IP�=Ͼ��8�0�*wO�]C�1
°�}���aRT+���C����~�ц�涻��Ⱦwx��3{'�q��a��0�*��۟vÈi��$!�@��M!���É1
°��;��q�IS���׺��8��o���f�Èq�$a�w����q&!XV���;�V�a�{��P�aP�G}ݽ���c
Ν?��0�k���F�kp�
°�/������Ȝ��:�o"��7�lG#v�xhi��p�]�����{����aXV{��C�*J�a|���'�
ϽϺ-�:��!��]��p{	e+u9�����9%�u\�É1
°��;��q�IP�<οt�8��T���z{C�1
°�f���
��o���[u�n�0�o�\֓F�[��
����~��8��@4�0�/�~����
��X_~���CL*J��wgw0���~�ou[�[8��E�㫭Wp�
°�/���hq��V������c
°�������aXy�s�8�L+<���햖�og�&ώ��d���%!Xw߳}hq�IP�>�_��q0�*��뮡Ę�CS�2"$A�`E H�D�BM���E$�upẃ�9ɝ��l��٫��n���i�Ա҂�hj� ��E�͂X�^2٦����Y�٥KY�1��6��+)�*4�%�(G\��-y�vq�و���jB&�]��&�6��R\��e��q��+5q62�i�� ���l=������
��ǣ�cs�avq�f���汻'�
����ޞ��LB�����Ǚr�ĵ�+��_Ώm�v:g�H�&�5ˬ���nw�C�%B��v�ݰ�aRT/����8����Q���g��s^�lC�"�ËIk���˚��͇T�
���w��B��*���8�0�+����IP�+s�>�0�J�t���LӚ���ͺs-��0�
��|���p�
°�/�g{�0�+
�ϻ�=�Ę�aX{߮���bJ�|u�Q�U�8�{�������IP�{�k�q�0�+�����+
°�;޹�q�aXV{���CV}��2��s�s{ޭ���]fl8��+s�����
��X}��CT��f��b�a�����/!g?~?3�#vyy6����:mÈc
���~�;�q&!XTrk�,iମ�0��5�n�2)�&�U��w�|����O/!g!x^��k�8�0�*����8����?͆vs���v|4�cK(+���h"�ͥ5�-д�K��Mm������ ����K�K ۉ�[��V)&vF��əMMZ�Q-�Y\K��83���F�,��k�5h�Ѧ��q�aXV�����c
°�߷��8�V�����Ì+
°��\�hq��V{~~�vۭWgk��k9���sa�aXV߻�naXV�����'�%C��w��8��+�s���*J��>�f�:��0�k��p֋�qaRT/}�5�8��+3����8¤�V����Èc
���~��É1
������X�[8�7�އ�ݹnÌ*J�a���q0�*Ͼ��I�V����w���aXy�w��8�V>{��̽ҹ��9��k�0ѻ��c
°�w��p�
°���*j�˭f��D�c�
1*�.0WG�j��!Ӹ���Z%���	��nMh�0��a�w�sp�
��{�v1��g�&�|�xUB�Y�sƳ5��ab��Z�s�LrRr�{�S�É1
°�=��XaRT+���v�	�6¤�{��O�I�V{��]Q���1�]W��݇T�
��{�=��ܒ�Є��a�����I�V����w��%B��{�k�8�0������en���2�h�u�6N0��a���É*�a�~ޞ��g�Fb��߷��0�%C����p�
³��[zV�vq���<�]k3a��aXy����!�+
����w0�J�a��]Ì+
���~��P�aY��>���og�'_5���r�OJrS�����=�𒜔�/|Z9ll4]�r�C�������5�j�.���}�5�8�V�}���$�+
�߾����%O�����&f�vyy;��A�f��3ڨl��WY�c���qaRT=�\��8�HV�Oo��T�
�Ͼ�݇ ~�� ��~�6�Y����uqn�%������p��Ͻ�����IP�{~��ĚB��/����T�
��߳]a�1�g}3�%�WK��.o��j�y�a�aXV����aXV���z{C�1�pH�A��a	H	'd�a�ι�(q��V��{�����g��Mz.�0��5u�72��aRT/�����M�XVw��ZaRT+z���'�Ђb���C�4�g�c�×X��0�����[���[0�*��gvN!�*J��k�y�-�\�5�.�Yy��*Z���ҙMc�����z��+�~�wC�*J�a�{�=��³��;U����z^�`	�妧.v̈́�.\5S4�kp�M�XV�w���
��Xy߷��8�V���w�a��a��]Ì+
��Lnw-ӭ�a���3u޵��c
°�v�ݡ�aXV����8°�+�~��CT�=�]tC�1
Ο}��&Qs{<9<^���V=�Ò�������l���1�IP�=s���M'� ��tϳ��`q�IP�=�v~�8�0��祷Gq�h��!����k�I�+
��{��C�*J�a�_���CT��o��8�HT:~�� PD`�󏞹�LmZ��kS]�끨��1iq5�ɀ%v�íVa�6d#h�h����9��J�Ћ�-�����ׄ8$Wb�a���
A]2[s,D�T��6�u�7r���:Uګ���`�u�Z��wYG �x.Z7l��J��o�䓓�y=�����J§�w�Gx9�˳�39����-��8�i*��뮺!�§�#��_�t�ep��t�1Ao0Y\l��J�w�}���O㒰�+��u�0�+
���ϻa�My����cY������Zx�U/�A16�t),]p����Y�,+
��~��Ì1�IP�����6°�<����8°�+{��]��V�|u��sE.�0��s3�unÌ8°�/���hq��V��ߵ���
��X{���8�0�*߾�u$�+=;���+vq�9�i�o2��T�
�����'�
���9���M!XV{�o�0�*���w�!����6�\5���CZ�י�u�5�q&!XV���C�*J�a|��ݰ�aRT/���p�0�~������Ì+
Ͽ�?k)�ffkgf��I���l8Ì+
���ٮ�yy�^B�� j7�M�K^6�f�3B�v6�P�\�f���7XV�a�z�ݡ�aXV���$��ߗ�;m֫��9�͞�y�`��~;)��",�����c�@H0H�DbXn	!#z�s�v�4RI�)���H>��"*�ɨd���"5�K�O4HȑTFDF	�l����� I�"0dF�FX)!�M�Æ���(D`e���@O}��H�1�����#�8hT%b�������L����b��x�;����l$f4��tm
����u�E�Y��UPUUVڪ�EU[m��m��q�*�mUAUT-շ,�֮jLiv�Iy��r�0�cSSBǙ�6kb�MM@�cM�(7,��\�!v1���/2��Q !
iC$f����)n4+*1�0�#�:6�E,�+U�LM�n�v�%�ҭ�IhJ�4L��A2Gr�+2n1m.
c�vv��;+v�5a��ce�TC!b�-A�i��٪GF��.K��+���앗3V�))IB�6�\8�	�n��$���[��1��]��,��6D��[���nkʉ���WK�[�f�@�ۥ����{��m�t��]t&����r9B������̶b�N+K,t3��]l t�8M�[,5�2��HO!$dܐ!�t�)7$P�z@��p�$!�$��$��`>��;�J�4S$�XbƵk��]��BBݝ@�&�Q�l�SF˂�0��t&5֚��h���c�j��F��sVթ$�{��w\��X�d��FW��*���'�*J�a{�����4¤�y����I�V�������%B��v�ݜ�9)���;�ld����%�Afw$��a�~���%B��߶k�!�*J��ﳻ�b�a߾�!�%N�����9Mf�0�ۛ��[�.��4°�=>���a��a��o����aX_=��hq��V���z{C�1�c�~\��^��8Úw�8hְ�8°�+�n}�a��a|��ݡĚB��;���8¤�V{ݝ6N!�+;ߵԮf]L��!�sy�h֍��q&��+}����B�B�'�ig��XM���Pq*y�a3]3e�
�Fw�~��vO��
����wp�M!XV}�o�0�*y����;�vq��71��[;�������m�A����4¤�y���p�LB��<���
IXT+�n}�!��
���ϻC�4³�������q��慴�8°�+=�|w08��@�1�a}�ٮ��°�=����8��XV�}�a�	 n����/�n�s�a�o8ۼ�k6a��a�{����
°�/���l�B��+3��u$�+
�ϻw��aXV}}��u�����q�j浸q�IP�/�߻�q0�*��붇T+
��u��0�+?B8�>�s���1�g~�S�юh˹�.s���oE��q%B��=�s���*J�L)�d�*T�6��M@[�r�]�[Q���}���'��^A%C���É1
°�{�wxaRR}�-g�1��<9*�_,�;ԕ�T1�a�3A�Ʃ��O	:rRr��ݻ�q%B��/�}�naXV��۟v�i�aXw߷��aXVw�:奧M.�0��|�k49�q�aXV�n}�a��a��6���aX}����q�IP�>;�����w�O��Wnf�Sz2㺯�w���/�߷r��2>@�Ld��H�K
X�$	 ��}��f�}�\�:�5=6��z,r�:@>��U ;ˬ���f@�nT��ܧI����{�w��v*ۦh�����n�̠\�vb�F�&�޽��;ָ˪��c|�9�ܝ�%#47jdYeZ!-LC�jn }z��[4>�� ���T�]uk�i��$��d�[�˹�h}�yb>��u7�)�66� �uV �[� ׫��\�+�{�4���V�l�`}�Y��q�\�9�Yl��J�����v/n'�t��[R]�]�v!41r+6\�Wff#��mL�BZX��P¤ř�↰�fܲŖ�#�H�5�%],�Y��NfX���F�7j�Bƀ&�f��3Wh��F��ڛW/R�T����*J��$�"�؎���5��v�Y�$$�����f׾�}�4��L�!'����,A��i�i���<����[
�,�Zi���w,�}�W��Um��ܙ�~&�̲�˿�9'�P:,ren4�060n��
'��߿������n[�@���x;�3U`(�f�oS�r�lз6� �������[��Ѧ���Mbz�zۓ {�����WHj{��Iǯ&=Y �\ޯ,A�ųC�[v�ͩ&�"��Ԗ���߻�#:N����-��`��#��l����<���o@�� �v�}ݻwt�ȵ�鿷Jt\�g�E4�.6Jv��[qJa]�ܸ���\�V�ԛ\�l0�q2Ćf��%��X�n����`��-p�nI�$e؂�֥Ќ.R�t.�%��{���<�,Yrs�[	/�s�Km��S�R2��"׫^��۰�<��.�C��v�jB�H�͛�7n5 =� /Z�ut�}���4��Di����bF����W� >-��b��^��	|��;����1�^�w����\�����۠;�RK�.�6��aٴ̸�[3�"ӯe��� >�m��z�M�NM՛iQQк�R�7&X]uk��}���4���� ��c>)Qq	�R �u7�Hz�G�!+�!޼ː��r�YjçP�4jN7�V�i�����d?�C|�[rk͹32e�n�iK��Cx�����k�>�t��٥�b[�4�ơ�9����-� ��${���vlt��(9�,t���5%tسMG������{����Y�/b���Pa������@�w46б.�@���:��ˬ���� }��hr��2�70W����Z�[4>T�4/�����؋��`n�{�u!(�ɡ���j��=>�jC��;�!H���١ޮ�<[��Sf��3`�Õ-q�^t��١���i�:��g=�w:�3�~�}��x�w��.;B��coH���$�,4[�D}��w� �ِ��zߓ���J:�w�l��`���έ؅.�qއ��~:��rxfV�����ZXn����(�������о�t�yu����{��$ĚJ9��kR���U =�l��������κ��
����67j�Wf�(�	�孶sv�/f����|��~F)�����kW9��m�f.�Z�;eV�!�]1Bx¥��Z!͌	�cXͥDl�����eյ���l��B��WY��R�f�9���4rH�3\��Z`s���^(ZM�*i�Nf]��\��te�M#��X�W+r��$!{O~���&���1��&z��wݠ��]��n�&��L��9��Q�I�G����n|��T ���[�a�m;�ߧ9$�'�Z�x͒4�Y�P����>P?{�� ��K�C�<��k�{�3V�c#�d�-����H��p��b��d��n�N=�<f��u�z�����˪�4��sjDjDF4jKb�� �x�h_g:@�����kZ��nD���q��4<��ݝ��ܑ�Eo,�-�迻�[2Ρ�E�KMhߟ��� �V��^X�x�k^���q���G�b���X��Ʈ"h�9��c�T�1cx�KT��]��*��L��Y���:�T)��\��e87G4�☴(�3ĺo�����rHt����\��`jmk���͹��z��C�Y��� �x�4��KV�C6Fl&,�{��up�[4>�Y��j��^#ww^27�7'�4>�<���p�R��Y�>�j��q]0�I�`�� �x�4>� �������mX�n�A95���Y�o߿t=�o�t+�-�"]*R;s^-���5`M��}�ߟ�[�,@}��-Ԑ�Bl��害�m��-V��GGmVm��� ��ވ����x|@���4�u,N���{��$朜����K-�{+�rs2�����Z:RR��G�ZlD@{���.�`z̀�"��U���Y�f�6ם �V����z��⦥�PxD�-Ǭ����شׯO�"�nR�CJMs��H��[����e�ܺ��[�.{�?�%�ղ��.�wT�j�n��X�݀� �^� �ΐ�.�K���׏`�	%& �z����Y�u��>�<�.\.�6,p�Gl��s&��3-YȄ���v�.%������ai��X$AD�j�
; J�h"���0�S��$H������

2$��'�5��!�0M���8"$�u,+"j���	D$�g	��%ɧa0J$#����F��܍��	��@A��K ��\�f4C$��_91�&�����J)PȔ�d(�!cA(%�,˃26 �(�I��I)i �B$�`z0
a#���D%DI�K0c(2$ID4k��D3�Ny�c2C� �2� 2J!Fi*

�&��e�����@@E�1H��"�"�&5ZK���(dI��#6h�D�f"FY<�s.Oq�:Ƽ�V��ĘnTAL��X%�!��-�4!e���qx�bV�`-���ukZֵ�ֵ�kZkZ�:��Lc.������Tؘ��4�����cʀ��1�`c�1�3�Arc�K�mX�P�l%ei�e��ΛV��j�͖�04б�8���\�s��&���3�L؋�)E49�x���h�c���w5��ELY��E�i��F�)�7f�P�T��m�Rk�e�Q
;[
#,l]x�F��]��:+�2�5\�.�3�5���$�c<0K��6PԖRU�˫�d�,4v�����B�̥D�@�⵰چ-(�[*�sBTqmZZ�WP6H�tS*�m�o�5��XB�͖	0Y7
@Р�MV"h:�B����Z��B`ι�ƎR��.H�`�;$5���bR�.!(5�GX��p3�҃W(a���kv�M\5�����5X;Za��+�r�&5�3mJ��v��j�1m5X�A�ɲe���B�7V�j��ukZī��)�-�u幂��݃5��V�v��[�K��ԈF�6-׊�4�a�X��c�8�B�k����#�D�(�f͋�`ҭai�d6SK`��^V�ҕ��ɨ�n�-&.�1�Ԕ
8WVg 1�q+���b\�ە��gEf�ۀ+KF��l��3)K0[kv���˵X�h�Fh˘�Qҹ��Oa���$>�jBHs�B��� ��$d��j�Bo�g�����kjq��~t�Z��Ȗ�K^�.�@���>�yb��Y���UK�mȘ����Y�hP5;��z�9Ш�T��f�#�[w1�ƹ2�����>]n�;�́�~;O�mnH�e�tX��jM�B2Rf(������� �]f��.�OuTI4�r`�=��s��;�p�] �]f��w[��4Ȅ�<�޶d �ݶ >��u�2��M11��ֆ��f�����] �}����s��|��>W6�-�Ůrgj�W]+r�q�T�Ơ\���vm����l@�jB+��*�b�P����m2����`�"��LX�n��)U&�R�A�6U��Z�s[�B�LEÊP�0�͚�M�Tv�����*6i\J[3��s�rrN>�o���9�f�`(��2-z��+fڼѥ��Řْ�*@����6���e�y�������vX���fgqQ#���Us���h>��dn���]5tyQ��-|�U�� }�٠{ˬ����Ët�wRq6���s@�[}�� >�l��S���ͨmG"cŢ{��]�{���]�yu�{ݵ�Ks[�j�?n1湡�����,@S��>�:@�F��jj7ɺ��4<���ٺR6��E2�i5��EI��l����� M��~����������u�KV�C6k��߳���^λ�j�.i�T0��!� �e.�Xhܭ+t%�%S�	.tԫ�;vv��ٹ;�ݳ�Qt�2��J�7'9�M@؊��9c-h6�@�x�1�����`ge�w�X~�Q��R�g7v�B�!ȍ��4��{� ܺ��:��t��˧䴻��di������W���m�yu�P�V=M�j$҈�D�ΐ�la������T!<��)�wSzF_�>��KWf�B�P1����S%��7,jZ6��6�y�߾ߠz�9^V#��:�k#n6�G�\�&��X6k�u�AR��9�ܹ����w��6!|��ۓ7fZ�Ғ�M��X�e�3��u	Gf~���<�d�����z�@�(��$�SV�&�k#W���W����D&���܆wim�1��`�T�nB�Ǩ ܺ��yb�W �S���v��\��[��7wb�] 
c��6K���V��DیbA�<�m�m�����^� �X���p/#�\7^=��Df�M_����{�[�f�6؂0�W� ��H�.�@�ݶ#ܭ��(=�x�% �S���� ��� {ˬ�ǅ�Q�ֶ8���̈����sp�!D(S=�R�a���ÜM��9cs[L�1�� {��wW �^�a�!DC����3G����J��sfν-�>}�o:ӵ�F:j`㖚� ka�a).���-��^A��v {�\Z�=Bi)$�P,6����v	`���A�� �z݀{����i}�u��n��H�S��� ���������i�uU�'�qűa�{ ָz��{�X���v�qv,��Q�m�5kr������޿����f��6�٬YS]����]���L�,��%pʪ&�Q��l3(f!�B����;z]�,�Y� �&m,L�6�e&B���.!)%���K��e�4�D*�v��k͈�db9̷WM �M��J�.��\����l%.e+�]r�A��'$��IȈ���m�s���uR�K���͢]U�}���p=zl��[�CqS��6��ʸ`�]+o�~�������<�-��I��f�u���vrda�T�l���@�w]�u�^�|�]�J+KZ�kؖ����`z��}����hr�+ݗk�F��rd��G�^�=������/u���lG���j�L�w7vJ��nm�����l�ܭ z���up:��n銆lsRN1�{��������P�c�,�"�	��4�W2�KpZ�����^�,A��#����7G�8�����:�����l�Z�Eb�X!ͨj-&���QtvH�4Ғ��X؜�Q
B�q�Rf�Z$�[rj�Lj��h֓@�0-��p�ͨʑ��J�+YkB��������{iby�v_�j���"RA<�{��ָ{�X��V�;�Zf��Q&�Q��<�ʝf�������X'�U�73.�\��>�o���m-�8������݋���7sCcH"�o�wn�۵5k��]�m(��2�\��響=��ws�|��4�wU�=��no�	]XF��GR��4q�>W��>����W ���o��Sf�V�ޮ[ށ��~z�NI'��9'�	B�Tv�K-��{�A�v���qL�1+��Ģ�z����Y�}mp��b�����G��H�	nL�[aBP��km�޽ې3�ʰ;���g�G~��^7D��J@������fN������R2�vM*XkX9V���l�gO��}?�C�����up=���`޽�kV鈁�m�f�7gF�&�:[����wW �W� �x�4���mk[&�J�P�yb��{�f@/����e�f�M���#N@>����y�z���
�0�@`0$� BH��5��Ǜ���~���~����-�Tѽz����h�Hg;XXj���f����5,tۻ��{�����_�����:��l�Ѓ�kZ�+#��M5Lغ����n�j�h}w�����x�{��u:��k͌��[,#FnROl�z�؃׬���Y�{��K��i����9��� =��hw�XX��,�N��%O���ْj���{3V��W�@=�^�^�2��5��z��`��u������گ�_~�9 9R���ADV�@�xcu2Db!�')�rY%�c���jʡ0Ba�sU�岴qV.�e��G3&�GV-�)�5�T��f5����
�ь5���㱛˭�B,l��a�-��d�ш��1��:��U���^&�)x�M��R!+SV�:�l\��2#���I��2B����{���1HL�uW7�wA\t/��wf�&�m��1
%6�b�M�-��nƭֲ}ˬ���H����r�Z�k��#L[�Ç���u���O&�F�̀|��h�lо�H�v��nl�я4#B١�s��������K�4���z�[I��)��K4�{۝f���b�f@>^�}�~|��+=e�wP4c��_�I�"{ܽ,�ݫ��yl؄�"�Z�g5n�hNj\ܖ�UЋ�>�̹�Gd����j[Y�U���f9DiM0[�7ﭿ��{���{z#��T�2���I	I'�d��$��䐐$��HHI,��$����$����$��HHI?ؐ�$��HHI��	I'����$��d��$��B@�Id��$����$����$����$����$����$����$��! I$�HHI?�b��L��7z�\ �|� � ����� ������ ��׼       >
ި�[}�.�<nw��׮g��j����pVr���4�ْ�,��64�١V���A�$+�v�ڇp���Sli�S6]�\ ��]c��^���kl�l֪����G�;�B��{m���=�l	����o   @ ����U*���U4 hɠ @�  )�L��*Bz��� A����h��UD$� �     ��SBT�hɁFL 	� �F�	�J�P�2 �d��i�A@��Di�І�z��S�L��4�L��顤��G���" ��I�V
=}��Py�� �Q ��6C������8G�����?�����P�Ŏ��Vxy�5�;�ۯ���7��F�sٞe�s�}3�J���bc��
5��ߤstq�oӖE Qި[����ӊ�tX��M˥J�E�A1�PKŹ�N=���o�������ٴ�{m�����jv��=Ge�N>M���<ꪊ�<�U��C:�:(�
���6�5��B��d��[H�b�@�PJh���^��3��
�r=m�.ԑ�j��r���V�1�ծM�@!F],h�X�X�JSx���U��H��|]�`��B�Hx��j�J�b�Q�i��S[�؅;����*Q)-�)1
��U��`c��6i!IHPE�700��H]#Q�cF$�ňA]\`��
	Y������ļ�]�a�+		*�!D�@\JqD
���v�QkX��좭}i)�`#E�P؄3%�B0�#;1��aV��(�J��Q#6����@#a�,X�.�1)H��)HD0
 ��� �@�̌ ����	$�I-"E���d���$V��E��XB,	R���u��7 d;H�&R�F�"B�`���M4l�
�1��|tB	�!!���1�0�[K5V.,\�tޚF��n��ꯛ�3�:����s�>����_��YB���V����{��%��p�\.a�a�a�a�a�j����a�a�a�a�a�a�a�a�a�a�a�ڣa���a�a�a�a�a�a�a��w���a�a�m�6ڣa�a�a�a�a�a�a�a�a�a�a�m�6ڣa�a�a�a�a�a�a�a�a�a�a�j��ڣa�a�a�a�a�a�a�a�a�a�a�j����a�a�a�a�a�a�a�a�a�a������6�mQ��0�0�0�0�0�0�0�0�0�0��F�mQ��0�0�0�0�0�0�0�0�0�0��F�Tl0�0�0�0�0�0�0�0�0�0�0��F�Tl0�0�0�0�0�0�0�0��a�a�a�a�a�a�c��9�p�nuxo��Pt��8h�L}�֞/�8�s�t=���M/��fo`cF�6&j��*qK�ӥ�S�$�stN�{U��u�wQ'w�K����<sN={�YSkf�IV�o��@m�ӈG"�֏fn5��y�T�ݘOw�#Bָ\!�s�'�P��&ofnc����;&s���Ӭ�3�kq&�,6Q��8���l���p�w�q�=��4r=�"ܮ�<\ �C!p����ɜyL�2�Ҋ����
$�L'�kZ[�T%N�)bB6-�;zD�;���Y����=����=Ǻb�C!p�w�q����� ���x�ڻ��Q���^�z��40�0�u���wt��tI$�)B�$���<H�.!�l�C�3Sm�m�x�����Y�'|����p�\.��� ��H�;������ʚ�%�rG��\�=&���\$�\4�k�q�=���2�tP�$�c�Iot�LFZ��}���p�7K	 ����#�$���n���=��}������IH�4I$nl�{����1]v�$���4�qYÏP
ʍ)��3_��E#!��ޑ�\q
��P�;{��  6�__�=07��������pQ��$'47�.����`e-��Ieq������>��E�@�R�:�D�i5�wq\�%>*bIk��l�wt��w ���.�|v�9kufVE���+�%��v�KY�8�ח���t|��uq��\s+1�&qe��0<�3?K빙��?,��$�s��i`JЦ��q6��9^n����a��Ea�]�.�� o���F2�-v�9����xѷ?������U���(�� �� *�E}i���������s`�QU:�k���uy�?_ì�'��Z{T�!䭅�)�*�#�0��hE�t��n�SAu ����3�� R�����WI �H@�6dbC(K�n�@��@
@�&P04!�h���,�v ��\$@�.��.���( �HHI? 8
f�7M�R�E����}Z5UZ5UV�U[UUmUU�UV�UZ5UZ5UV�UU��V^�tW[Qa���u �$�(�Q�96LVu�*����N�Jo}}�rn-q�"i6�p����ͯk�����kvK�Ì�ݮ�������/f����OY}�E-D��}��i0b� {�D"s��{�6���9���b�����k���)�v|�
�����{{�@�h�;r�pc	�&L��}ŗ�zpt6���-qz�@�Z�y��Wb�d���wj�������aD��T�l2s���Z"��0�8H#&cn�C�+g�G$����ɋ2�{� G�I���6��KJR*��IA�FS\T��R�Fw���s��������T���7e���\�{�~$�~���$����nV���cs3�f
�1�2*�@S�(����Y��/[S�}#ΐ(�ړ=�ϗh�Bx��  B`��
n�J�`˺��=8:GV������<�A��M���>˙wa�r��pJ.*���Nt_�%H}������쏦I��I��b�۵�qąKPv�\U�'���^�n������Ry����b��6��99���4�=M�R%�锝N���P�Y�����N�BZBZ[P�X�\��aeR�ᛶuwכ�^��nf^r���37jb�ٙ����ع�֤�V���K���V�J����}��(��QAwGH���2U�a�x�k4�n��9��9����o���ٿ���G�h�������#�$�!��,��4�Ls���٫�� ����"""" ����"""#h�����""" ����"""" ����"""""D��9y�9�����r���x���a�u%qmEqG"��8��ګ�G�5q�M٭�����b��H�P��%IP
jj��4�&�m�rкT�U83m��8�ړ&��r�ff/�@ު�wb�`��d����@��!z�9&���W��|�3�3��C��͞�-��PЉQ�O�ZZֵ��[�ҿ?  `���PX�h p���7�EH�{7�Rz��ЊQ�ffu`���3'����춐���������HQ7U�2�z�7�g}䯖+���Dߛ���d�~fw'�ݿ���1UU=c�+�����>
�>K\�������b�J�7ͯ�`U=��*�B�iQ�,���'��P[[]8��ྐྵ���UW�[��J�'~Z�0�a��"�����~�۪/t�_O{<�O�LL��ɯ�w&�����i4��j�#�ވ����!6���nj(�Ě/}gX @�1~8�܅Sqo�p8EW7㖯m�|�!�yr�~Vȣ������z���=3�S$�S$�r��3���o��k�k���9�����328]@��mz7��!_}Uù>u]���^�S�I�}פl���b�wL����fg�w��W�{L��T#C��Y�4	=m�U��*��ĚY��#��io�SNb�4����]�oS�����~��a>t�< ���旻=���jK�k}�ԕҵ]��}Z�?UI�{U>[�����S5U�������@>M��|���3&s�Cm�Fɲ;V��Y�F�7���@�E�����Ɔ���W׉���RO.{�u���"!L�Oɯ�޹��P@y���z�ﮧ��W6��5�����u�o��t��m��{��I���Ez)���z�F�Y	AHI-i����x<�j����z��Ͼ������H9�#\������t�ް^�<�b����`�X*�W^��t�<���M�ѱ��t�����^���C�		!p	��0���ܚ*�� �+�xw��s��Y�kk�Uz���ڪ�j������j�������ڪ��[a�ҥ��q:�a��]����Nq��{��(��:��r��E���	��4�\9�����?0��W���뚪��ݵ48A^^�?���+t)-?E�Ef���`�)��g��-a�5�z��.>�?��Cη$�Q�����̕�j�cY�w��\�]r�_�bV�^8Z/TWʥ਱`�[���c]�k�[k�f(5�w�E�R8^��i�7d�0�/E�C�X���`��`�[�u�-<*#ZO���S��l�3��c�Qeח}v/��1)'�Q֠�`�rn� �I<�<�f����±��8�`�x+,��}Լy�w��Џ�S1L�1L�Fݜ�yv�x֢�F%{��sw9�_���d��o��p�s}b�(��^<*�b���C�ذTYu�{������X�d,�<����"�M>���/������K)P�τ��"#|��픠����!{�=`�)��g��`��`�^��yJ����V+VԖ5��(y5cG3[k��3�:��Zl�^O
�u�T,Ԓ/!�W�~��x�^���&��`��o�}�.��z���ͪ��57���1�<,��z�����_FL\�X)&�>jtXY�k�v/��b�麉�t��(�)Lǻ]�����i�S�+"&׎���2�~d�-����7�ʥ���s�e<>+!�鏽55�S$�S;m[n�wR�n������-{˼�k��I�v&��W�ks2��JՍV�Up��3�^އ�r�*,X)$X+ϧzbV�ñt�*���o�"`q?C���t]�s�q77��e-�%����!%�j�mҲ�hSz�X�:k���*x+,X+?:���+�±]�~��j�cX���N�d]z��$#<")�k)p���M�V5vk�\��e��z�jRKST�^�����v/{Ӽb��k��m��_H��� �0#���~=�7�R6���^�}1r�`�x*�W\��c�?>���!$�Z[ֻ�.դ��ޖ�ݿ)JJDDDm�DDDDDDD@ DDDDDDDF��t��+:6��^�6�e�61	yH�г��f!��t&�%�����(��l3nj�r<�b�z�������Uz����paC��4.<��"v�g��T-,�~پ����z�z��Ǭۣ��ˬn���ɸ�uR��ZxV9�Sb�E�����z�x�^�5d&��hb�y�������ߤ��f*)��I��еƞΜW]vj���S�e�Q�/4�����'�X����ƀ��[�^</�*�K$�b���LJ�C��V.��P<B�����D��r��2���\��y�wwz��}E3�v���Db*�|ЬV�axX?}
��}?yB��Z:#��hX:
����饣�h�U==D<���g�LL(�t?��7�"V���x��^CZ�Jpr,�'�z-���]3�5Ǣ�{ ����;�pLw������6)��B������T��*�i#Eb�ɾ����h�tz+�`��"*'�I���C��ȣJ�Z<��jxX+
���m��X�t/M�B
�c]Z_$֒_}�K)l���[,��L�����KV�h��YkNٮ�\�ʺ���	Ѓ��]k吠
p�2�
G��F�s�%h�Z:]u)
���ou���C�xv>�������}j�ƹ90���E3�[Z$��"3��m*�V�x-
)wT�b�Ѿ��饣�h�U��0�R<�������R&^E��kow�e������p���P�V|����2�T=�U-EBC�f�L�@�z!��Z+�[�p�PJ��x*�u(�X+
���;*��A��X�h�vz/���k�E;�Z����$���@�qX�DAOC����m��شt�f�D��W�j�gd;�5�q��}Jf)�f)��۳�\m������r�Z~jQ�%k�<��T'sQ�5�q��|`���GB��R�a�L��^�����ȴt>��S�аT/ONqG�m3�#�U����V
�eB;�����y盏1�s��v�UZ5UZ5UV�U[UUmUU�UV�U[UUh�UTmU�,��8gNuKc2�S���<çT6���'ms�9"�6HmL�X, p��@�i��կW��h�|'��l��R|��9�B�
ǣ�z2릖�ţ�Q�3s#�X��{7�P�t/]�G�"#�	RFۡ`�:v�P�4�r=�
�ea��X�V*��ꥣ��^�b5��<���=w�=T���#�T��PD
T��ذT.쓲��Ш^�������4�q�eR���T8�S��v�DTr�SOc�����$$�.��E��zo� X|���s盛�z,�֪~�x:
�K����f*)��I��v�O^j��c�X�@�aQe��_uM��Uy�易8��ˡ�k2�F�XՏF�^�-�GC��X*
����!�Z:R��`���ff<�o�V���s��e������YU���b�H�
6�1c�z�X�ݗ�R<��h��%B�},B�t��^��GK�A3��x*��-B �����[q�ꥦ$�I
ţ�wF��
G��T��]�G��֬��f��<׭M�q�̏�8����h�tz+�`�x+T�X�  �m�[�a�b9��������וU�ޱ���@�K�H��±]{��W�����O�C�`���z�h�zbu��1SSE3�S$�r��;mt���*������ֵ�N53xT����舏�X���r?{{u X+�Z<����P,B���!�Z:R�ł�o��R���G}�""����������C��T>,�*�X蛖�}���6�6�&��\z�~��nE��h�^.�dX*
����f��k�U���SX�Nt82I���-lf�@TNUZ���T.��d<)�ɴ�X�xd��]�G��Ъ}=B�X�twd��OD陘�*I��T?�Q"���X)
����z-o�{��!��H�c��:,H����DDDD@ DDDDDDDF�DDDD@ DDDDDL���K�nD/<{-V]���m�&�Ƌ����8D�q������GLӭ������qu�4v���<y3�'l�H>}W��l�)q=�����}}`�v=��* X.و�L�B��;�'r�hV�(���h�Q賦e`�x*z:/U-�GB��ł��_>���I��I��b�i����Y�	ԕ�N�<﯎���m��?v��3hzǭ�����b��z,���>!h�Z:R��`�x*�1]u=G���f����OH�y�ƺ���g���7L�%��'<s����l���8�D+�_�/EC�P��p���i��\�)�z�cU�l��j�Mw� j�R"4T<db�(.�`�x:*y{�ŧ�ġh�<NOEK�X�T-����Z<x����計pS7�E��������q֧���$�0z,O�z�h�Gb�Ϫ Z*5Z���z.=?t�Uce�[z�EB�9S+b�P���z�h�Z:OGRX;�Z9����Y?MET�S$�S$�m���\�.u���An�@��ǫ���}﬐�D�c��aU�jދ��E(�
ǂ���������TwM�<�b�Wl�GǢfg��=.E�����-Ѝ�>[>g�6���2"����G��{�;�-�GB�Ob�Z+��w��~5�t/E�щ�4����|j�Ƭ��m�!Q4�x-
���R��Q����E��T�����诩`�x+��޵� C�uFlQ��E� �B���^��Z;��龨C�P�#E��/����X������k��
J��EY2�A�kG"�Ъz'����������h�}=��
���y���|{d��f)�f)��t�h]/����l狝>�^wb�ɘ�u��|Ω�U�X@D
L�
ǂ�{��Դt=
�雘X)
��ٸ�ţ�x��c]��I�/sX��d��q&i12���F��HRB�l4������9����[UUmUU�UV�U[UUmUU�UU�UUmUU�UU`�#-�<c�:�+��m6X���mɼ�����:�i6���L�ɗ
n����W�z�Z����5�Y�.ki<��mm��|g"��^��V���m����R-�1Y"��S��v-�阈���ذW8�*?�%
��{�(z}��T�bM(X-����J�P�T*we�E�I��~���T���E�^Nf��"��EB��T!�x:*w�:�h��4v(�dGL-�B��ɧ�7�":`!E`�x+��P�C�ذV-Z|�b��V?��T�T<?N|B�$����1L�1L�2M��Vmûr�6i.�s5������~��\k�}�l>MX��5����m���]�=�;�J�z�A�3A�*�s�n6C�.lZZ��!-!--�Զ9qJ蛖�-$�m��3k��*�-��Uzyҷ�����UQ"T�u��<ʤ=2�m6�F�f���R�B!�I�5k���Kt_Z���;�Y�t	'�`(v���ڈ�!�x�P�o�Z*���}X�F�B�<�;��+(T�r�j*�ݟ��ԜR�W�Y���E�fO
z�{�$�p�FDS1m�u�9�e��c�U�]�]%������HG��ܹ�m�"��b�aE4�AЪX���� 5���skϜ�R���[c�9e�XQ�+cm����wطk����}�{�J����@��L��O1}���p�2d�����ҩkH�Qn�I�iΊ�A�){��ffz��B{|�g4�8�ta�^G��f�>������M�a ����[U��p����"""" �����"""#h����""" ����"""" ����"""""S(.�4�Z��� ��踢.�Ŝ������{H[��譵�\:�j��ch"�\��{u�G��qo5cak��b��J��%��R���m�K�c����E�{ח��X��陘�T�^��
���Z�d�h�bt��������z�O���f*)��I�۩ر��Q�{i��g2��Ie�̗��I$�mȚ933.�s뵈>ٸ���X�v�� +�E�� ������{BI����k����"���X���Dk뻳��z���V�3��Z�p�[;f�	���1ܑ�����Z\>����K�qr�t�|,�!�x�� P.�3��K.�}�EjRmL�kG���������Ob���7�93l˻��,wAKP��9Z:MLd��1L�E3�ݬ�z�c$�P��5����K��y���j;�e�dU�A���C��� +�Dsjn$��ˡbX��Ei{�_n�^�^�h�b�"\��͐h��쬳Wa�C=S�j�QBv�0�;}���$��x��!4�`a^���0O:{T~��ob����}T�Ξ������س��N6O��x���ƽT���=[�T����pGL!��R����h�;q׌c�7�Y����\��h( $3
*��p�FA�D�E2���s������E��=��7.a�� y6框���ww��Z���d[�a^�$���X��{���< ���<rY��x֯4��_wz�|{���ڪ�j������j�������ڪ�j���l�p�f�ܗ���iw-�e�z�m�k��"�Q��+4J�m
%,Pk]H�KI].%�/i$��i	il��A�'ch��kIA�&���N}|\�=�V��#��A�LQ���,B�w��E5�ܽ7��疴��K����}��ߎg"�K�}��9���$�_E&�iv��D��3mom�fٷ 9
@7��;adA� �#�S�i `�+cD�A���������A�ێ/kL�J�$��'Bi��V$����Q:����������!�8�u��d������r�*��� � �� m�q��PF�QB�����<�������E3�3�[t���؃4�!��̯xhu-��� �9����V+���V˼A�A�g4���m�4Q$�v�6�;A�Ŝ_�, � � � �m�l,ز������aq* � � � �^�q��A�ڸ�*�<^�+�A�ƴ���I�ܲ����[Յ�E*j� i�$!T"m$�i;OD��C�)s&8���� ���8�uo uo+�X8��usuo7��k"����UQD�Z\$��'�id�l[`H�K � � � �^��u������#����[R�����b���R�N-��� �A�A����q� �
o��UW�*�q��#h$�M-�ݶ `��OD����`�m���DD�@�6�q{qu�uq�1@A�,��k �quo6�b�ߋ��6��*#�(�si|&�n�$A_����~o�P�o� �EH%_W����;���{�>ئb���d�����	��Sط<���}/���>t86I�ɑ|������''9�o�)b�֢2T�j�0�� 3�)���z���)��F�����vyi��!8�g}{rd~���[��R(<2e(�3 ج��+qhB���e�����Cꦞ?W�^�V�}����S�zWj��f +3 �m�['.�ɝ���Obʬ�E�tnߚ�+R�Дd�%���Y�%�0$*Ģ�w��  6�D"bE�o\W���DDDF�� ����"""" ����"""6������"""6�����""#�""�ҙ��s��I���hw���W��h̝��:�3�O6�ň\kL@��!w$���6^g�3��+�͝YJD�Ċ�U�[%�Z���ik�_WҪ��T�Ϙ���#�\陀`�+1kF��Yv+��]������W�%�s~93�Z��z/��ae��YKb��gn�`��#4�De��Jsk{��t ���3�߹�>;�Wy������IR��!�Q���b���u��=z7tq�.�BZ[&*���w`��Lr��UQ��^�kj�H^l�I�'B)Ty���/,����cz��0²���:YO}_Wo��a�>t���Y��;5���62�#��ڞ����5��.��������� �����M��Uէ����@�[1��澯u�����阦I��b���m=v�=t�M=I���ke9f��g�@�L�o+�݋��%H^�H� GR�Q���=6\��=*�s�8^.i%9e-�%�����V-������ǿ�EH^l�I�'B)j���ݼ�ΒxR�8�� �".�&���y�����.��`��N�� �`�żU��y�M�m2>#�E�"�8:[��ﾥ�{�{�f���f�tj�vpݜA�l�>�����n��Y�/lY���=kZ�4ք��3%$��)l�TS$�s]W)�����C5Q$xnoz����?	��71s�7�c����]ʌ	�������c���	����U*<Z�������q�������$�I'�  
5j��� ��H��A����_���ƫL>6(�ܗ�@Sh �lG���#כX���{83`@h���d�87�c0�Ê�?�uB�@q�T��?�}ӗV?����'@U��=��Ϳ�����_ŧ�7g�F�}m�巍�}��}�$#�(�z6.X���U`�>s��6���̣�&��_�^��}���� ܻ������z�@Q���2aso��y���';'h|�ƀ��0x�M�ϻ��zj�����vz�
������k��������F{��	���l[��+��b2D�&z�н��D�O�ж�mv�x�.�<������~>��msh�o}�j"vm=�����j��aV mD�۫(�(�z`8���z-b���ŜA�U�X8�=~���@@r���k�	�5��y��q�6�4����|�������;s�׫�����>��6��i=S��U6�zr�}�\P�����KM��t�t��^)����?�Ƌם���x��a|7C�1&�}�E��9;��v�=���<s��}���:��4�~l_�>{���xZ{~92x� ����N����|<O�c>�v��yjv�{}��D��[�Q;� Q�
:�����ȇ�U,2n�/t��X�4e��<􀂍�PǪ9���ȱE��j���tM ��������bB������B<�R� bCP<QDw��`m/���[�N�2R��E'�]/��<yW����6G����PG���=��~9��'�������2Ʃ<?_���y��t��w�n}K븾�O����7;o��|���� �?��'���zM~ؠ�r��o|����9�� ��
)����
n�����xLX�:�>��:�c�ˬ����4�i�>a�r�:̆�e>ꇿ�|�!r�:md��.��c}ӗ���c��t�����Ю1�aѰ_���tx�&� (�����ͳn��B�%��m����o6�m�9���0�!����{v`�.'e��r/a�����P���;��0D�����e~���
<��=ncՠ�nC��~��6��mlp���Ϻ�CD$�~���g`���"�(HT�� 