BZh91AY&SYf�� B߀Px���������P�:81��i	D��!�h��4hѴ�I� 4 hz��h�        ��MS#�Q�4l�@b1�ѡ���A�ɓ&F�L�LD�"4�&*~�M'�y@�j46�@�#)�!	*��(B~��l��� ?�?�VhGk�;��%h�����g��B�U�����~�d��)�40��Y1��r]��)#���@�8�lᄊ��G����aԓ�"!njky�f��!,0� �>e�9�p c7#�CZ
]���e�T��oL�IRkC�-�g����ZX�� m
���F��.tG2�1
&M�Ҙ!�l���e\�CJ{�A͖�1PtAPE�s$3�Z��+i�p�V���h��$;IT�%�%���"���C�d�F�ddD���׹�Rmsv�
�;����&h��
���
I$� &#|��wbd� ;��t޻T�B���Ҋ�H�W,�TZbe���bI�1�z2���A,/k�Ť�����/�<�o�j�$�kJ�	\0������e�~��~���D��Rb%Z�����o^�a40���3)a�q��GI>���WD���&d0�TUA>��1žE�'nQ�P�dt� ��|�k7�g�^��,��(d(t#D�&��k��%b���M��8f=��������f�%#9�T5,�ҝ� �oZZpA ӭmC,�>$U\"�3OY�� `@24��kΚ�v����Hd�x��TQ��Ow��N�	�@[Y�E~�"�:���M[�QK/!�V�$w��'N����rb�G�&cs�4 \j�� `0fs~�uF=�)�	J(RJ�"Q���*s ���S&&2�������eE��&H��yCE.2�l����Q�#"�n��1���r��X��sʪ�TC5�ˀ&��mD� �
��i�^(���T�]��J�;�Q�V����0]�#��� $�b������f�c�~�p2�;�T0Ug%��&o��|Ml�v�f�9�,V9$W�o�v+)J�6{�W&���&0�Hڦ~��k�tj]�Å|X�כ���?��
�iW��&u,����l��N��t*�ɼ��	�RA�����H�
ӹ�`