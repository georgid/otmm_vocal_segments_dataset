BZh91AY&SY1� )_�Py���������`}�(i���     d ��WF�P+ZXDC3I䧩�D�P$����42O 5�S�0     2dɈ��	�����%=$��z�L�      (�	OD�2'�&OS5���@���!�mD��!��'�(�� 4�q�N|*((ڊ�x?�UFS���PI$$TO؊
��{��I%�����(����H+t�-��Mv�f���-��d�I��ͧ9Ͷ���m����oYm����m�m�M��i��0܆�-�u��ǧ�]=�ޮ��i�Ye��-�m�ލ��v;�{!���� g�g�m��Cm���[m���m�m�m�M�-����=�W\H14���Em|
�S�OnH�B0���m�n����3V]q�E5f���8PY(4��r�����8Li���H��0v�E�fNօod��V Q���2���\�K���;ͼQ�2�^�'T��-��w�P�6��0�obʻ�bF+�13�̣b*]f�%H;����v�ė�.b��KmC���}��k�.�<gfK�R$Lq��y�2j����0"l������,d--��Kq�1�c$��.{��=x�ZQ��9?��L�,T���Q�9���Nt�i�v����3?��ۻ����wwm��m��m��lcP�[J+�K�' Xv�f#���r��Vwu@�n&a�A����z���bgCc �2��2"��C>*	E��ǃV@U&�3�<�Jґ�*�  `���	Q���A��{WyW`��Gg��`�F��f��&�4��;�uT9��5��~�Q���ol	2��������ҩt��*~�ڋ`��k����V�KX��+�m�vfid�#"�
̛kek���΃�S�c������xr�q���|���� I�>$��g�E����Z�ɘ� �"I\�B<��Dk�� g�b`�&x{��m^!���U��<G�4G��-oR]2�*Z� #�=5[P"��Y���9 x�U524�����K=�y�w�d�4G�� 3/��fFK�_}US覺@��B�P�S��p�
-2NE��Qp�9�b0�L��n�JL\x�_���_"Ց_. �ɐ<C:D�bwsB��h�<
�A���S<��DG0�5�B9�q|y�����]�R����e�7�a] ���<�����r!C�A�a�8&���؆u3n�z�C�1�:y}��x����Rw��(V	�d#.�0btt��O+�О?fW ۼ	�+�y�9���t(���� �cĬ��]�^�rO)�־A"��ͥL?�Md�5� i���H?��������uߪ�Q�0oU��`�|�(Q���u3
o��6��[����ڮs]E���r���j���Sq4-u-���p<ܛ /��uX�t���;sJ���*�IdE�;�X��������;YU�z2rt>���X�M�Ws��s�:<�(鼑���~��e�����;Lĺ��7��"mV������xp%w�3�c2�Oe\�w�1Q�C�Y>؟����R
&L��������Wl��*��X���A���D~�$�W^P~���;�5b�X��E+���I5����%�y�U�ͼ����X�}���������ƅ���o�x� ^��r&�4�vg�o��������뾬�ȔDK�T���iH�����܃6�oB���LYR7���8";�+�M$���^��W��14Ay�&cH�w������}7�4����þ�>);��o��{��ﾬ��V�,�;U��͓v��]"��sDNB��=�8(�fY�N�x�=>�-�jED&bc�VWb~�{=�?��@�V���,��{_N��� ����G|���{�X�ց:�M�g�WiVv痕a��>ڱ�������Mf���_pa���P�遻�R���ԅ�����V9=�5�-gG�gۂ����z��,��� iha�*�ȵ�����Egn��A��
r��ط1�	�O8®�����߽Q!�s�E5�����)�<��V�\�GMZ��jӚßKH�K�U$�E���xÇ0��q(����./�����QS&�6V,ը�d��4j�αB1UE�*�"���EQZ05��V�TUUTTX"�������ETꨘ�V��j��-P�*bD��D�p�-��!h�7!$�8����b-�-(2�����YRЪ���R�\�,R9D}�-��\@Љ��(��|��8A!IP�M�u��*������ynX�
'T8U��wB����,�@"�j��,�7�~��b�(D�~~PXLu}�¡�]"�!�v��-=�Ё���zQU�`��h�	%0�x�u�}���H�<c+Dz��&@V�8=d4u��Nt��֞��EO�
���?Jy���� @�4�/@S��!O2w���"�$ H��2����d�%Z����4�׶X
�7N�V���-e�qL|s�v�L�`B�D
�Ҕ(Q�DA�F�iV�Z��!�*�	!$���f\��������l��X�'q}���4�;@Xdj�RRAI$�%|�ͼ:s12Ƃ�O*9��`̥�.%�0ݙ�9ؓ������s�"�>�eK=��ǟ�>ӣ��7�#b� �V2��ߔ�V�����&�1�15:�ɾ�^&ޜ|$���r��Z
�?�D��x2��-칵�&I�gIC#O�F�yL��<a�rv�-��7^b���U���b0�6�X�݀��&(~7�z���m��Y�h����C1��7x�-����7�#�Z��}�T
0B�뿋׸t�zP<~b����cT@v����t^�v���d̼������ݴ��k���;�:��Gk���\b��!��p@�<��\g7f��]�W�l�;�hc˪�ȑ�8�5b�0�Җ3�xP-4�5bdg�g�ՌG��
�\��m�%��K��a�g�����#���7�(Ko�!���nw�w�k���*��"�p����0�3	[�1�����a���s�W8+���w����SBP�aA���,ۑ*o6]�O��+!��eU�A��k�[���H�
=�@